VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO scan_wrapper_lesson_1
  CLASS BLOCK ;
  FOREIGN scan_wrapper_lesson_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 70.000 BY 70.000 ;
  PIN clk_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.570 66.000 68.130 70.000 ;
    END
  END clk_in
  PIN clk_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 0.000 32.710 4.000 ;
    END
  END clk_out
  PIN data_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 66.000 33.740 70.000 34.940 ;
    END
  END data_in
  PIN data_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.740 4.000 34.940 ;
    END
  END data_out
  PIN latch_enable_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -0.050 0.000 0.510 4.000 ;
    END
  END latch_enable_in
  PIN latch_enable_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -0.050 66.000 0.510 70.000 ;
    END
  END latch_enable_out
  PIN scan_select_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.370 66.000 35.930 70.000 ;
    END
  END scan_select_in
  PIN scan_select_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.570 0.000 68.130 4.000 ;
    END
  END scan_select_out
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 14.550 10.640 16.150 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 34.200 10.640 35.800 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 53.855 10.640 55.455 57.360 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.370 10.640 25.970 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 44.025 10.640 45.625 57.360 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 64.400 57.205 ;
      LAYER met1 ;
        RECT 0.070 10.640 68.010 57.360 ;
      LAYER met2 ;
        RECT 0.790 65.720 35.090 66.000 ;
        RECT 36.210 65.720 67.290 66.000 ;
        RECT 0.100 4.280 67.980 65.720 ;
        RECT 0.790 4.000 31.870 4.280 ;
        RECT 32.990 4.000 67.290 4.280 ;
      LAYER met3 ;
        RECT 4.000 35.340 66.000 57.285 ;
        RECT 4.400 33.340 65.600 35.340 ;
        RECT 4.000 10.715 66.000 33.340 ;
      LAYER met4 ;
        RECT 16.550 10.640 23.970 57.360 ;
        RECT 26.370 10.640 33.800 57.360 ;
        RECT 36.200 10.640 43.625 57.360 ;
        RECT 46.025 10.640 53.455 57.360 ;
  END
END scan_wrapper_lesson_1
END LIBRARY

