magic
tech sky130A
magscale 1 2
timestamp 1656598884
<< obsli1 >>
rect 17104 18159 547860 681425
<< obsm1 >>
rect 14 13064 580506 700732
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< obsm2 >>
rect 20 703464 8030 703610
rect 8254 703464 24222 703610
rect 24446 703464 40414 703610
rect 40638 703464 56698 703610
rect 56922 703464 72890 703610
rect 73114 703464 89082 703610
rect 89306 703464 105366 703610
rect 105590 703464 121558 703610
rect 121782 703464 137750 703610
rect 137974 703464 154034 703610
rect 154258 703464 170226 703610
rect 170450 703464 186418 703610
rect 186642 703464 202702 703610
rect 202926 703464 218894 703610
rect 219118 703464 235086 703610
rect 235310 703464 251370 703610
rect 251594 703464 267562 703610
rect 267786 703464 283754 703610
rect 283978 703464 300038 703610
rect 300262 703464 316230 703610
rect 316454 703464 332422 703610
rect 332646 703464 348706 703610
rect 348930 703464 364898 703610
rect 365122 703464 381090 703610
rect 381314 703464 397374 703610
rect 397598 703464 413566 703610
rect 413790 703464 429758 703610
rect 429982 703464 446042 703610
rect 446266 703464 462234 703610
rect 462458 703464 478426 703610
rect 478650 703464 494710 703610
rect 494934 703464 510902 703610
rect 511126 703464 527094 703610
rect 527318 703464 543378 703610
rect 543602 703464 559570 703610
rect 559794 703464 575762 703610
rect 575986 703464 580502 703610
rect 20 536 580502 703464
rect 20 326 486 536
rect 710 326 1590 536
rect 1814 326 2786 536
rect 3010 326 3982 536
rect 4206 326 5178 536
rect 5402 326 6374 536
rect 6598 326 7570 536
rect 7794 326 8674 536
rect 8898 326 9870 536
rect 10094 326 11066 536
rect 11290 326 12262 536
rect 12486 326 13458 536
rect 13682 326 14654 536
rect 14878 326 15850 536
rect 16074 326 16954 536
rect 17178 326 18150 536
rect 18374 326 19346 536
rect 19570 326 20542 536
rect 20766 326 21738 536
rect 21962 326 22934 536
rect 23158 326 24130 536
rect 24354 326 25234 536
rect 25458 326 26430 536
rect 26654 326 27626 536
rect 27850 326 28822 536
rect 29046 326 30018 536
rect 30242 326 31214 536
rect 31438 326 32318 536
rect 32542 326 33514 536
rect 33738 326 34710 536
rect 34934 326 35906 536
rect 36130 326 37102 536
rect 37326 326 38298 536
rect 38522 326 39494 536
rect 39718 326 40598 536
rect 40822 326 41794 536
rect 42018 326 42990 536
rect 43214 326 44186 536
rect 44410 326 45382 536
rect 45606 326 46578 536
rect 46802 326 47774 536
rect 47998 326 48878 536
rect 49102 326 50074 536
rect 50298 326 51270 536
rect 51494 326 52466 536
rect 52690 326 53662 536
rect 53886 326 54858 536
rect 55082 326 55962 536
rect 56186 326 57158 536
rect 57382 326 58354 536
rect 58578 326 59550 536
rect 59774 326 60746 536
rect 60970 326 61942 536
rect 62166 326 63138 536
rect 63362 326 64242 536
rect 64466 326 65438 536
rect 65662 326 66634 536
rect 66858 326 67830 536
rect 68054 326 69026 536
rect 69250 326 70222 536
rect 70446 326 71418 536
rect 71642 326 72522 536
rect 72746 326 73718 536
rect 73942 326 74914 536
rect 75138 326 76110 536
rect 76334 326 77306 536
rect 77530 326 78502 536
rect 78726 326 79606 536
rect 79830 326 80802 536
rect 81026 326 81998 536
rect 82222 326 83194 536
rect 83418 326 84390 536
rect 84614 326 85586 536
rect 85810 326 86782 536
rect 87006 326 87886 536
rect 88110 326 89082 536
rect 89306 326 90278 536
rect 90502 326 91474 536
rect 91698 326 92670 536
rect 92894 326 93866 536
rect 94090 326 95062 536
rect 95286 326 96166 536
rect 96390 326 97362 536
rect 97586 326 98558 536
rect 98782 326 99754 536
rect 99978 326 100950 536
rect 101174 326 102146 536
rect 102370 326 103250 536
rect 103474 326 104446 536
rect 104670 326 105642 536
rect 105866 326 106838 536
rect 107062 326 108034 536
rect 108258 326 109230 536
rect 109454 326 110426 536
rect 110650 326 111530 536
rect 111754 326 112726 536
rect 112950 326 113922 536
rect 114146 326 115118 536
rect 115342 326 116314 536
rect 116538 326 117510 536
rect 117734 326 118706 536
rect 118930 326 119810 536
rect 120034 326 121006 536
rect 121230 326 122202 536
rect 122426 326 123398 536
rect 123622 326 124594 536
rect 124818 326 125790 536
rect 126014 326 126894 536
rect 127118 326 128090 536
rect 128314 326 129286 536
rect 129510 326 130482 536
rect 130706 326 131678 536
rect 131902 326 132874 536
rect 133098 326 134070 536
rect 134294 326 135174 536
rect 135398 326 136370 536
rect 136594 326 137566 536
rect 137790 326 138762 536
rect 138986 326 139958 536
rect 140182 326 141154 536
rect 141378 326 142350 536
rect 142574 326 143454 536
rect 143678 326 144650 536
rect 144874 326 145846 536
rect 146070 326 147042 536
rect 147266 326 148238 536
rect 148462 326 149434 536
rect 149658 326 150538 536
rect 150762 326 151734 536
rect 151958 326 152930 536
rect 153154 326 154126 536
rect 154350 326 155322 536
rect 155546 326 156518 536
rect 156742 326 157714 536
rect 157938 326 158818 536
rect 159042 326 160014 536
rect 160238 326 161210 536
rect 161434 326 162406 536
rect 162630 326 163602 536
rect 163826 326 164798 536
rect 165022 326 165994 536
rect 166218 326 167098 536
rect 167322 326 168294 536
rect 168518 326 169490 536
rect 169714 326 170686 536
rect 170910 326 171882 536
rect 172106 326 173078 536
rect 173302 326 174182 536
rect 174406 326 175378 536
rect 175602 326 176574 536
rect 176798 326 177770 536
rect 177994 326 178966 536
rect 179190 326 180162 536
rect 180386 326 181358 536
rect 181582 326 182462 536
rect 182686 326 183658 536
rect 183882 326 184854 536
rect 185078 326 186050 536
rect 186274 326 187246 536
rect 187470 326 188442 536
rect 188666 326 189638 536
rect 189862 326 190742 536
rect 190966 326 191938 536
rect 192162 326 193134 536
rect 193358 326 194330 536
rect 194554 326 195526 536
rect 195750 326 196722 536
rect 196946 326 197826 536
rect 198050 326 199022 536
rect 199246 326 200218 536
rect 200442 326 201414 536
rect 201638 326 202610 536
rect 202834 326 203806 536
rect 204030 326 205002 536
rect 205226 326 206106 536
rect 206330 326 207302 536
rect 207526 326 208498 536
rect 208722 326 209694 536
rect 209918 326 210890 536
rect 211114 326 212086 536
rect 212310 326 213282 536
rect 213506 326 214386 536
rect 214610 326 215582 536
rect 215806 326 216778 536
rect 217002 326 217974 536
rect 218198 326 219170 536
rect 219394 326 220366 536
rect 220590 326 221470 536
rect 221694 326 222666 536
rect 222890 326 223862 536
rect 224086 326 225058 536
rect 225282 326 226254 536
rect 226478 326 227450 536
rect 227674 326 228646 536
rect 228870 326 229750 536
rect 229974 326 230946 536
rect 231170 326 232142 536
rect 232366 326 233338 536
rect 233562 326 234534 536
rect 234758 326 235730 536
rect 235954 326 236926 536
rect 237150 326 238030 536
rect 238254 326 239226 536
rect 239450 326 240422 536
rect 240646 326 241618 536
rect 241842 326 242814 536
rect 243038 326 244010 536
rect 244234 326 245114 536
rect 245338 326 246310 536
rect 246534 326 247506 536
rect 247730 326 248702 536
rect 248926 326 249898 536
rect 250122 326 251094 536
rect 251318 326 252290 536
rect 252514 326 253394 536
rect 253618 326 254590 536
rect 254814 326 255786 536
rect 256010 326 256982 536
rect 257206 326 258178 536
rect 258402 326 259374 536
rect 259598 326 260570 536
rect 260794 326 261674 536
rect 261898 326 262870 536
rect 263094 326 264066 536
rect 264290 326 265262 536
rect 265486 326 266458 536
rect 266682 326 267654 536
rect 267878 326 268758 536
rect 268982 326 269954 536
rect 270178 326 271150 536
rect 271374 326 272346 536
rect 272570 326 273542 536
rect 273766 326 274738 536
rect 274962 326 275934 536
rect 276158 326 277038 536
rect 277262 326 278234 536
rect 278458 326 279430 536
rect 279654 326 280626 536
rect 280850 326 281822 536
rect 282046 326 283018 536
rect 283242 326 284214 536
rect 284438 326 285318 536
rect 285542 326 286514 536
rect 286738 326 287710 536
rect 287934 326 288906 536
rect 289130 326 290102 536
rect 290326 326 291298 536
rect 291522 326 292494 536
rect 292718 326 293598 536
rect 293822 326 294794 536
rect 295018 326 295990 536
rect 296214 326 297186 536
rect 297410 326 298382 536
rect 298606 326 299578 536
rect 299802 326 300682 536
rect 300906 326 301878 536
rect 302102 326 303074 536
rect 303298 326 304270 536
rect 304494 326 305466 536
rect 305690 326 306662 536
rect 306886 326 307858 536
rect 308082 326 308962 536
rect 309186 326 310158 536
rect 310382 326 311354 536
rect 311578 326 312550 536
rect 312774 326 313746 536
rect 313970 326 314942 536
rect 315166 326 316138 536
rect 316362 326 317242 536
rect 317466 326 318438 536
rect 318662 326 319634 536
rect 319858 326 320830 536
rect 321054 326 322026 536
rect 322250 326 323222 536
rect 323446 326 324326 536
rect 324550 326 325522 536
rect 325746 326 326718 536
rect 326942 326 327914 536
rect 328138 326 329110 536
rect 329334 326 330306 536
rect 330530 326 331502 536
rect 331726 326 332606 536
rect 332830 326 333802 536
rect 334026 326 334998 536
rect 335222 326 336194 536
rect 336418 326 337390 536
rect 337614 326 338586 536
rect 338810 326 339782 536
rect 340006 326 340886 536
rect 341110 326 342082 536
rect 342306 326 343278 536
rect 343502 326 344474 536
rect 344698 326 345670 536
rect 345894 326 346866 536
rect 347090 326 347970 536
rect 348194 326 349166 536
rect 349390 326 350362 536
rect 350586 326 351558 536
rect 351782 326 352754 536
rect 352978 326 353950 536
rect 354174 326 355146 536
rect 355370 326 356250 536
rect 356474 326 357446 536
rect 357670 326 358642 536
rect 358866 326 359838 536
rect 360062 326 361034 536
rect 361258 326 362230 536
rect 362454 326 363426 536
rect 363650 326 364530 536
rect 364754 326 365726 536
rect 365950 326 366922 536
rect 367146 326 368118 536
rect 368342 326 369314 536
rect 369538 326 370510 536
rect 370734 326 371614 536
rect 371838 326 372810 536
rect 373034 326 374006 536
rect 374230 326 375202 536
rect 375426 326 376398 536
rect 376622 326 377594 536
rect 377818 326 378790 536
rect 379014 326 379894 536
rect 380118 326 381090 536
rect 381314 326 382286 536
rect 382510 326 383482 536
rect 383706 326 384678 536
rect 384902 326 385874 536
rect 386098 326 387070 536
rect 387294 326 388174 536
rect 388398 326 389370 536
rect 389594 326 390566 536
rect 390790 326 391762 536
rect 391986 326 392958 536
rect 393182 326 394154 536
rect 394378 326 395258 536
rect 395482 326 396454 536
rect 396678 326 397650 536
rect 397874 326 398846 536
rect 399070 326 400042 536
rect 400266 326 401238 536
rect 401462 326 402434 536
rect 402658 326 403538 536
rect 403762 326 404734 536
rect 404958 326 405930 536
rect 406154 326 407126 536
rect 407350 326 408322 536
rect 408546 326 409518 536
rect 409742 326 410714 536
rect 410938 326 411818 536
rect 412042 326 413014 536
rect 413238 326 414210 536
rect 414434 326 415406 536
rect 415630 326 416602 536
rect 416826 326 417798 536
rect 418022 326 418902 536
rect 419126 326 420098 536
rect 420322 326 421294 536
rect 421518 326 422490 536
rect 422714 326 423686 536
rect 423910 326 424882 536
rect 425106 326 426078 536
rect 426302 326 427182 536
rect 427406 326 428378 536
rect 428602 326 429574 536
rect 429798 326 430770 536
rect 430994 326 431966 536
rect 432190 326 433162 536
rect 433386 326 434358 536
rect 434582 326 435462 536
rect 435686 326 436658 536
rect 436882 326 437854 536
rect 438078 326 439050 536
rect 439274 326 440246 536
rect 440470 326 441442 536
rect 441666 326 442546 536
rect 442770 326 443742 536
rect 443966 326 444938 536
rect 445162 326 446134 536
rect 446358 326 447330 536
rect 447554 326 448526 536
rect 448750 326 449722 536
rect 449946 326 450826 536
rect 451050 326 452022 536
rect 452246 326 453218 536
rect 453442 326 454414 536
rect 454638 326 455610 536
rect 455834 326 456806 536
rect 457030 326 458002 536
rect 458226 326 459106 536
rect 459330 326 460302 536
rect 460526 326 461498 536
rect 461722 326 462694 536
rect 462918 326 463890 536
rect 464114 326 465086 536
rect 465310 326 466190 536
rect 466414 326 467386 536
rect 467610 326 468582 536
rect 468806 326 469778 536
rect 470002 326 470974 536
rect 471198 326 472170 536
rect 472394 326 473366 536
rect 473590 326 474470 536
rect 474694 326 475666 536
rect 475890 326 476862 536
rect 477086 326 478058 536
rect 478282 326 479254 536
rect 479478 326 480450 536
rect 480674 326 481646 536
rect 481870 326 482750 536
rect 482974 326 483946 536
rect 484170 326 485142 536
rect 485366 326 486338 536
rect 486562 326 487534 536
rect 487758 326 488730 536
rect 488954 326 489834 536
rect 490058 326 491030 536
rect 491254 326 492226 536
rect 492450 326 493422 536
rect 493646 326 494618 536
rect 494842 326 495814 536
rect 496038 326 497010 536
rect 497234 326 498114 536
rect 498338 326 499310 536
rect 499534 326 500506 536
rect 500730 326 501702 536
rect 501926 326 502898 536
rect 503122 326 504094 536
rect 504318 326 505290 536
rect 505514 326 506394 536
rect 506618 326 507590 536
rect 507814 326 508786 536
rect 509010 326 509982 536
rect 510206 326 511178 536
rect 511402 326 512374 536
rect 512598 326 513478 536
rect 513702 326 514674 536
rect 514898 326 515870 536
rect 516094 326 517066 536
rect 517290 326 518262 536
rect 518486 326 519458 536
rect 519682 326 520654 536
rect 520878 326 521758 536
rect 521982 326 522954 536
rect 523178 326 524150 536
rect 524374 326 525346 536
rect 525570 326 526542 536
rect 526766 326 527738 536
rect 527962 326 528934 536
rect 529158 326 530038 536
rect 530262 326 531234 536
rect 531458 326 532430 536
rect 532654 326 533626 536
rect 533850 326 534822 536
rect 535046 326 536018 536
rect 536242 326 537122 536
rect 537346 326 538318 536
rect 538542 326 539514 536
rect 539738 326 540710 536
rect 540934 326 541906 536
rect 542130 326 543102 536
rect 543326 326 544298 536
rect 544522 326 545402 536
rect 545626 326 546598 536
rect 546822 326 547794 536
rect 548018 326 548990 536
rect 549214 326 550186 536
rect 550410 326 551382 536
rect 551606 326 552578 536
rect 552802 326 553682 536
rect 553906 326 554878 536
rect 555102 326 556074 536
rect 556298 326 557270 536
rect 557494 326 558466 536
rect 558690 326 559662 536
rect 559886 326 560766 536
rect 560990 326 561962 536
rect 562186 326 563158 536
rect 563382 326 564354 536
rect 564578 326 565550 536
rect 565774 326 566746 536
rect 566970 326 567942 536
rect 568166 326 569046 536
rect 569270 326 570242 536
rect 570466 326 571438 536
rect 571662 326 572634 536
rect 572858 326 573830 536
rect 574054 326 575026 536
rect 575250 326 576222 536
rect 576446 326 577326 536
rect 577550 326 578522 536
rect 578746 326 579718 536
rect 579942 326 580502 536
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 583520 298604 584960 298844
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 583520 6476 584960 6716
<< obsm3 >>
rect 560 684084 583520 684317
rect 480 684076 583520 684084
rect 480 683676 583440 684076
rect 480 671428 583520 683676
rect 560 671028 583520 671428
rect 480 670884 583520 671028
rect 480 670484 583440 670884
rect 480 658372 583520 670484
rect 560 657972 583520 658372
rect 480 657556 583520 657972
rect 480 657156 583440 657556
rect 480 645316 583520 657156
rect 560 644916 583520 645316
rect 480 644228 583520 644916
rect 480 643828 583440 644228
rect 480 632260 583520 643828
rect 560 631860 583520 632260
rect 480 631036 583520 631860
rect 480 630636 583440 631036
rect 480 619340 583520 630636
rect 560 618940 583520 619340
rect 480 617708 583520 618940
rect 480 617308 583440 617708
rect 480 606284 583520 617308
rect 560 605884 583520 606284
rect 480 604380 583520 605884
rect 480 603980 583440 604380
rect 480 593228 583520 603980
rect 560 592828 583520 593228
rect 480 591188 583520 592828
rect 480 590788 583440 591188
rect 480 580172 583520 590788
rect 560 579772 583520 580172
rect 480 577860 583520 579772
rect 480 577460 583440 577860
rect 480 567116 583520 577460
rect 560 566716 583520 567116
rect 480 564532 583520 566716
rect 480 564132 583440 564532
rect 480 554060 583520 564132
rect 560 553660 583520 554060
rect 480 551340 583520 553660
rect 480 550940 583440 551340
rect 480 541004 583520 550940
rect 560 540604 583520 541004
rect 480 538012 583520 540604
rect 480 537612 583440 538012
rect 480 528084 583520 537612
rect 560 527684 583520 528084
rect 480 524684 583520 527684
rect 480 524284 583440 524684
rect 480 515028 583520 524284
rect 560 514628 583520 515028
rect 480 511492 583520 514628
rect 480 511092 583440 511492
rect 480 501972 583520 511092
rect 560 501572 583520 501972
rect 480 498164 583520 501572
rect 480 497764 583440 498164
rect 480 488916 583520 497764
rect 560 488516 583520 488916
rect 480 484836 583520 488516
rect 480 484436 583440 484836
rect 480 475860 583520 484436
rect 560 475460 583520 475860
rect 480 471644 583520 475460
rect 480 471244 583440 471644
rect 480 462804 583520 471244
rect 560 462404 583520 462804
rect 480 458316 583520 462404
rect 480 457916 583440 458316
rect 480 449748 583520 457916
rect 560 449348 583520 449748
rect 480 444988 583520 449348
rect 480 444588 583440 444988
rect 480 436828 583520 444588
rect 560 436428 583520 436828
rect 480 431796 583520 436428
rect 480 431396 583440 431796
rect 480 423772 583520 431396
rect 560 423372 583520 423772
rect 480 418468 583520 423372
rect 480 418068 583440 418468
rect 480 410716 583520 418068
rect 560 410316 583520 410716
rect 480 405140 583520 410316
rect 480 404740 583440 405140
rect 480 397660 583520 404740
rect 560 397260 583520 397660
rect 480 391948 583520 397260
rect 480 391548 583440 391948
rect 480 384604 583520 391548
rect 560 384204 583520 384604
rect 480 378620 583520 384204
rect 480 378220 583440 378620
rect 480 371548 583520 378220
rect 560 371148 583520 371548
rect 480 365292 583520 371148
rect 480 364892 583440 365292
rect 480 358628 583520 364892
rect 560 358228 583520 358628
rect 480 352100 583520 358228
rect 480 351700 583440 352100
rect 480 345572 583520 351700
rect 560 345172 583520 345572
rect 480 338772 583520 345172
rect 480 338372 583440 338772
rect 480 332516 583520 338372
rect 560 332116 583520 332516
rect 480 325444 583520 332116
rect 480 325044 583440 325444
rect 480 319460 583520 325044
rect 560 319060 583520 319460
rect 480 312252 583520 319060
rect 480 311852 583440 312252
rect 480 306404 583520 311852
rect 560 306004 583520 306404
rect 480 298924 583520 306004
rect 480 298524 583440 298924
rect 480 293348 583520 298524
rect 560 292948 583520 293348
rect 480 285596 583520 292948
rect 480 285196 583440 285596
rect 480 280292 583520 285196
rect 560 279892 583520 280292
rect 480 272404 583520 279892
rect 480 272004 583440 272404
rect 480 267372 583520 272004
rect 560 266972 583520 267372
rect 480 259076 583520 266972
rect 480 258676 583440 259076
rect 480 254316 583520 258676
rect 560 253916 583520 254316
rect 480 245748 583520 253916
rect 480 245348 583440 245748
rect 480 241260 583520 245348
rect 560 240860 583520 241260
rect 480 232556 583520 240860
rect 480 232156 583440 232556
rect 480 228204 583520 232156
rect 560 227804 583520 228204
rect 480 219228 583520 227804
rect 480 218828 583440 219228
rect 480 215148 583520 218828
rect 560 214748 583520 215148
rect 480 205900 583520 214748
rect 480 205500 583440 205900
rect 480 202092 583520 205500
rect 560 201692 583520 202092
rect 480 192708 583520 201692
rect 480 192308 583440 192708
rect 480 189036 583520 192308
rect 560 188636 583520 189036
rect 480 179380 583520 188636
rect 480 178980 583440 179380
rect 480 176116 583520 178980
rect 560 175716 583520 176116
rect 480 166052 583520 175716
rect 480 165652 583440 166052
rect 480 163060 583520 165652
rect 560 162660 583520 163060
rect 480 152860 583520 162660
rect 480 152460 583440 152860
rect 480 150004 583520 152460
rect 560 149604 583520 150004
rect 480 139532 583520 149604
rect 480 139132 583440 139532
rect 480 136948 583520 139132
rect 560 136548 583520 136948
rect 480 126204 583520 136548
rect 480 125804 583440 126204
rect 480 123892 583520 125804
rect 560 123492 583520 123892
rect 480 113012 583520 123492
rect 480 112612 583440 113012
rect 480 110836 583520 112612
rect 560 110436 583520 110836
rect 480 99684 583520 110436
rect 480 99284 583440 99684
rect 480 97780 583520 99284
rect 560 97380 583520 97780
rect 480 86356 583520 97380
rect 480 85956 583440 86356
rect 480 84860 583520 85956
rect 560 84460 583520 84860
rect 480 73164 583520 84460
rect 480 72764 583440 73164
rect 480 71804 583520 72764
rect 560 71404 583520 71804
rect 480 59836 583520 71404
rect 480 59436 583440 59836
rect 480 58748 583520 59436
rect 560 58348 583520 58748
rect 480 46508 583520 58348
rect 480 46108 583440 46508
rect 480 45692 583520 46108
rect 560 45292 583520 45692
rect 480 33316 583520 45292
rect 480 32916 583440 33316
rect 480 32636 583520 32916
rect 560 32236 583520 32636
rect 480 19988 583520 32236
rect 480 19588 583440 19988
rect 480 19580 583520 19588
rect 560 19180 583520 19580
rect 480 6796 583520 19180
rect 480 6660 583440 6796
rect 560 6427 583440 6660
<< metal4 >>
rect -2966 -1894 -2346 705830
rect -2006 -934 -1386 704870
rect 1794 -1894 2414 705830
rect 10794 -1894 11414 705830
rect 19794 686000 20414 705830
rect 28794 686000 29414 705830
rect 37794 686000 38414 705830
rect 46794 686000 47414 705830
rect 55794 686000 56414 705830
rect 64794 686000 65414 705830
rect 73794 686000 74414 705830
rect 82794 686000 83414 705830
rect 91794 686000 92414 705830
rect 100794 686000 101414 705830
rect 109794 686000 110414 705830
rect 118794 686000 119414 705830
rect 127794 686000 128414 705830
rect 136794 686000 137414 705830
rect 145794 686000 146414 705830
rect 154794 686000 155414 705830
rect 163794 686000 164414 705830
rect 172794 686000 173414 705830
rect 181794 686000 182414 705830
rect 190794 686000 191414 705830
rect 199794 686000 200414 705830
rect 208794 686000 209414 705830
rect 217794 686000 218414 705830
rect 226794 686000 227414 705830
rect 235794 686000 236414 705830
rect 244794 686000 245414 705830
rect 253794 686000 254414 705830
rect 262794 686000 263414 705830
rect 271794 686000 272414 705830
rect 280794 686000 281414 705830
rect 289794 686000 290414 705830
rect 298794 686000 299414 705830
rect 307794 686000 308414 705830
rect 316794 686000 317414 705830
rect 325794 686000 326414 705830
rect 334794 686000 335414 705830
rect 343794 686000 344414 705830
rect 352794 686000 353414 705830
rect 361794 686000 362414 705830
rect 370794 686000 371414 705830
rect 379794 686000 380414 705830
rect 388794 686000 389414 705830
rect 397794 686000 398414 705830
rect 406794 686000 407414 705830
rect 415794 686000 416414 705830
rect 424794 686000 425414 705830
rect 433794 686000 434414 705830
rect 442794 686000 443414 705830
rect 451794 686000 452414 705830
rect 460794 686000 461414 705830
rect 469794 686000 470414 705830
rect 478794 686000 479414 705830
rect 487794 686000 488414 705830
rect 496794 686000 497414 705830
rect 505794 686000 506414 705830
rect 514794 686000 515414 705830
rect 523794 686000 524414 705830
rect 532794 686000 533414 705830
rect 541794 686000 542414 705830
rect 550794 686000 551414 705830
rect 19794 659000 20414 662000
rect 28794 659000 29414 662000
rect 37794 659000 38414 662000
rect 46794 659000 47414 662000
rect 55794 659000 56414 662000
rect 64794 659000 65414 662000
rect 73794 659000 74414 662000
rect 82794 659000 83414 662000
rect 91794 659000 92414 662000
rect 100794 659000 101414 662000
rect 109794 659000 110414 662000
rect 118794 659000 119414 662000
rect 127794 659000 128414 662000
rect 136794 659000 137414 662000
rect 145794 659000 146414 662000
rect 154794 659000 155414 662000
rect 163794 659000 164414 662000
rect 172794 659000 173414 662000
rect 181794 659000 182414 662000
rect 190794 659000 191414 662000
rect 199794 659000 200414 662000
rect 208794 659000 209414 662000
rect 217794 659000 218414 662000
rect 226794 659000 227414 662000
rect 235794 659000 236414 662000
rect 244794 659000 245414 662000
rect 253794 659000 254414 662000
rect 262794 659000 263414 662000
rect 271794 659000 272414 662000
rect 280794 659000 281414 662000
rect 289794 659000 290414 662000
rect 298794 659000 299414 662000
rect 307794 659000 308414 662000
rect 316794 659000 317414 662000
rect 325794 659000 326414 662000
rect 334794 659000 335414 662000
rect 343794 659000 344414 662000
rect 352794 659000 353414 662000
rect 361794 659000 362414 662000
rect 370794 659000 371414 662000
rect 379794 659000 380414 662000
rect 388794 659000 389414 662000
rect 397794 659000 398414 662000
rect 406794 659000 407414 662000
rect 415794 659000 416414 662000
rect 424794 659000 425414 662000
rect 433794 659000 434414 662000
rect 442794 659000 443414 662000
rect 451794 659000 452414 662000
rect 460794 659000 461414 662000
rect 469794 659000 470414 662000
rect 478794 659000 479414 662000
rect 487794 659000 488414 662000
rect 496794 659000 497414 662000
rect 505794 659000 506414 662000
rect 514794 659000 515414 662000
rect 523794 659000 524414 662000
rect 532794 659000 533414 662000
rect 541794 659000 542414 662000
rect 550794 659000 551414 662000
rect 19794 632000 20414 635000
rect 28794 632000 29414 635000
rect 37794 632000 38414 635000
rect 46794 632000 47414 635000
rect 55794 632000 56414 635000
rect 64794 632000 65414 635000
rect 73794 632000 74414 635000
rect 82794 632000 83414 635000
rect 91794 632000 92414 635000
rect 100794 632000 101414 635000
rect 109794 632000 110414 635000
rect 118794 632000 119414 635000
rect 127794 632000 128414 635000
rect 136794 632000 137414 635000
rect 145794 632000 146414 635000
rect 154794 632000 155414 635000
rect 163794 632000 164414 635000
rect 172794 632000 173414 635000
rect 181794 632000 182414 635000
rect 190794 632000 191414 635000
rect 199794 632000 200414 635000
rect 208794 632000 209414 635000
rect 217794 632000 218414 635000
rect 226794 632000 227414 635000
rect 235794 632000 236414 635000
rect 244794 632000 245414 635000
rect 253794 632000 254414 635000
rect 262794 632000 263414 635000
rect 271794 632000 272414 635000
rect 280794 632000 281414 635000
rect 289794 632000 290414 635000
rect 298794 632000 299414 635000
rect 307794 632000 308414 635000
rect 316794 632000 317414 635000
rect 325794 632000 326414 635000
rect 334794 632000 335414 635000
rect 343794 632000 344414 635000
rect 352794 632000 353414 635000
rect 361794 632000 362414 635000
rect 370794 632000 371414 635000
rect 379794 632000 380414 635000
rect 388794 632000 389414 635000
rect 397794 632000 398414 635000
rect 406794 632000 407414 635000
rect 415794 632000 416414 635000
rect 424794 632000 425414 635000
rect 433794 632000 434414 635000
rect 442794 632000 443414 635000
rect 451794 632000 452414 635000
rect 460794 632000 461414 635000
rect 469794 632000 470414 635000
rect 478794 632000 479414 635000
rect 487794 632000 488414 635000
rect 496794 632000 497414 635000
rect 505794 632000 506414 635000
rect 514794 632000 515414 635000
rect 523794 632000 524414 635000
rect 532794 632000 533414 635000
rect 541794 632000 542414 635000
rect 550794 632000 551414 635000
rect 19794 605000 20414 608000
rect 28794 605000 29414 608000
rect 37794 605000 38414 608000
rect 46794 605000 47414 608000
rect 55794 605000 56414 608000
rect 64794 605000 65414 608000
rect 73794 605000 74414 608000
rect 82794 605000 83414 608000
rect 91794 605000 92414 608000
rect 100794 605000 101414 608000
rect 109794 605000 110414 608000
rect 118794 605000 119414 608000
rect 127794 605000 128414 608000
rect 136794 605000 137414 608000
rect 145794 605000 146414 608000
rect 154794 605000 155414 608000
rect 163794 605000 164414 608000
rect 172794 605000 173414 608000
rect 181794 605000 182414 608000
rect 190794 605000 191414 608000
rect 199794 605000 200414 608000
rect 208794 605000 209414 608000
rect 217794 605000 218414 608000
rect 226794 605000 227414 608000
rect 235794 605000 236414 608000
rect 244794 605000 245414 608000
rect 253794 605000 254414 608000
rect 262794 605000 263414 608000
rect 271794 605000 272414 608000
rect 280794 605000 281414 608000
rect 289794 605000 290414 608000
rect 298794 605000 299414 608000
rect 307794 605000 308414 608000
rect 316794 605000 317414 608000
rect 325794 605000 326414 608000
rect 334794 605000 335414 608000
rect 343794 605000 344414 608000
rect 352794 605000 353414 608000
rect 361794 605000 362414 608000
rect 370794 605000 371414 608000
rect 379794 605000 380414 608000
rect 388794 605000 389414 608000
rect 397794 605000 398414 608000
rect 406794 605000 407414 608000
rect 415794 605000 416414 608000
rect 424794 605000 425414 608000
rect 433794 605000 434414 608000
rect 442794 605000 443414 608000
rect 451794 605000 452414 608000
rect 460794 605000 461414 608000
rect 469794 605000 470414 608000
rect 478794 605000 479414 608000
rect 487794 605000 488414 608000
rect 496794 605000 497414 608000
rect 505794 605000 506414 608000
rect 514794 605000 515414 608000
rect 523794 605000 524414 608000
rect 532794 605000 533414 608000
rect 541794 605000 542414 608000
rect 550794 605000 551414 608000
rect 19794 578000 20414 581000
rect 28794 578000 29414 581000
rect 37794 578000 38414 581000
rect 46794 578000 47414 581000
rect 55794 578000 56414 581000
rect 64794 578000 65414 581000
rect 73794 578000 74414 581000
rect 82794 578000 83414 581000
rect 91794 578000 92414 581000
rect 100794 578000 101414 581000
rect 109794 578000 110414 581000
rect 118794 578000 119414 581000
rect 127794 578000 128414 581000
rect 136794 578000 137414 581000
rect 145794 578000 146414 581000
rect 154794 578000 155414 581000
rect 163794 578000 164414 581000
rect 172794 578000 173414 581000
rect 181794 578000 182414 581000
rect 190794 578000 191414 581000
rect 199794 578000 200414 581000
rect 208794 578000 209414 581000
rect 217794 578000 218414 581000
rect 226794 578000 227414 581000
rect 235794 578000 236414 581000
rect 244794 578000 245414 581000
rect 253794 578000 254414 581000
rect 262794 578000 263414 581000
rect 271794 578000 272414 581000
rect 280794 578000 281414 581000
rect 289794 578000 290414 581000
rect 298794 578000 299414 581000
rect 307794 578000 308414 581000
rect 316794 578000 317414 581000
rect 325794 578000 326414 581000
rect 334794 578000 335414 581000
rect 343794 578000 344414 581000
rect 352794 578000 353414 581000
rect 361794 578000 362414 581000
rect 370794 578000 371414 581000
rect 379794 578000 380414 581000
rect 388794 578000 389414 581000
rect 397794 578000 398414 581000
rect 406794 578000 407414 581000
rect 415794 578000 416414 581000
rect 424794 578000 425414 581000
rect 433794 578000 434414 581000
rect 442794 578000 443414 581000
rect 451794 578000 452414 581000
rect 460794 578000 461414 581000
rect 469794 578000 470414 581000
rect 478794 578000 479414 581000
rect 487794 578000 488414 581000
rect 496794 578000 497414 581000
rect 505794 578000 506414 581000
rect 514794 578000 515414 581000
rect 523794 578000 524414 581000
rect 532794 578000 533414 581000
rect 541794 578000 542414 581000
rect 550794 578000 551414 581000
rect 19794 551000 20414 554000
rect 28794 551000 29414 554000
rect 37794 551000 38414 554000
rect 46794 551000 47414 554000
rect 55794 551000 56414 554000
rect 64794 551000 65414 554000
rect 73794 551000 74414 554000
rect 82794 551000 83414 554000
rect 91794 551000 92414 554000
rect 100794 551000 101414 554000
rect 109794 551000 110414 554000
rect 118794 551000 119414 554000
rect 127794 551000 128414 554000
rect 136794 551000 137414 554000
rect 145794 551000 146414 554000
rect 154794 551000 155414 554000
rect 163794 551000 164414 554000
rect 172794 551000 173414 554000
rect 181794 551000 182414 554000
rect 190794 551000 191414 554000
rect 199794 551000 200414 554000
rect 208794 551000 209414 554000
rect 217794 551000 218414 554000
rect 226794 551000 227414 554000
rect 235794 551000 236414 554000
rect 244794 551000 245414 554000
rect 253794 551000 254414 554000
rect 262794 551000 263414 554000
rect 271794 551000 272414 554000
rect 280794 551000 281414 554000
rect 289794 551000 290414 554000
rect 298794 551000 299414 554000
rect 307794 551000 308414 554000
rect 316794 551000 317414 554000
rect 325794 551000 326414 554000
rect 334794 551000 335414 554000
rect 343794 551000 344414 554000
rect 352794 551000 353414 554000
rect 361794 551000 362414 554000
rect 370794 551000 371414 554000
rect 379794 551000 380414 554000
rect 388794 551000 389414 554000
rect 397794 551000 398414 554000
rect 406794 551000 407414 554000
rect 415794 551000 416414 554000
rect 424794 551000 425414 554000
rect 433794 551000 434414 554000
rect 442794 551000 443414 554000
rect 451794 551000 452414 554000
rect 460794 551000 461414 554000
rect 469794 551000 470414 554000
rect 478794 551000 479414 554000
rect 487794 551000 488414 554000
rect 496794 551000 497414 554000
rect 505794 551000 506414 554000
rect 514794 551000 515414 554000
rect 523794 551000 524414 554000
rect 532794 551000 533414 554000
rect 541794 551000 542414 554000
rect 550794 551000 551414 554000
rect 19794 524000 20414 527000
rect 28794 524000 29414 527000
rect 37794 524000 38414 527000
rect 46794 524000 47414 527000
rect 55794 524000 56414 527000
rect 64794 524000 65414 527000
rect 73794 524000 74414 527000
rect 82794 524000 83414 527000
rect 91794 524000 92414 527000
rect 100794 524000 101414 527000
rect 109794 524000 110414 527000
rect 118794 524000 119414 527000
rect 127794 524000 128414 527000
rect 136794 524000 137414 527000
rect 145794 524000 146414 527000
rect 154794 524000 155414 527000
rect 163794 524000 164414 527000
rect 172794 524000 173414 527000
rect 181794 524000 182414 527000
rect 190794 524000 191414 527000
rect 199794 524000 200414 527000
rect 208794 524000 209414 527000
rect 217794 524000 218414 527000
rect 226794 524000 227414 527000
rect 235794 524000 236414 527000
rect 244794 524000 245414 527000
rect 253794 524000 254414 527000
rect 262794 524000 263414 527000
rect 271794 524000 272414 527000
rect 280794 524000 281414 527000
rect 289794 524000 290414 527000
rect 298794 524000 299414 527000
rect 307794 524000 308414 527000
rect 316794 524000 317414 527000
rect 325794 524000 326414 527000
rect 334794 524000 335414 527000
rect 343794 524000 344414 527000
rect 352794 524000 353414 527000
rect 361794 524000 362414 527000
rect 370794 524000 371414 527000
rect 379794 524000 380414 527000
rect 388794 524000 389414 527000
rect 397794 524000 398414 527000
rect 406794 524000 407414 527000
rect 415794 524000 416414 527000
rect 424794 524000 425414 527000
rect 433794 524000 434414 527000
rect 442794 524000 443414 527000
rect 451794 524000 452414 527000
rect 460794 524000 461414 527000
rect 469794 524000 470414 527000
rect 478794 524000 479414 527000
rect 487794 524000 488414 527000
rect 496794 524000 497414 527000
rect 505794 524000 506414 527000
rect 514794 524000 515414 527000
rect 523794 524000 524414 527000
rect 532794 524000 533414 527000
rect 541794 524000 542414 527000
rect 550794 524000 551414 527000
rect 19794 497000 20414 500000
rect 28794 497000 29414 500000
rect 37794 497000 38414 500000
rect 46794 497000 47414 500000
rect 55794 497000 56414 500000
rect 64794 497000 65414 500000
rect 73794 497000 74414 500000
rect 82794 497000 83414 500000
rect 91794 497000 92414 500000
rect 100794 497000 101414 500000
rect 109794 497000 110414 500000
rect 118794 497000 119414 500000
rect 127794 497000 128414 500000
rect 136794 497000 137414 500000
rect 145794 497000 146414 500000
rect 154794 497000 155414 500000
rect 163794 497000 164414 500000
rect 172794 497000 173414 500000
rect 181794 497000 182414 500000
rect 190794 497000 191414 500000
rect 199794 497000 200414 500000
rect 208794 497000 209414 500000
rect 217794 497000 218414 500000
rect 226794 497000 227414 500000
rect 235794 497000 236414 500000
rect 244794 497000 245414 500000
rect 253794 497000 254414 500000
rect 262794 497000 263414 500000
rect 271794 497000 272414 500000
rect 280794 497000 281414 500000
rect 289794 497000 290414 500000
rect 298794 497000 299414 500000
rect 307794 497000 308414 500000
rect 316794 497000 317414 500000
rect 325794 497000 326414 500000
rect 334794 497000 335414 500000
rect 343794 497000 344414 500000
rect 352794 497000 353414 500000
rect 361794 497000 362414 500000
rect 370794 497000 371414 500000
rect 379794 497000 380414 500000
rect 388794 497000 389414 500000
rect 397794 497000 398414 500000
rect 406794 497000 407414 500000
rect 415794 497000 416414 500000
rect 424794 497000 425414 500000
rect 433794 497000 434414 500000
rect 442794 497000 443414 500000
rect 451794 497000 452414 500000
rect 460794 497000 461414 500000
rect 469794 497000 470414 500000
rect 478794 497000 479414 500000
rect 487794 497000 488414 500000
rect 496794 497000 497414 500000
rect 505794 497000 506414 500000
rect 514794 497000 515414 500000
rect 523794 497000 524414 500000
rect 532794 497000 533414 500000
rect 541794 497000 542414 500000
rect 550794 497000 551414 500000
rect 19794 470000 20414 473000
rect 28794 470000 29414 473000
rect 37794 470000 38414 473000
rect 46794 470000 47414 473000
rect 55794 470000 56414 473000
rect 64794 470000 65414 473000
rect 73794 470000 74414 473000
rect 82794 470000 83414 473000
rect 91794 470000 92414 473000
rect 100794 470000 101414 473000
rect 109794 470000 110414 473000
rect 118794 470000 119414 473000
rect 127794 470000 128414 473000
rect 136794 470000 137414 473000
rect 145794 470000 146414 473000
rect 154794 470000 155414 473000
rect 163794 470000 164414 473000
rect 172794 470000 173414 473000
rect 181794 470000 182414 473000
rect 190794 470000 191414 473000
rect 199794 470000 200414 473000
rect 208794 470000 209414 473000
rect 217794 470000 218414 473000
rect 226794 470000 227414 473000
rect 235794 470000 236414 473000
rect 244794 470000 245414 473000
rect 253794 470000 254414 473000
rect 262794 470000 263414 473000
rect 271794 470000 272414 473000
rect 280794 470000 281414 473000
rect 289794 470000 290414 473000
rect 298794 470000 299414 473000
rect 307794 470000 308414 473000
rect 316794 470000 317414 473000
rect 325794 470000 326414 473000
rect 334794 470000 335414 473000
rect 343794 470000 344414 473000
rect 352794 470000 353414 473000
rect 361794 470000 362414 473000
rect 370794 470000 371414 473000
rect 379794 470000 380414 473000
rect 388794 470000 389414 473000
rect 397794 470000 398414 473000
rect 406794 470000 407414 473000
rect 415794 470000 416414 473000
rect 424794 470000 425414 473000
rect 433794 470000 434414 473000
rect 442794 470000 443414 473000
rect 451794 470000 452414 473000
rect 460794 470000 461414 473000
rect 469794 470000 470414 473000
rect 478794 470000 479414 473000
rect 487794 470000 488414 473000
rect 496794 470000 497414 473000
rect 505794 470000 506414 473000
rect 514794 470000 515414 473000
rect 523794 470000 524414 473000
rect 532794 470000 533414 473000
rect 541794 470000 542414 473000
rect 550794 470000 551414 473000
rect 19794 443000 20414 446000
rect 28794 443000 29414 446000
rect 37794 443000 38414 446000
rect 46794 443000 47414 446000
rect 55794 443000 56414 446000
rect 64794 443000 65414 446000
rect 73794 443000 74414 446000
rect 82794 443000 83414 446000
rect 91794 443000 92414 446000
rect 100794 443000 101414 446000
rect 109794 443000 110414 446000
rect 118794 443000 119414 446000
rect 127794 443000 128414 446000
rect 136794 443000 137414 446000
rect 145794 443000 146414 446000
rect 154794 443000 155414 446000
rect 163794 443000 164414 446000
rect 172794 443000 173414 446000
rect 181794 443000 182414 446000
rect 190794 443000 191414 446000
rect 199794 443000 200414 446000
rect 208794 443000 209414 446000
rect 217794 443000 218414 446000
rect 226794 443000 227414 446000
rect 235794 443000 236414 446000
rect 244794 443000 245414 446000
rect 253794 443000 254414 446000
rect 262794 443000 263414 446000
rect 271794 443000 272414 446000
rect 280794 443000 281414 446000
rect 289794 443000 290414 446000
rect 298794 443000 299414 446000
rect 307794 443000 308414 446000
rect 316794 443000 317414 446000
rect 325794 443000 326414 446000
rect 334794 443000 335414 446000
rect 343794 443000 344414 446000
rect 352794 443000 353414 446000
rect 361794 443000 362414 446000
rect 370794 443000 371414 446000
rect 379794 443000 380414 446000
rect 388794 443000 389414 446000
rect 397794 443000 398414 446000
rect 406794 443000 407414 446000
rect 415794 443000 416414 446000
rect 424794 443000 425414 446000
rect 433794 443000 434414 446000
rect 442794 443000 443414 446000
rect 451794 443000 452414 446000
rect 460794 443000 461414 446000
rect 469794 443000 470414 446000
rect 478794 443000 479414 446000
rect 487794 443000 488414 446000
rect 496794 443000 497414 446000
rect 505794 443000 506414 446000
rect 514794 443000 515414 446000
rect 523794 443000 524414 446000
rect 532794 443000 533414 446000
rect 541794 443000 542414 446000
rect 550794 443000 551414 446000
rect 19794 416000 20414 419000
rect 28794 416000 29414 419000
rect 37794 416000 38414 419000
rect 46794 416000 47414 419000
rect 55794 416000 56414 419000
rect 64794 416000 65414 419000
rect 73794 416000 74414 419000
rect 82794 416000 83414 419000
rect 91794 416000 92414 419000
rect 100794 416000 101414 419000
rect 109794 416000 110414 419000
rect 118794 416000 119414 419000
rect 127794 416000 128414 419000
rect 136794 416000 137414 419000
rect 145794 416000 146414 419000
rect 154794 416000 155414 419000
rect 163794 416000 164414 419000
rect 172794 416000 173414 419000
rect 181794 416000 182414 419000
rect 190794 416000 191414 419000
rect 199794 416000 200414 419000
rect 208794 416000 209414 419000
rect 217794 416000 218414 419000
rect 226794 416000 227414 419000
rect 235794 416000 236414 419000
rect 244794 416000 245414 419000
rect 253794 416000 254414 419000
rect 262794 416000 263414 419000
rect 271794 416000 272414 419000
rect 280794 416000 281414 419000
rect 289794 416000 290414 419000
rect 298794 416000 299414 419000
rect 307794 416000 308414 419000
rect 316794 416000 317414 419000
rect 325794 416000 326414 419000
rect 334794 416000 335414 419000
rect 343794 416000 344414 419000
rect 352794 416000 353414 419000
rect 361794 416000 362414 419000
rect 370794 416000 371414 419000
rect 379794 416000 380414 419000
rect 388794 416000 389414 419000
rect 397794 416000 398414 419000
rect 406794 416000 407414 419000
rect 415794 416000 416414 419000
rect 424794 416000 425414 419000
rect 433794 416000 434414 419000
rect 442794 416000 443414 419000
rect 451794 416000 452414 419000
rect 460794 416000 461414 419000
rect 469794 416000 470414 419000
rect 478794 416000 479414 419000
rect 487794 416000 488414 419000
rect 496794 416000 497414 419000
rect 505794 416000 506414 419000
rect 514794 416000 515414 419000
rect 523794 416000 524414 419000
rect 532794 416000 533414 419000
rect 541794 416000 542414 419000
rect 550794 416000 551414 419000
rect 19794 389000 20414 392000
rect 28794 389000 29414 392000
rect 37794 389000 38414 392000
rect 46794 389000 47414 392000
rect 55794 389000 56414 392000
rect 64794 389000 65414 392000
rect 73794 389000 74414 392000
rect 82794 389000 83414 392000
rect 91794 389000 92414 392000
rect 100794 389000 101414 392000
rect 109794 389000 110414 392000
rect 118794 389000 119414 392000
rect 127794 389000 128414 392000
rect 136794 389000 137414 392000
rect 145794 389000 146414 392000
rect 154794 389000 155414 392000
rect 163794 389000 164414 392000
rect 172794 389000 173414 392000
rect 181794 389000 182414 392000
rect 190794 389000 191414 392000
rect 199794 389000 200414 392000
rect 208794 389000 209414 392000
rect 217794 389000 218414 392000
rect 226794 389000 227414 392000
rect 235794 389000 236414 392000
rect 244794 389000 245414 392000
rect 253794 389000 254414 392000
rect 262794 389000 263414 392000
rect 271794 389000 272414 392000
rect 280794 389000 281414 392000
rect 289794 389000 290414 392000
rect 298794 389000 299414 392000
rect 307794 389000 308414 392000
rect 316794 389000 317414 392000
rect 325794 389000 326414 392000
rect 334794 389000 335414 392000
rect 343794 389000 344414 392000
rect 352794 389000 353414 392000
rect 361794 389000 362414 392000
rect 370794 389000 371414 392000
rect 379794 389000 380414 392000
rect 388794 389000 389414 392000
rect 397794 389000 398414 392000
rect 406794 389000 407414 392000
rect 415794 389000 416414 392000
rect 424794 389000 425414 392000
rect 433794 389000 434414 392000
rect 442794 389000 443414 392000
rect 451794 389000 452414 392000
rect 460794 389000 461414 392000
rect 469794 389000 470414 392000
rect 478794 389000 479414 392000
rect 487794 389000 488414 392000
rect 496794 389000 497414 392000
rect 505794 389000 506414 392000
rect 514794 389000 515414 392000
rect 523794 389000 524414 392000
rect 532794 389000 533414 392000
rect 541794 389000 542414 392000
rect 550794 389000 551414 392000
rect 19794 362000 20414 365000
rect 28794 362000 29414 365000
rect 37794 362000 38414 365000
rect 46794 362000 47414 365000
rect 55794 362000 56414 365000
rect 64794 362000 65414 365000
rect 73794 362000 74414 365000
rect 82794 362000 83414 365000
rect 91794 362000 92414 365000
rect 100794 362000 101414 365000
rect 109794 362000 110414 365000
rect 118794 362000 119414 365000
rect 127794 362000 128414 365000
rect 136794 362000 137414 365000
rect 145794 362000 146414 365000
rect 154794 362000 155414 365000
rect 163794 362000 164414 365000
rect 172794 362000 173414 365000
rect 181794 362000 182414 365000
rect 190794 362000 191414 365000
rect 199794 362000 200414 365000
rect 208794 362000 209414 365000
rect 217794 362000 218414 365000
rect 226794 362000 227414 365000
rect 235794 362000 236414 365000
rect 244794 362000 245414 365000
rect 253794 362000 254414 365000
rect 262794 362000 263414 365000
rect 271794 362000 272414 365000
rect 280794 362000 281414 365000
rect 289794 362000 290414 365000
rect 298794 362000 299414 365000
rect 307794 362000 308414 365000
rect 316794 362000 317414 365000
rect 325794 362000 326414 365000
rect 334794 362000 335414 365000
rect 343794 362000 344414 365000
rect 352794 362000 353414 365000
rect 361794 362000 362414 365000
rect 370794 362000 371414 365000
rect 379794 362000 380414 365000
rect 388794 362000 389414 365000
rect 397794 362000 398414 365000
rect 406794 362000 407414 365000
rect 415794 362000 416414 365000
rect 424794 362000 425414 365000
rect 433794 362000 434414 365000
rect 442794 362000 443414 365000
rect 451794 362000 452414 365000
rect 460794 362000 461414 365000
rect 469794 362000 470414 365000
rect 478794 362000 479414 365000
rect 487794 362000 488414 365000
rect 496794 362000 497414 365000
rect 505794 362000 506414 365000
rect 514794 362000 515414 365000
rect 523794 362000 524414 365000
rect 532794 362000 533414 365000
rect 541794 362000 542414 365000
rect 550794 362000 551414 365000
rect 19794 335000 20414 338000
rect 28794 335000 29414 338000
rect 37794 335000 38414 338000
rect 46794 335000 47414 338000
rect 55794 335000 56414 338000
rect 64794 335000 65414 338000
rect 73794 335000 74414 338000
rect 82794 335000 83414 338000
rect 91794 335000 92414 338000
rect 100794 335000 101414 338000
rect 109794 335000 110414 338000
rect 118794 335000 119414 338000
rect 127794 335000 128414 338000
rect 136794 335000 137414 338000
rect 145794 335000 146414 338000
rect 154794 335000 155414 338000
rect 163794 335000 164414 338000
rect 172794 335000 173414 338000
rect 181794 335000 182414 338000
rect 190794 335000 191414 338000
rect 199794 335000 200414 338000
rect 208794 335000 209414 338000
rect 217794 335000 218414 338000
rect 226794 335000 227414 338000
rect 235794 335000 236414 338000
rect 244794 335000 245414 338000
rect 253794 335000 254414 338000
rect 262794 335000 263414 338000
rect 271794 335000 272414 338000
rect 280794 335000 281414 338000
rect 289794 335000 290414 338000
rect 298794 335000 299414 338000
rect 307794 335000 308414 338000
rect 316794 335000 317414 338000
rect 325794 335000 326414 338000
rect 334794 335000 335414 338000
rect 343794 335000 344414 338000
rect 352794 335000 353414 338000
rect 361794 335000 362414 338000
rect 370794 335000 371414 338000
rect 379794 335000 380414 338000
rect 388794 335000 389414 338000
rect 397794 335000 398414 338000
rect 406794 335000 407414 338000
rect 415794 335000 416414 338000
rect 424794 335000 425414 338000
rect 433794 335000 434414 338000
rect 442794 335000 443414 338000
rect 451794 335000 452414 338000
rect 460794 335000 461414 338000
rect 469794 335000 470414 338000
rect 478794 335000 479414 338000
rect 487794 335000 488414 338000
rect 496794 335000 497414 338000
rect 505794 335000 506414 338000
rect 514794 335000 515414 338000
rect 523794 335000 524414 338000
rect 532794 335000 533414 338000
rect 541794 335000 542414 338000
rect 550794 335000 551414 338000
rect 19794 308000 20414 311000
rect 28794 308000 29414 311000
rect 37794 308000 38414 311000
rect 46794 308000 47414 311000
rect 55794 308000 56414 311000
rect 64794 308000 65414 311000
rect 73794 308000 74414 311000
rect 82794 308000 83414 311000
rect 91794 308000 92414 311000
rect 100794 308000 101414 311000
rect 109794 308000 110414 311000
rect 118794 308000 119414 311000
rect 127794 308000 128414 311000
rect 136794 308000 137414 311000
rect 145794 308000 146414 311000
rect 154794 308000 155414 311000
rect 163794 308000 164414 311000
rect 172794 308000 173414 311000
rect 181794 308000 182414 311000
rect 190794 308000 191414 311000
rect 199794 308000 200414 311000
rect 208794 308000 209414 311000
rect 217794 308000 218414 311000
rect 226794 308000 227414 311000
rect 235794 308000 236414 311000
rect 244794 308000 245414 311000
rect 253794 308000 254414 311000
rect 262794 308000 263414 311000
rect 271794 308000 272414 311000
rect 280794 308000 281414 311000
rect 289794 308000 290414 311000
rect 298794 308000 299414 311000
rect 307794 308000 308414 311000
rect 316794 308000 317414 311000
rect 325794 308000 326414 311000
rect 334794 308000 335414 311000
rect 343794 308000 344414 311000
rect 352794 308000 353414 311000
rect 361794 308000 362414 311000
rect 370794 308000 371414 311000
rect 379794 308000 380414 311000
rect 388794 308000 389414 311000
rect 397794 308000 398414 311000
rect 406794 308000 407414 311000
rect 415794 308000 416414 311000
rect 424794 308000 425414 311000
rect 433794 308000 434414 311000
rect 442794 308000 443414 311000
rect 451794 308000 452414 311000
rect 460794 308000 461414 311000
rect 469794 308000 470414 311000
rect 478794 308000 479414 311000
rect 487794 308000 488414 311000
rect 496794 308000 497414 311000
rect 505794 308000 506414 311000
rect 514794 308000 515414 311000
rect 523794 308000 524414 311000
rect 532794 308000 533414 311000
rect 541794 308000 542414 311000
rect 550794 308000 551414 311000
rect 19794 281000 20414 284000
rect 28794 281000 29414 284000
rect 37794 281000 38414 284000
rect 46794 281000 47414 284000
rect 55794 281000 56414 284000
rect 64794 281000 65414 284000
rect 73794 281000 74414 284000
rect 82794 281000 83414 284000
rect 91794 281000 92414 284000
rect 100794 281000 101414 284000
rect 109794 281000 110414 284000
rect 118794 281000 119414 284000
rect 127794 281000 128414 284000
rect 136794 281000 137414 284000
rect 145794 281000 146414 284000
rect 154794 281000 155414 284000
rect 163794 281000 164414 284000
rect 172794 281000 173414 284000
rect 181794 281000 182414 284000
rect 190794 281000 191414 284000
rect 199794 281000 200414 284000
rect 208794 281000 209414 284000
rect 217794 281000 218414 284000
rect 226794 281000 227414 284000
rect 235794 281000 236414 284000
rect 244794 281000 245414 284000
rect 253794 281000 254414 284000
rect 262794 281000 263414 284000
rect 271794 281000 272414 284000
rect 280794 281000 281414 284000
rect 289794 281000 290414 284000
rect 298794 281000 299414 284000
rect 307794 281000 308414 284000
rect 316794 281000 317414 284000
rect 325794 281000 326414 284000
rect 334794 281000 335414 284000
rect 343794 281000 344414 284000
rect 352794 281000 353414 284000
rect 361794 281000 362414 284000
rect 370794 281000 371414 284000
rect 379794 281000 380414 284000
rect 388794 281000 389414 284000
rect 397794 281000 398414 284000
rect 406794 281000 407414 284000
rect 415794 281000 416414 284000
rect 424794 281000 425414 284000
rect 433794 281000 434414 284000
rect 442794 281000 443414 284000
rect 451794 281000 452414 284000
rect 460794 281000 461414 284000
rect 469794 281000 470414 284000
rect 478794 281000 479414 284000
rect 487794 281000 488414 284000
rect 496794 281000 497414 284000
rect 505794 281000 506414 284000
rect 514794 281000 515414 284000
rect 523794 281000 524414 284000
rect 532794 281000 533414 284000
rect 541794 281000 542414 284000
rect 550794 281000 551414 284000
rect 19794 254000 20414 257000
rect 28794 254000 29414 257000
rect 37794 254000 38414 257000
rect 46794 254000 47414 257000
rect 55794 254000 56414 257000
rect 64794 254000 65414 257000
rect 73794 254000 74414 257000
rect 82794 254000 83414 257000
rect 91794 254000 92414 257000
rect 100794 254000 101414 257000
rect 109794 254000 110414 257000
rect 118794 254000 119414 257000
rect 127794 254000 128414 257000
rect 136794 254000 137414 257000
rect 145794 254000 146414 257000
rect 154794 254000 155414 257000
rect 163794 254000 164414 257000
rect 172794 254000 173414 257000
rect 181794 254000 182414 257000
rect 190794 254000 191414 257000
rect 199794 254000 200414 257000
rect 208794 254000 209414 257000
rect 217794 254000 218414 257000
rect 226794 254000 227414 257000
rect 235794 254000 236414 257000
rect 244794 254000 245414 257000
rect 253794 254000 254414 257000
rect 262794 254000 263414 257000
rect 271794 254000 272414 257000
rect 280794 254000 281414 257000
rect 289794 254000 290414 257000
rect 298794 254000 299414 257000
rect 307794 254000 308414 257000
rect 316794 254000 317414 257000
rect 325794 254000 326414 257000
rect 334794 254000 335414 257000
rect 343794 254000 344414 257000
rect 352794 254000 353414 257000
rect 361794 254000 362414 257000
rect 370794 254000 371414 257000
rect 379794 254000 380414 257000
rect 388794 254000 389414 257000
rect 397794 254000 398414 257000
rect 406794 254000 407414 257000
rect 415794 254000 416414 257000
rect 424794 254000 425414 257000
rect 433794 254000 434414 257000
rect 442794 254000 443414 257000
rect 451794 254000 452414 257000
rect 460794 254000 461414 257000
rect 469794 254000 470414 257000
rect 478794 254000 479414 257000
rect 487794 254000 488414 257000
rect 496794 254000 497414 257000
rect 505794 254000 506414 257000
rect 514794 254000 515414 257000
rect 523794 254000 524414 257000
rect 532794 254000 533414 257000
rect 541794 254000 542414 257000
rect 550794 254000 551414 257000
rect 19794 227000 20414 230000
rect 28794 227000 29414 230000
rect 37794 227000 38414 230000
rect 46794 227000 47414 230000
rect 55794 227000 56414 230000
rect 64794 227000 65414 230000
rect 73794 227000 74414 230000
rect 82794 227000 83414 230000
rect 91794 227000 92414 230000
rect 100794 227000 101414 230000
rect 109794 227000 110414 230000
rect 118794 227000 119414 230000
rect 127794 227000 128414 230000
rect 136794 227000 137414 230000
rect 145794 227000 146414 230000
rect 154794 227000 155414 230000
rect 163794 227000 164414 230000
rect 172794 227000 173414 230000
rect 181794 227000 182414 230000
rect 190794 227000 191414 230000
rect 199794 227000 200414 230000
rect 208794 227000 209414 230000
rect 217794 227000 218414 230000
rect 226794 227000 227414 230000
rect 235794 227000 236414 230000
rect 244794 227000 245414 230000
rect 253794 227000 254414 230000
rect 262794 227000 263414 230000
rect 271794 227000 272414 230000
rect 280794 227000 281414 230000
rect 289794 227000 290414 230000
rect 298794 227000 299414 230000
rect 307794 227000 308414 230000
rect 316794 227000 317414 230000
rect 325794 227000 326414 230000
rect 334794 227000 335414 230000
rect 343794 227000 344414 230000
rect 352794 227000 353414 230000
rect 361794 227000 362414 230000
rect 370794 227000 371414 230000
rect 379794 227000 380414 230000
rect 388794 227000 389414 230000
rect 397794 227000 398414 230000
rect 406794 227000 407414 230000
rect 415794 227000 416414 230000
rect 424794 227000 425414 230000
rect 433794 227000 434414 230000
rect 442794 227000 443414 230000
rect 451794 227000 452414 230000
rect 460794 227000 461414 230000
rect 469794 227000 470414 230000
rect 478794 227000 479414 230000
rect 487794 227000 488414 230000
rect 496794 227000 497414 230000
rect 505794 227000 506414 230000
rect 514794 227000 515414 230000
rect 523794 227000 524414 230000
rect 532794 227000 533414 230000
rect 541794 227000 542414 230000
rect 550794 227000 551414 230000
rect 19794 200000 20414 203000
rect 28794 200000 29414 203000
rect 37794 200000 38414 203000
rect 46794 200000 47414 203000
rect 55794 200000 56414 203000
rect 64794 200000 65414 203000
rect 73794 200000 74414 203000
rect 82794 200000 83414 203000
rect 91794 200000 92414 203000
rect 100794 200000 101414 203000
rect 109794 200000 110414 203000
rect 118794 200000 119414 203000
rect 127794 200000 128414 203000
rect 136794 200000 137414 203000
rect 145794 200000 146414 203000
rect 154794 200000 155414 203000
rect 163794 200000 164414 203000
rect 172794 200000 173414 203000
rect 181794 200000 182414 203000
rect 190794 200000 191414 203000
rect 199794 200000 200414 203000
rect 208794 200000 209414 203000
rect 217794 200000 218414 203000
rect 226794 200000 227414 203000
rect 235794 200000 236414 203000
rect 244794 200000 245414 203000
rect 253794 200000 254414 203000
rect 262794 200000 263414 203000
rect 271794 200000 272414 203000
rect 280794 200000 281414 203000
rect 289794 200000 290414 203000
rect 298794 200000 299414 203000
rect 307794 200000 308414 203000
rect 316794 200000 317414 203000
rect 325794 200000 326414 203000
rect 334794 200000 335414 203000
rect 343794 200000 344414 203000
rect 352794 200000 353414 203000
rect 361794 200000 362414 203000
rect 370794 200000 371414 203000
rect 379794 200000 380414 203000
rect 388794 200000 389414 203000
rect 397794 200000 398414 203000
rect 406794 200000 407414 203000
rect 415794 200000 416414 203000
rect 424794 200000 425414 203000
rect 433794 200000 434414 203000
rect 442794 200000 443414 203000
rect 451794 200000 452414 203000
rect 460794 200000 461414 203000
rect 469794 200000 470414 203000
rect 478794 200000 479414 203000
rect 487794 200000 488414 203000
rect 496794 200000 497414 203000
rect 505794 200000 506414 203000
rect 514794 200000 515414 203000
rect 523794 200000 524414 203000
rect 532794 200000 533414 203000
rect 541794 200000 542414 203000
rect 550794 200000 551414 203000
rect 19794 173000 20414 176000
rect 28794 173000 29414 176000
rect 37794 173000 38414 176000
rect 46794 173000 47414 176000
rect 55794 173000 56414 176000
rect 64794 173000 65414 176000
rect 73794 173000 74414 176000
rect 82794 173000 83414 176000
rect 91794 173000 92414 176000
rect 100794 173000 101414 176000
rect 109794 173000 110414 176000
rect 118794 173000 119414 176000
rect 127794 173000 128414 176000
rect 136794 173000 137414 176000
rect 145794 173000 146414 176000
rect 154794 173000 155414 176000
rect 163794 173000 164414 176000
rect 172794 173000 173414 176000
rect 181794 173000 182414 176000
rect 190794 173000 191414 176000
rect 199794 173000 200414 176000
rect 208794 173000 209414 176000
rect 217794 173000 218414 176000
rect 226794 173000 227414 176000
rect 235794 173000 236414 176000
rect 244794 173000 245414 176000
rect 253794 173000 254414 176000
rect 262794 173000 263414 176000
rect 271794 173000 272414 176000
rect 280794 173000 281414 176000
rect 289794 173000 290414 176000
rect 298794 173000 299414 176000
rect 307794 173000 308414 176000
rect 316794 173000 317414 176000
rect 325794 173000 326414 176000
rect 334794 173000 335414 176000
rect 343794 173000 344414 176000
rect 352794 173000 353414 176000
rect 361794 173000 362414 176000
rect 370794 173000 371414 176000
rect 379794 173000 380414 176000
rect 388794 173000 389414 176000
rect 397794 173000 398414 176000
rect 406794 173000 407414 176000
rect 415794 173000 416414 176000
rect 424794 173000 425414 176000
rect 433794 173000 434414 176000
rect 442794 173000 443414 176000
rect 451794 173000 452414 176000
rect 460794 173000 461414 176000
rect 469794 173000 470414 176000
rect 478794 173000 479414 176000
rect 487794 173000 488414 176000
rect 496794 173000 497414 176000
rect 505794 173000 506414 176000
rect 514794 173000 515414 176000
rect 523794 173000 524414 176000
rect 532794 173000 533414 176000
rect 541794 173000 542414 176000
rect 550794 173000 551414 176000
rect 19794 146000 20414 149000
rect 28794 146000 29414 149000
rect 37794 146000 38414 149000
rect 46794 146000 47414 149000
rect 55794 146000 56414 149000
rect 64794 146000 65414 149000
rect 73794 146000 74414 149000
rect 82794 146000 83414 149000
rect 91794 146000 92414 149000
rect 100794 146000 101414 149000
rect 109794 146000 110414 149000
rect 118794 146000 119414 149000
rect 127794 146000 128414 149000
rect 136794 146000 137414 149000
rect 145794 146000 146414 149000
rect 154794 146000 155414 149000
rect 163794 146000 164414 149000
rect 172794 146000 173414 149000
rect 181794 146000 182414 149000
rect 190794 146000 191414 149000
rect 199794 146000 200414 149000
rect 208794 146000 209414 149000
rect 217794 146000 218414 149000
rect 226794 146000 227414 149000
rect 235794 146000 236414 149000
rect 244794 146000 245414 149000
rect 253794 146000 254414 149000
rect 262794 146000 263414 149000
rect 271794 146000 272414 149000
rect 280794 146000 281414 149000
rect 289794 146000 290414 149000
rect 298794 146000 299414 149000
rect 307794 146000 308414 149000
rect 316794 146000 317414 149000
rect 325794 146000 326414 149000
rect 334794 146000 335414 149000
rect 343794 146000 344414 149000
rect 352794 146000 353414 149000
rect 361794 146000 362414 149000
rect 370794 146000 371414 149000
rect 379794 146000 380414 149000
rect 388794 146000 389414 149000
rect 397794 146000 398414 149000
rect 406794 146000 407414 149000
rect 415794 146000 416414 149000
rect 424794 146000 425414 149000
rect 433794 146000 434414 149000
rect 442794 146000 443414 149000
rect 451794 146000 452414 149000
rect 460794 146000 461414 149000
rect 469794 146000 470414 149000
rect 478794 146000 479414 149000
rect 487794 146000 488414 149000
rect 496794 146000 497414 149000
rect 505794 146000 506414 149000
rect 514794 146000 515414 149000
rect 523794 146000 524414 149000
rect 532794 146000 533414 149000
rect 541794 146000 542414 149000
rect 550794 146000 551414 149000
rect 19794 119000 20414 122000
rect 28794 119000 29414 122000
rect 37794 119000 38414 122000
rect 46794 119000 47414 122000
rect 55794 119000 56414 122000
rect 64794 119000 65414 122000
rect 73794 119000 74414 122000
rect 82794 119000 83414 122000
rect 91794 119000 92414 122000
rect 100794 119000 101414 122000
rect 109794 119000 110414 122000
rect 118794 119000 119414 122000
rect 127794 119000 128414 122000
rect 136794 119000 137414 122000
rect 145794 119000 146414 122000
rect 154794 119000 155414 122000
rect 163794 119000 164414 122000
rect 172794 119000 173414 122000
rect 181794 119000 182414 122000
rect 190794 119000 191414 122000
rect 199794 119000 200414 122000
rect 208794 119000 209414 122000
rect 217794 119000 218414 122000
rect 226794 119000 227414 122000
rect 235794 119000 236414 122000
rect 244794 119000 245414 122000
rect 253794 119000 254414 122000
rect 262794 119000 263414 122000
rect 271794 119000 272414 122000
rect 280794 119000 281414 122000
rect 289794 119000 290414 122000
rect 298794 119000 299414 122000
rect 307794 119000 308414 122000
rect 316794 119000 317414 122000
rect 325794 119000 326414 122000
rect 334794 119000 335414 122000
rect 343794 119000 344414 122000
rect 352794 119000 353414 122000
rect 361794 119000 362414 122000
rect 370794 119000 371414 122000
rect 379794 119000 380414 122000
rect 388794 119000 389414 122000
rect 397794 119000 398414 122000
rect 406794 119000 407414 122000
rect 415794 119000 416414 122000
rect 424794 119000 425414 122000
rect 433794 119000 434414 122000
rect 442794 119000 443414 122000
rect 451794 119000 452414 122000
rect 460794 119000 461414 122000
rect 469794 119000 470414 122000
rect 478794 119000 479414 122000
rect 487794 119000 488414 122000
rect 496794 119000 497414 122000
rect 505794 119000 506414 122000
rect 514794 119000 515414 122000
rect 523794 119000 524414 122000
rect 532794 119000 533414 122000
rect 541794 119000 542414 122000
rect 550794 119000 551414 122000
rect 19794 92000 20414 95000
rect 28794 92000 29414 95000
rect 37794 92000 38414 95000
rect 46794 92000 47414 95000
rect 55794 92000 56414 95000
rect 64794 92000 65414 95000
rect 73794 92000 74414 95000
rect 82794 92000 83414 95000
rect 91794 92000 92414 95000
rect 100794 92000 101414 95000
rect 109794 92000 110414 95000
rect 118794 92000 119414 95000
rect 127794 92000 128414 95000
rect 136794 92000 137414 95000
rect 145794 92000 146414 95000
rect 154794 92000 155414 95000
rect 163794 92000 164414 95000
rect 172794 92000 173414 95000
rect 181794 92000 182414 95000
rect 190794 92000 191414 95000
rect 199794 92000 200414 95000
rect 208794 92000 209414 95000
rect 217794 92000 218414 95000
rect 226794 92000 227414 95000
rect 235794 92000 236414 95000
rect 244794 92000 245414 95000
rect 253794 92000 254414 95000
rect 262794 92000 263414 95000
rect 271794 92000 272414 95000
rect 280794 92000 281414 95000
rect 289794 92000 290414 95000
rect 298794 92000 299414 95000
rect 307794 92000 308414 95000
rect 316794 92000 317414 95000
rect 325794 92000 326414 95000
rect 334794 92000 335414 95000
rect 343794 92000 344414 95000
rect 352794 92000 353414 95000
rect 361794 92000 362414 95000
rect 370794 92000 371414 95000
rect 379794 92000 380414 95000
rect 388794 92000 389414 95000
rect 397794 92000 398414 95000
rect 406794 92000 407414 95000
rect 415794 92000 416414 95000
rect 424794 92000 425414 95000
rect 433794 92000 434414 95000
rect 442794 92000 443414 95000
rect 451794 92000 452414 95000
rect 460794 92000 461414 95000
rect 469794 92000 470414 95000
rect 478794 92000 479414 95000
rect 487794 92000 488414 95000
rect 496794 92000 497414 95000
rect 505794 92000 506414 95000
rect 514794 92000 515414 95000
rect 523794 92000 524414 95000
rect 532794 92000 533414 95000
rect 541794 92000 542414 95000
rect 550794 92000 551414 95000
rect 19794 65000 20414 68000
rect 28794 65000 29414 68000
rect 37794 65000 38414 68000
rect 46794 65000 47414 68000
rect 55794 65000 56414 68000
rect 64794 65000 65414 68000
rect 73794 65000 74414 68000
rect 82794 65000 83414 68000
rect 91794 65000 92414 68000
rect 100794 65000 101414 68000
rect 109794 65000 110414 68000
rect 118794 65000 119414 68000
rect 127794 65000 128414 68000
rect 136794 65000 137414 68000
rect 145794 65000 146414 68000
rect 154794 65000 155414 68000
rect 163794 65000 164414 68000
rect 172794 65000 173414 68000
rect 181794 65000 182414 68000
rect 190794 65000 191414 68000
rect 199794 65000 200414 68000
rect 208794 65000 209414 68000
rect 217794 65000 218414 68000
rect 226794 65000 227414 68000
rect 235794 65000 236414 68000
rect 244794 65000 245414 68000
rect 253794 65000 254414 68000
rect 262794 65000 263414 68000
rect 271794 65000 272414 68000
rect 280794 65000 281414 68000
rect 289794 65000 290414 68000
rect 298794 65000 299414 68000
rect 307794 65000 308414 68000
rect 316794 65000 317414 68000
rect 325794 65000 326414 68000
rect 334794 65000 335414 68000
rect 343794 65000 344414 68000
rect 352794 65000 353414 68000
rect 361794 65000 362414 68000
rect 370794 65000 371414 68000
rect 379794 65000 380414 68000
rect 388794 65000 389414 68000
rect 397794 65000 398414 68000
rect 406794 65000 407414 68000
rect 415794 65000 416414 68000
rect 424794 65000 425414 68000
rect 433794 65000 434414 68000
rect 442794 65000 443414 68000
rect 451794 65000 452414 68000
rect 460794 65000 461414 68000
rect 469794 65000 470414 68000
rect 478794 65000 479414 68000
rect 487794 65000 488414 68000
rect 496794 65000 497414 68000
rect 505794 65000 506414 68000
rect 514794 65000 515414 68000
rect 523794 65000 524414 68000
rect 532794 65000 533414 68000
rect 541794 65000 542414 68000
rect 550794 65000 551414 68000
rect 19794 38000 20414 41000
rect 28794 38000 29414 41000
rect 37794 38000 38414 41000
rect 46794 38000 47414 41000
rect 55794 38000 56414 41000
rect 19794 -1894 20414 14000
rect 28794 -1894 29414 14000
rect 37794 -1894 38414 14000
rect 46794 -1894 47414 14000
rect 55794 -1894 56414 14000
rect 64794 -1894 65414 41000
rect 73794 38000 74414 41000
rect 82794 38000 83414 41000
rect 91794 38000 92414 41000
rect 100794 38000 101414 41000
rect 109794 38000 110414 41000
rect 118794 38000 119414 41000
rect 127794 38000 128414 41000
rect 136794 38000 137414 41000
rect 145794 38000 146414 41000
rect 154794 38000 155414 41000
rect 163794 38000 164414 41000
rect 172794 38000 173414 41000
rect 181794 38000 182414 41000
rect 190794 38000 191414 41000
rect 199794 38000 200414 41000
rect 208794 38000 209414 41000
rect 217794 38000 218414 41000
rect 226794 38000 227414 41000
rect 235794 38000 236414 41000
rect 244794 38000 245414 41000
rect 253794 38000 254414 41000
rect 262794 38000 263414 41000
rect 271794 38000 272414 41000
rect 280794 38000 281414 41000
rect 289794 38000 290414 41000
rect 298794 38000 299414 41000
rect 307794 38000 308414 41000
rect 316794 38000 317414 41000
rect 325794 38000 326414 41000
rect 334794 38000 335414 41000
rect 343794 38000 344414 41000
rect 352794 38000 353414 41000
rect 361794 38000 362414 41000
rect 370794 38000 371414 41000
rect 379794 38000 380414 41000
rect 388794 38000 389414 41000
rect 397794 38000 398414 41000
rect 406794 38000 407414 41000
rect 415794 38000 416414 41000
rect 424794 38000 425414 41000
rect 433794 38000 434414 41000
rect 442794 38000 443414 41000
rect 451794 38000 452414 41000
rect 460794 38000 461414 41000
rect 469794 38000 470414 41000
rect 478794 38000 479414 41000
rect 487794 38000 488414 41000
rect 496794 38000 497414 41000
rect 505794 38000 506414 41000
rect 514794 38000 515414 41000
rect 523794 38000 524414 41000
rect 532794 38000 533414 41000
rect 541794 38000 542414 41000
rect 550794 38000 551414 41000
rect 73794 -1894 74414 14000
rect 82794 -1894 83414 14000
rect 91794 -1894 92414 14000
rect 100794 -1894 101414 14000
rect 109794 -1894 110414 14000
rect 118794 -1894 119414 14000
rect 127794 -1894 128414 14000
rect 136794 -1894 137414 14000
rect 145794 -1894 146414 14000
rect 154794 -1894 155414 14000
rect 163794 -1894 164414 14000
rect 172794 -1894 173414 14000
rect 181794 -1894 182414 14000
rect 190794 -1894 191414 14000
rect 199794 -1894 200414 14000
rect 208794 -1894 209414 14000
rect 217794 -1894 218414 14000
rect 226794 -1894 227414 14000
rect 235794 -1894 236414 14000
rect 244794 -1894 245414 14000
rect 253794 -1894 254414 14000
rect 262794 -1894 263414 14000
rect 271794 -1894 272414 14000
rect 280794 -1894 281414 14000
rect 289794 -1894 290414 14000
rect 298794 -1894 299414 14000
rect 307794 -1894 308414 14000
rect 316794 -1894 317414 14000
rect 325794 -1894 326414 14000
rect 334794 -1894 335414 14000
rect 343794 -1894 344414 14000
rect 352794 -1894 353414 14000
rect 361794 -1894 362414 14000
rect 370794 -1894 371414 14000
rect 379794 -1894 380414 14000
rect 388794 -1894 389414 14000
rect 397794 -1894 398414 14000
rect 406794 -1894 407414 14000
rect 415794 -1894 416414 14000
rect 424794 -1894 425414 14000
rect 433794 -1894 434414 14000
rect 442794 -1894 443414 14000
rect 451794 -1894 452414 14000
rect 460794 -1894 461414 14000
rect 469794 -1894 470414 14000
rect 478794 -1894 479414 14000
rect 487794 -1894 488414 14000
rect 496794 -1894 497414 14000
rect 505794 -1894 506414 14000
rect 514794 -1894 515414 14000
rect 523794 -1894 524414 14000
rect 532794 -1894 533414 14000
rect 541794 -1894 542414 14000
rect 550794 -1894 551414 14000
rect 559794 -1894 560414 705830
rect 568794 -1894 569414 705830
rect 577794 -1894 578414 705830
rect 585310 -934 585930 704870
rect 586270 -1894 586890 705830
<< obsm4 >>
rect 19910 662080 545091 681456
rect 20494 658920 28714 662080
rect 29494 658920 37714 662080
rect 38494 658920 46714 662080
rect 47494 658920 55714 662080
rect 56494 658920 64714 662080
rect 65494 658920 73714 662080
rect 74494 658920 82714 662080
rect 83494 658920 91714 662080
rect 92494 658920 100714 662080
rect 101494 658920 109714 662080
rect 110494 658920 118714 662080
rect 119494 658920 127714 662080
rect 128494 658920 136714 662080
rect 137494 658920 145714 662080
rect 146494 658920 154714 662080
rect 155494 658920 163714 662080
rect 164494 658920 172714 662080
rect 173494 658920 181714 662080
rect 182494 658920 190714 662080
rect 191494 658920 199714 662080
rect 200494 658920 208714 662080
rect 209494 658920 217714 662080
rect 218494 658920 226714 662080
rect 227494 658920 235714 662080
rect 236494 658920 244714 662080
rect 245494 658920 253714 662080
rect 254494 658920 262714 662080
rect 263494 658920 271714 662080
rect 272494 658920 280714 662080
rect 281494 658920 289714 662080
rect 290494 658920 298714 662080
rect 299494 658920 307714 662080
rect 308494 658920 316714 662080
rect 317494 658920 325714 662080
rect 326494 658920 334714 662080
rect 335494 658920 343714 662080
rect 344494 658920 352714 662080
rect 353494 658920 361714 662080
rect 362494 658920 370714 662080
rect 371494 658920 379714 662080
rect 380494 658920 388714 662080
rect 389494 658920 397714 662080
rect 398494 658920 406714 662080
rect 407494 658920 415714 662080
rect 416494 658920 424714 662080
rect 425494 658920 433714 662080
rect 434494 658920 442714 662080
rect 443494 658920 451714 662080
rect 452494 658920 460714 662080
rect 461494 658920 469714 662080
rect 470494 658920 478714 662080
rect 479494 658920 487714 662080
rect 488494 658920 496714 662080
rect 497494 658920 505714 662080
rect 506494 658920 514714 662080
rect 515494 658920 523714 662080
rect 524494 658920 532714 662080
rect 533494 658920 541714 662080
rect 542494 658920 545091 662080
rect 19910 635080 545091 658920
rect 20494 631920 28714 635080
rect 29494 631920 37714 635080
rect 38494 631920 46714 635080
rect 47494 631920 55714 635080
rect 56494 631920 64714 635080
rect 65494 631920 73714 635080
rect 74494 631920 82714 635080
rect 83494 631920 91714 635080
rect 92494 631920 100714 635080
rect 101494 631920 109714 635080
rect 110494 631920 118714 635080
rect 119494 631920 127714 635080
rect 128494 631920 136714 635080
rect 137494 631920 145714 635080
rect 146494 631920 154714 635080
rect 155494 631920 163714 635080
rect 164494 631920 172714 635080
rect 173494 631920 181714 635080
rect 182494 631920 190714 635080
rect 191494 631920 199714 635080
rect 200494 631920 208714 635080
rect 209494 631920 217714 635080
rect 218494 631920 226714 635080
rect 227494 631920 235714 635080
rect 236494 631920 244714 635080
rect 245494 631920 253714 635080
rect 254494 631920 262714 635080
rect 263494 631920 271714 635080
rect 272494 631920 280714 635080
rect 281494 631920 289714 635080
rect 290494 631920 298714 635080
rect 299494 631920 307714 635080
rect 308494 631920 316714 635080
rect 317494 631920 325714 635080
rect 326494 631920 334714 635080
rect 335494 631920 343714 635080
rect 344494 631920 352714 635080
rect 353494 631920 361714 635080
rect 362494 631920 370714 635080
rect 371494 631920 379714 635080
rect 380494 631920 388714 635080
rect 389494 631920 397714 635080
rect 398494 631920 406714 635080
rect 407494 631920 415714 635080
rect 416494 631920 424714 635080
rect 425494 631920 433714 635080
rect 434494 631920 442714 635080
rect 443494 631920 451714 635080
rect 452494 631920 460714 635080
rect 461494 631920 469714 635080
rect 470494 631920 478714 635080
rect 479494 631920 487714 635080
rect 488494 631920 496714 635080
rect 497494 631920 505714 635080
rect 506494 631920 514714 635080
rect 515494 631920 523714 635080
rect 524494 631920 532714 635080
rect 533494 631920 541714 635080
rect 542494 631920 545091 635080
rect 19910 608080 545091 631920
rect 20494 604920 28714 608080
rect 29494 604920 37714 608080
rect 38494 604920 46714 608080
rect 47494 604920 55714 608080
rect 56494 604920 64714 608080
rect 65494 604920 73714 608080
rect 74494 604920 82714 608080
rect 83494 604920 91714 608080
rect 92494 604920 100714 608080
rect 101494 604920 109714 608080
rect 110494 604920 118714 608080
rect 119494 604920 127714 608080
rect 128494 604920 136714 608080
rect 137494 604920 145714 608080
rect 146494 604920 154714 608080
rect 155494 604920 163714 608080
rect 164494 604920 172714 608080
rect 173494 604920 181714 608080
rect 182494 604920 190714 608080
rect 191494 604920 199714 608080
rect 200494 604920 208714 608080
rect 209494 604920 217714 608080
rect 218494 604920 226714 608080
rect 227494 604920 235714 608080
rect 236494 604920 244714 608080
rect 245494 604920 253714 608080
rect 254494 604920 262714 608080
rect 263494 604920 271714 608080
rect 272494 604920 280714 608080
rect 281494 604920 289714 608080
rect 290494 604920 298714 608080
rect 299494 604920 307714 608080
rect 308494 604920 316714 608080
rect 317494 604920 325714 608080
rect 326494 604920 334714 608080
rect 335494 604920 343714 608080
rect 344494 604920 352714 608080
rect 353494 604920 361714 608080
rect 362494 604920 370714 608080
rect 371494 604920 379714 608080
rect 380494 604920 388714 608080
rect 389494 604920 397714 608080
rect 398494 604920 406714 608080
rect 407494 604920 415714 608080
rect 416494 604920 424714 608080
rect 425494 604920 433714 608080
rect 434494 604920 442714 608080
rect 443494 604920 451714 608080
rect 452494 604920 460714 608080
rect 461494 604920 469714 608080
rect 470494 604920 478714 608080
rect 479494 604920 487714 608080
rect 488494 604920 496714 608080
rect 497494 604920 505714 608080
rect 506494 604920 514714 608080
rect 515494 604920 523714 608080
rect 524494 604920 532714 608080
rect 533494 604920 541714 608080
rect 542494 604920 545091 608080
rect 19910 581080 545091 604920
rect 20494 577920 28714 581080
rect 29494 577920 37714 581080
rect 38494 577920 46714 581080
rect 47494 577920 55714 581080
rect 56494 577920 64714 581080
rect 65494 577920 73714 581080
rect 74494 577920 82714 581080
rect 83494 577920 91714 581080
rect 92494 577920 100714 581080
rect 101494 577920 109714 581080
rect 110494 577920 118714 581080
rect 119494 577920 127714 581080
rect 128494 577920 136714 581080
rect 137494 577920 145714 581080
rect 146494 577920 154714 581080
rect 155494 577920 163714 581080
rect 164494 577920 172714 581080
rect 173494 577920 181714 581080
rect 182494 577920 190714 581080
rect 191494 577920 199714 581080
rect 200494 577920 208714 581080
rect 209494 577920 217714 581080
rect 218494 577920 226714 581080
rect 227494 577920 235714 581080
rect 236494 577920 244714 581080
rect 245494 577920 253714 581080
rect 254494 577920 262714 581080
rect 263494 577920 271714 581080
rect 272494 577920 280714 581080
rect 281494 577920 289714 581080
rect 290494 577920 298714 581080
rect 299494 577920 307714 581080
rect 308494 577920 316714 581080
rect 317494 577920 325714 581080
rect 326494 577920 334714 581080
rect 335494 577920 343714 581080
rect 344494 577920 352714 581080
rect 353494 577920 361714 581080
rect 362494 577920 370714 581080
rect 371494 577920 379714 581080
rect 380494 577920 388714 581080
rect 389494 577920 397714 581080
rect 398494 577920 406714 581080
rect 407494 577920 415714 581080
rect 416494 577920 424714 581080
rect 425494 577920 433714 581080
rect 434494 577920 442714 581080
rect 443494 577920 451714 581080
rect 452494 577920 460714 581080
rect 461494 577920 469714 581080
rect 470494 577920 478714 581080
rect 479494 577920 487714 581080
rect 488494 577920 496714 581080
rect 497494 577920 505714 581080
rect 506494 577920 514714 581080
rect 515494 577920 523714 581080
rect 524494 577920 532714 581080
rect 533494 577920 541714 581080
rect 542494 577920 545091 581080
rect 19910 554080 545091 577920
rect 20494 550920 28714 554080
rect 29494 550920 37714 554080
rect 38494 550920 46714 554080
rect 47494 550920 55714 554080
rect 56494 550920 64714 554080
rect 65494 550920 73714 554080
rect 74494 550920 82714 554080
rect 83494 550920 91714 554080
rect 92494 550920 100714 554080
rect 101494 550920 109714 554080
rect 110494 550920 118714 554080
rect 119494 550920 127714 554080
rect 128494 550920 136714 554080
rect 137494 550920 145714 554080
rect 146494 550920 154714 554080
rect 155494 550920 163714 554080
rect 164494 550920 172714 554080
rect 173494 550920 181714 554080
rect 182494 550920 190714 554080
rect 191494 550920 199714 554080
rect 200494 550920 208714 554080
rect 209494 550920 217714 554080
rect 218494 550920 226714 554080
rect 227494 550920 235714 554080
rect 236494 550920 244714 554080
rect 245494 550920 253714 554080
rect 254494 550920 262714 554080
rect 263494 550920 271714 554080
rect 272494 550920 280714 554080
rect 281494 550920 289714 554080
rect 290494 550920 298714 554080
rect 299494 550920 307714 554080
rect 308494 550920 316714 554080
rect 317494 550920 325714 554080
rect 326494 550920 334714 554080
rect 335494 550920 343714 554080
rect 344494 550920 352714 554080
rect 353494 550920 361714 554080
rect 362494 550920 370714 554080
rect 371494 550920 379714 554080
rect 380494 550920 388714 554080
rect 389494 550920 397714 554080
rect 398494 550920 406714 554080
rect 407494 550920 415714 554080
rect 416494 550920 424714 554080
rect 425494 550920 433714 554080
rect 434494 550920 442714 554080
rect 443494 550920 451714 554080
rect 452494 550920 460714 554080
rect 461494 550920 469714 554080
rect 470494 550920 478714 554080
rect 479494 550920 487714 554080
rect 488494 550920 496714 554080
rect 497494 550920 505714 554080
rect 506494 550920 514714 554080
rect 515494 550920 523714 554080
rect 524494 550920 532714 554080
rect 533494 550920 541714 554080
rect 542494 550920 545091 554080
rect 19910 527080 545091 550920
rect 20494 523920 28714 527080
rect 29494 523920 37714 527080
rect 38494 523920 46714 527080
rect 47494 523920 55714 527080
rect 56494 523920 64714 527080
rect 65494 523920 73714 527080
rect 74494 523920 82714 527080
rect 83494 523920 91714 527080
rect 92494 523920 100714 527080
rect 101494 523920 109714 527080
rect 110494 523920 118714 527080
rect 119494 523920 127714 527080
rect 128494 523920 136714 527080
rect 137494 523920 145714 527080
rect 146494 523920 154714 527080
rect 155494 523920 163714 527080
rect 164494 523920 172714 527080
rect 173494 523920 181714 527080
rect 182494 523920 190714 527080
rect 191494 523920 199714 527080
rect 200494 523920 208714 527080
rect 209494 523920 217714 527080
rect 218494 523920 226714 527080
rect 227494 523920 235714 527080
rect 236494 523920 244714 527080
rect 245494 523920 253714 527080
rect 254494 523920 262714 527080
rect 263494 523920 271714 527080
rect 272494 523920 280714 527080
rect 281494 523920 289714 527080
rect 290494 523920 298714 527080
rect 299494 523920 307714 527080
rect 308494 523920 316714 527080
rect 317494 523920 325714 527080
rect 326494 523920 334714 527080
rect 335494 523920 343714 527080
rect 344494 523920 352714 527080
rect 353494 523920 361714 527080
rect 362494 523920 370714 527080
rect 371494 523920 379714 527080
rect 380494 523920 388714 527080
rect 389494 523920 397714 527080
rect 398494 523920 406714 527080
rect 407494 523920 415714 527080
rect 416494 523920 424714 527080
rect 425494 523920 433714 527080
rect 434494 523920 442714 527080
rect 443494 523920 451714 527080
rect 452494 523920 460714 527080
rect 461494 523920 469714 527080
rect 470494 523920 478714 527080
rect 479494 523920 487714 527080
rect 488494 523920 496714 527080
rect 497494 523920 505714 527080
rect 506494 523920 514714 527080
rect 515494 523920 523714 527080
rect 524494 523920 532714 527080
rect 533494 523920 541714 527080
rect 542494 523920 545091 527080
rect 19910 500080 545091 523920
rect 20494 496920 28714 500080
rect 29494 496920 37714 500080
rect 38494 496920 46714 500080
rect 47494 496920 55714 500080
rect 56494 496920 64714 500080
rect 65494 496920 73714 500080
rect 74494 496920 82714 500080
rect 83494 496920 91714 500080
rect 92494 496920 100714 500080
rect 101494 496920 109714 500080
rect 110494 496920 118714 500080
rect 119494 496920 127714 500080
rect 128494 496920 136714 500080
rect 137494 496920 145714 500080
rect 146494 496920 154714 500080
rect 155494 496920 163714 500080
rect 164494 496920 172714 500080
rect 173494 496920 181714 500080
rect 182494 496920 190714 500080
rect 191494 496920 199714 500080
rect 200494 496920 208714 500080
rect 209494 496920 217714 500080
rect 218494 496920 226714 500080
rect 227494 496920 235714 500080
rect 236494 496920 244714 500080
rect 245494 496920 253714 500080
rect 254494 496920 262714 500080
rect 263494 496920 271714 500080
rect 272494 496920 280714 500080
rect 281494 496920 289714 500080
rect 290494 496920 298714 500080
rect 299494 496920 307714 500080
rect 308494 496920 316714 500080
rect 317494 496920 325714 500080
rect 326494 496920 334714 500080
rect 335494 496920 343714 500080
rect 344494 496920 352714 500080
rect 353494 496920 361714 500080
rect 362494 496920 370714 500080
rect 371494 496920 379714 500080
rect 380494 496920 388714 500080
rect 389494 496920 397714 500080
rect 398494 496920 406714 500080
rect 407494 496920 415714 500080
rect 416494 496920 424714 500080
rect 425494 496920 433714 500080
rect 434494 496920 442714 500080
rect 443494 496920 451714 500080
rect 452494 496920 460714 500080
rect 461494 496920 469714 500080
rect 470494 496920 478714 500080
rect 479494 496920 487714 500080
rect 488494 496920 496714 500080
rect 497494 496920 505714 500080
rect 506494 496920 514714 500080
rect 515494 496920 523714 500080
rect 524494 496920 532714 500080
rect 533494 496920 541714 500080
rect 542494 496920 545091 500080
rect 19910 473080 545091 496920
rect 20494 469920 28714 473080
rect 29494 469920 37714 473080
rect 38494 469920 46714 473080
rect 47494 469920 55714 473080
rect 56494 469920 64714 473080
rect 65494 469920 73714 473080
rect 74494 469920 82714 473080
rect 83494 469920 91714 473080
rect 92494 469920 100714 473080
rect 101494 469920 109714 473080
rect 110494 469920 118714 473080
rect 119494 469920 127714 473080
rect 128494 469920 136714 473080
rect 137494 469920 145714 473080
rect 146494 469920 154714 473080
rect 155494 469920 163714 473080
rect 164494 469920 172714 473080
rect 173494 469920 181714 473080
rect 182494 469920 190714 473080
rect 191494 469920 199714 473080
rect 200494 469920 208714 473080
rect 209494 469920 217714 473080
rect 218494 469920 226714 473080
rect 227494 469920 235714 473080
rect 236494 469920 244714 473080
rect 245494 469920 253714 473080
rect 254494 469920 262714 473080
rect 263494 469920 271714 473080
rect 272494 469920 280714 473080
rect 281494 469920 289714 473080
rect 290494 469920 298714 473080
rect 299494 469920 307714 473080
rect 308494 469920 316714 473080
rect 317494 469920 325714 473080
rect 326494 469920 334714 473080
rect 335494 469920 343714 473080
rect 344494 469920 352714 473080
rect 353494 469920 361714 473080
rect 362494 469920 370714 473080
rect 371494 469920 379714 473080
rect 380494 469920 388714 473080
rect 389494 469920 397714 473080
rect 398494 469920 406714 473080
rect 407494 469920 415714 473080
rect 416494 469920 424714 473080
rect 425494 469920 433714 473080
rect 434494 469920 442714 473080
rect 443494 469920 451714 473080
rect 452494 469920 460714 473080
rect 461494 469920 469714 473080
rect 470494 469920 478714 473080
rect 479494 469920 487714 473080
rect 488494 469920 496714 473080
rect 497494 469920 505714 473080
rect 506494 469920 514714 473080
rect 515494 469920 523714 473080
rect 524494 469920 532714 473080
rect 533494 469920 541714 473080
rect 542494 469920 545091 473080
rect 19910 446080 545091 469920
rect 20494 442920 28714 446080
rect 29494 442920 37714 446080
rect 38494 442920 46714 446080
rect 47494 442920 55714 446080
rect 56494 442920 64714 446080
rect 65494 442920 73714 446080
rect 74494 442920 82714 446080
rect 83494 442920 91714 446080
rect 92494 442920 100714 446080
rect 101494 442920 109714 446080
rect 110494 442920 118714 446080
rect 119494 442920 127714 446080
rect 128494 442920 136714 446080
rect 137494 442920 145714 446080
rect 146494 442920 154714 446080
rect 155494 442920 163714 446080
rect 164494 442920 172714 446080
rect 173494 442920 181714 446080
rect 182494 442920 190714 446080
rect 191494 442920 199714 446080
rect 200494 442920 208714 446080
rect 209494 442920 217714 446080
rect 218494 442920 226714 446080
rect 227494 442920 235714 446080
rect 236494 442920 244714 446080
rect 245494 442920 253714 446080
rect 254494 442920 262714 446080
rect 263494 442920 271714 446080
rect 272494 442920 280714 446080
rect 281494 442920 289714 446080
rect 290494 442920 298714 446080
rect 299494 442920 307714 446080
rect 308494 442920 316714 446080
rect 317494 442920 325714 446080
rect 326494 442920 334714 446080
rect 335494 442920 343714 446080
rect 344494 442920 352714 446080
rect 353494 442920 361714 446080
rect 362494 442920 370714 446080
rect 371494 442920 379714 446080
rect 380494 442920 388714 446080
rect 389494 442920 397714 446080
rect 398494 442920 406714 446080
rect 407494 442920 415714 446080
rect 416494 442920 424714 446080
rect 425494 442920 433714 446080
rect 434494 442920 442714 446080
rect 443494 442920 451714 446080
rect 452494 442920 460714 446080
rect 461494 442920 469714 446080
rect 470494 442920 478714 446080
rect 479494 442920 487714 446080
rect 488494 442920 496714 446080
rect 497494 442920 505714 446080
rect 506494 442920 514714 446080
rect 515494 442920 523714 446080
rect 524494 442920 532714 446080
rect 533494 442920 541714 446080
rect 542494 442920 545091 446080
rect 19910 419080 545091 442920
rect 20494 415920 28714 419080
rect 29494 415920 37714 419080
rect 38494 415920 46714 419080
rect 47494 415920 55714 419080
rect 56494 415920 64714 419080
rect 65494 415920 73714 419080
rect 74494 415920 82714 419080
rect 83494 415920 91714 419080
rect 92494 415920 100714 419080
rect 101494 415920 109714 419080
rect 110494 415920 118714 419080
rect 119494 415920 127714 419080
rect 128494 415920 136714 419080
rect 137494 415920 145714 419080
rect 146494 415920 154714 419080
rect 155494 415920 163714 419080
rect 164494 415920 172714 419080
rect 173494 415920 181714 419080
rect 182494 415920 190714 419080
rect 191494 415920 199714 419080
rect 200494 415920 208714 419080
rect 209494 415920 217714 419080
rect 218494 415920 226714 419080
rect 227494 415920 235714 419080
rect 236494 415920 244714 419080
rect 245494 415920 253714 419080
rect 254494 415920 262714 419080
rect 263494 415920 271714 419080
rect 272494 415920 280714 419080
rect 281494 415920 289714 419080
rect 290494 415920 298714 419080
rect 299494 415920 307714 419080
rect 308494 415920 316714 419080
rect 317494 415920 325714 419080
rect 326494 415920 334714 419080
rect 335494 415920 343714 419080
rect 344494 415920 352714 419080
rect 353494 415920 361714 419080
rect 362494 415920 370714 419080
rect 371494 415920 379714 419080
rect 380494 415920 388714 419080
rect 389494 415920 397714 419080
rect 398494 415920 406714 419080
rect 407494 415920 415714 419080
rect 416494 415920 424714 419080
rect 425494 415920 433714 419080
rect 434494 415920 442714 419080
rect 443494 415920 451714 419080
rect 452494 415920 460714 419080
rect 461494 415920 469714 419080
rect 470494 415920 478714 419080
rect 479494 415920 487714 419080
rect 488494 415920 496714 419080
rect 497494 415920 505714 419080
rect 506494 415920 514714 419080
rect 515494 415920 523714 419080
rect 524494 415920 532714 419080
rect 533494 415920 541714 419080
rect 542494 415920 545091 419080
rect 19910 392080 545091 415920
rect 20494 388920 28714 392080
rect 29494 388920 37714 392080
rect 38494 388920 46714 392080
rect 47494 388920 55714 392080
rect 56494 388920 64714 392080
rect 65494 388920 73714 392080
rect 74494 388920 82714 392080
rect 83494 388920 91714 392080
rect 92494 388920 100714 392080
rect 101494 388920 109714 392080
rect 110494 388920 118714 392080
rect 119494 388920 127714 392080
rect 128494 388920 136714 392080
rect 137494 388920 145714 392080
rect 146494 388920 154714 392080
rect 155494 388920 163714 392080
rect 164494 388920 172714 392080
rect 173494 388920 181714 392080
rect 182494 388920 190714 392080
rect 191494 388920 199714 392080
rect 200494 388920 208714 392080
rect 209494 388920 217714 392080
rect 218494 388920 226714 392080
rect 227494 388920 235714 392080
rect 236494 388920 244714 392080
rect 245494 388920 253714 392080
rect 254494 388920 262714 392080
rect 263494 388920 271714 392080
rect 272494 388920 280714 392080
rect 281494 388920 289714 392080
rect 290494 388920 298714 392080
rect 299494 388920 307714 392080
rect 308494 388920 316714 392080
rect 317494 388920 325714 392080
rect 326494 388920 334714 392080
rect 335494 388920 343714 392080
rect 344494 388920 352714 392080
rect 353494 388920 361714 392080
rect 362494 388920 370714 392080
rect 371494 388920 379714 392080
rect 380494 388920 388714 392080
rect 389494 388920 397714 392080
rect 398494 388920 406714 392080
rect 407494 388920 415714 392080
rect 416494 388920 424714 392080
rect 425494 388920 433714 392080
rect 434494 388920 442714 392080
rect 443494 388920 451714 392080
rect 452494 388920 460714 392080
rect 461494 388920 469714 392080
rect 470494 388920 478714 392080
rect 479494 388920 487714 392080
rect 488494 388920 496714 392080
rect 497494 388920 505714 392080
rect 506494 388920 514714 392080
rect 515494 388920 523714 392080
rect 524494 388920 532714 392080
rect 533494 388920 541714 392080
rect 542494 388920 545091 392080
rect 19910 365080 545091 388920
rect 20494 361920 28714 365080
rect 29494 361920 37714 365080
rect 38494 361920 46714 365080
rect 47494 361920 55714 365080
rect 56494 361920 64714 365080
rect 65494 361920 73714 365080
rect 74494 361920 82714 365080
rect 83494 361920 91714 365080
rect 92494 361920 100714 365080
rect 101494 361920 109714 365080
rect 110494 361920 118714 365080
rect 119494 361920 127714 365080
rect 128494 361920 136714 365080
rect 137494 361920 145714 365080
rect 146494 361920 154714 365080
rect 155494 361920 163714 365080
rect 164494 361920 172714 365080
rect 173494 361920 181714 365080
rect 182494 361920 190714 365080
rect 191494 361920 199714 365080
rect 200494 361920 208714 365080
rect 209494 361920 217714 365080
rect 218494 361920 226714 365080
rect 227494 361920 235714 365080
rect 236494 361920 244714 365080
rect 245494 361920 253714 365080
rect 254494 361920 262714 365080
rect 263494 361920 271714 365080
rect 272494 361920 280714 365080
rect 281494 361920 289714 365080
rect 290494 361920 298714 365080
rect 299494 361920 307714 365080
rect 308494 361920 316714 365080
rect 317494 361920 325714 365080
rect 326494 361920 334714 365080
rect 335494 361920 343714 365080
rect 344494 361920 352714 365080
rect 353494 361920 361714 365080
rect 362494 361920 370714 365080
rect 371494 361920 379714 365080
rect 380494 361920 388714 365080
rect 389494 361920 397714 365080
rect 398494 361920 406714 365080
rect 407494 361920 415714 365080
rect 416494 361920 424714 365080
rect 425494 361920 433714 365080
rect 434494 361920 442714 365080
rect 443494 361920 451714 365080
rect 452494 361920 460714 365080
rect 461494 361920 469714 365080
rect 470494 361920 478714 365080
rect 479494 361920 487714 365080
rect 488494 361920 496714 365080
rect 497494 361920 505714 365080
rect 506494 361920 514714 365080
rect 515494 361920 523714 365080
rect 524494 361920 532714 365080
rect 533494 361920 541714 365080
rect 542494 361920 545091 365080
rect 19910 338080 545091 361920
rect 20494 334920 28714 338080
rect 29494 334920 37714 338080
rect 38494 334920 46714 338080
rect 47494 334920 55714 338080
rect 56494 334920 64714 338080
rect 65494 334920 73714 338080
rect 74494 334920 82714 338080
rect 83494 334920 91714 338080
rect 92494 334920 100714 338080
rect 101494 334920 109714 338080
rect 110494 334920 118714 338080
rect 119494 334920 127714 338080
rect 128494 334920 136714 338080
rect 137494 334920 145714 338080
rect 146494 334920 154714 338080
rect 155494 334920 163714 338080
rect 164494 334920 172714 338080
rect 173494 334920 181714 338080
rect 182494 334920 190714 338080
rect 191494 334920 199714 338080
rect 200494 334920 208714 338080
rect 209494 334920 217714 338080
rect 218494 334920 226714 338080
rect 227494 334920 235714 338080
rect 236494 334920 244714 338080
rect 245494 334920 253714 338080
rect 254494 334920 262714 338080
rect 263494 334920 271714 338080
rect 272494 334920 280714 338080
rect 281494 334920 289714 338080
rect 290494 334920 298714 338080
rect 299494 334920 307714 338080
rect 308494 334920 316714 338080
rect 317494 334920 325714 338080
rect 326494 334920 334714 338080
rect 335494 334920 343714 338080
rect 344494 334920 352714 338080
rect 353494 334920 361714 338080
rect 362494 334920 370714 338080
rect 371494 334920 379714 338080
rect 380494 334920 388714 338080
rect 389494 334920 397714 338080
rect 398494 334920 406714 338080
rect 407494 334920 415714 338080
rect 416494 334920 424714 338080
rect 425494 334920 433714 338080
rect 434494 334920 442714 338080
rect 443494 334920 451714 338080
rect 452494 334920 460714 338080
rect 461494 334920 469714 338080
rect 470494 334920 478714 338080
rect 479494 334920 487714 338080
rect 488494 334920 496714 338080
rect 497494 334920 505714 338080
rect 506494 334920 514714 338080
rect 515494 334920 523714 338080
rect 524494 334920 532714 338080
rect 533494 334920 541714 338080
rect 542494 334920 545091 338080
rect 19910 311080 545091 334920
rect 20494 307920 28714 311080
rect 29494 307920 37714 311080
rect 38494 307920 46714 311080
rect 47494 307920 55714 311080
rect 56494 307920 64714 311080
rect 65494 307920 73714 311080
rect 74494 307920 82714 311080
rect 83494 307920 91714 311080
rect 92494 307920 100714 311080
rect 101494 307920 109714 311080
rect 110494 307920 118714 311080
rect 119494 307920 127714 311080
rect 128494 307920 136714 311080
rect 137494 307920 145714 311080
rect 146494 307920 154714 311080
rect 155494 307920 163714 311080
rect 164494 307920 172714 311080
rect 173494 307920 181714 311080
rect 182494 307920 190714 311080
rect 191494 307920 199714 311080
rect 200494 307920 208714 311080
rect 209494 307920 217714 311080
rect 218494 307920 226714 311080
rect 227494 307920 235714 311080
rect 236494 307920 244714 311080
rect 245494 307920 253714 311080
rect 254494 307920 262714 311080
rect 263494 307920 271714 311080
rect 272494 307920 280714 311080
rect 281494 307920 289714 311080
rect 290494 307920 298714 311080
rect 299494 307920 307714 311080
rect 308494 307920 316714 311080
rect 317494 307920 325714 311080
rect 326494 307920 334714 311080
rect 335494 307920 343714 311080
rect 344494 307920 352714 311080
rect 353494 307920 361714 311080
rect 362494 307920 370714 311080
rect 371494 307920 379714 311080
rect 380494 307920 388714 311080
rect 389494 307920 397714 311080
rect 398494 307920 406714 311080
rect 407494 307920 415714 311080
rect 416494 307920 424714 311080
rect 425494 307920 433714 311080
rect 434494 307920 442714 311080
rect 443494 307920 451714 311080
rect 452494 307920 460714 311080
rect 461494 307920 469714 311080
rect 470494 307920 478714 311080
rect 479494 307920 487714 311080
rect 488494 307920 496714 311080
rect 497494 307920 505714 311080
rect 506494 307920 514714 311080
rect 515494 307920 523714 311080
rect 524494 307920 532714 311080
rect 533494 307920 541714 311080
rect 542494 307920 545091 311080
rect 19910 284080 545091 307920
rect 20494 280920 28714 284080
rect 29494 280920 37714 284080
rect 38494 280920 46714 284080
rect 47494 280920 55714 284080
rect 56494 280920 64714 284080
rect 65494 280920 73714 284080
rect 74494 280920 82714 284080
rect 83494 280920 91714 284080
rect 92494 280920 100714 284080
rect 101494 280920 109714 284080
rect 110494 280920 118714 284080
rect 119494 280920 127714 284080
rect 128494 280920 136714 284080
rect 137494 280920 145714 284080
rect 146494 280920 154714 284080
rect 155494 280920 163714 284080
rect 164494 280920 172714 284080
rect 173494 280920 181714 284080
rect 182494 280920 190714 284080
rect 191494 280920 199714 284080
rect 200494 280920 208714 284080
rect 209494 280920 217714 284080
rect 218494 280920 226714 284080
rect 227494 280920 235714 284080
rect 236494 280920 244714 284080
rect 245494 280920 253714 284080
rect 254494 280920 262714 284080
rect 263494 280920 271714 284080
rect 272494 280920 280714 284080
rect 281494 280920 289714 284080
rect 290494 280920 298714 284080
rect 299494 280920 307714 284080
rect 308494 280920 316714 284080
rect 317494 280920 325714 284080
rect 326494 280920 334714 284080
rect 335494 280920 343714 284080
rect 344494 280920 352714 284080
rect 353494 280920 361714 284080
rect 362494 280920 370714 284080
rect 371494 280920 379714 284080
rect 380494 280920 388714 284080
rect 389494 280920 397714 284080
rect 398494 280920 406714 284080
rect 407494 280920 415714 284080
rect 416494 280920 424714 284080
rect 425494 280920 433714 284080
rect 434494 280920 442714 284080
rect 443494 280920 451714 284080
rect 452494 280920 460714 284080
rect 461494 280920 469714 284080
rect 470494 280920 478714 284080
rect 479494 280920 487714 284080
rect 488494 280920 496714 284080
rect 497494 280920 505714 284080
rect 506494 280920 514714 284080
rect 515494 280920 523714 284080
rect 524494 280920 532714 284080
rect 533494 280920 541714 284080
rect 542494 280920 545091 284080
rect 19910 257080 545091 280920
rect 20494 253920 28714 257080
rect 29494 253920 37714 257080
rect 38494 253920 46714 257080
rect 47494 253920 55714 257080
rect 56494 253920 64714 257080
rect 65494 253920 73714 257080
rect 74494 253920 82714 257080
rect 83494 253920 91714 257080
rect 92494 253920 100714 257080
rect 101494 253920 109714 257080
rect 110494 253920 118714 257080
rect 119494 253920 127714 257080
rect 128494 253920 136714 257080
rect 137494 253920 145714 257080
rect 146494 253920 154714 257080
rect 155494 253920 163714 257080
rect 164494 253920 172714 257080
rect 173494 253920 181714 257080
rect 182494 253920 190714 257080
rect 191494 253920 199714 257080
rect 200494 253920 208714 257080
rect 209494 253920 217714 257080
rect 218494 253920 226714 257080
rect 227494 253920 235714 257080
rect 236494 253920 244714 257080
rect 245494 253920 253714 257080
rect 254494 253920 262714 257080
rect 263494 253920 271714 257080
rect 272494 253920 280714 257080
rect 281494 253920 289714 257080
rect 290494 253920 298714 257080
rect 299494 253920 307714 257080
rect 308494 253920 316714 257080
rect 317494 253920 325714 257080
rect 326494 253920 334714 257080
rect 335494 253920 343714 257080
rect 344494 253920 352714 257080
rect 353494 253920 361714 257080
rect 362494 253920 370714 257080
rect 371494 253920 379714 257080
rect 380494 253920 388714 257080
rect 389494 253920 397714 257080
rect 398494 253920 406714 257080
rect 407494 253920 415714 257080
rect 416494 253920 424714 257080
rect 425494 253920 433714 257080
rect 434494 253920 442714 257080
rect 443494 253920 451714 257080
rect 452494 253920 460714 257080
rect 461494 253920 469714 257080
rect 470494 253920 478714 257080
rect 479494 253920 487714 257080
rect 488494 253920 496714 257080
rect 497494 253920 505714 257080
rect 506494 253920 514714 257080
rect 515494 253920 523714 257080
rect 524494 253920 532714 257080
rect 533494 253920 541714 257080
rect 542494 253920 545091 257080
rect 19910 230080 545091 253920
rect 20494 226920 28714 230080
rect 29494 226920 37714 230080
rect 38494 226920 46714 230080
rect 47494 226920 55714 230080
rect 56494 226920 64714 230080
rect 65494 226920 73714 230080
rect 74494 226920 82714 230080
rect 83494 226920 91714 230080
rect 92494 226920 100714 230080
rect 101494 226920 109714 230080
rect 110494 226920 118714 230080
rect 119494 226920 127714 230080
rect 128494 226920 136714 230080
rect 137494 226920 145714 230080
rect 146494 226920 154714 230080
rect 155494 226920 163714 230080
rect 164494 226920 172714 230080
rect 173494 226920 181714 230080
rect 182494 226920 190714 230080
rect 191494 226920 199714 230080
rect 200494 226920 208714 230080
rect 209494 226920 217714 230080
rect 218494 226920 226714 230080
rect 227494 226920 235714 230080
rect 236494 226920 244714 230080
rect 245494 226920 253714 230080
rect 254494 226920 262714 230080
rect 263494 226920 271714 230080
rect 272494 226920 280714 230080
rect 281494 226920 289714 230080
rect 290494 226920 298714 230080
rect 299494 226920 307714 230080
rect 308494 226920 316714 230080
rect 317494 226920 325714 230080
rect 326494 226920 334714 230080
rect 335494 226920 343714 230080
rect 344494 226920 352714 230080
rect 353494 226920 361714 230080
rect 362494 226920 370714 230080
rect 371494 226920 379714 230080
rect 380494 226920 388714 230080
rect 389494 226920 397714 230080
rect 398494 226920 406714 230080
rect 407494 226920 415714 230080
rect 416494 226920 424714 230080
rect 425494 226920 433714 230080
rect 434494 226920 442714 230080
rect 443494 226920 451714 230080
rect 452494 226920 460714 230080
rect 461494 226920 469714 230080
rect 470494 226920 478714 230080
rect 479494 226920 487714 230080
rect 488494 226920 496714 230080
rect 497494 226920 505714 230080
rect 506494 226920 514714 230080
rect 515494 226920 523714 230080
rect 524494 226920 532714 230080
rect 533494 226920 541714 230080
rect 542494 226920 545091 230080
rect 19910 203080 545091 226920
rect 20494 199920 28714 203080
rect 29494 199920 37714 203080
rect 38494 199920 46714 203080
rect 47494 199920 55714 203080
rect 56494 199920 64714 203080
rect 65494 199920 73714 203080
rect 74494 199920 82714 203080
rect 83494 199920 91714 203080
rect 92494 199920 100714 203080
rect 101494 199920 109714 203080
rect 110494 199920 118714 203080
rect 119494 199920 127714 203080
rect 128494 199920 136714 203080
rect 137494 199920 145714 203080
rect 146494 199920 154714 203080
rect 155494 199920 163714 203080
rect 164494 199920 172714 203080
rect 173494 199920 181714 203080
rect 182494 199920 190714 203080
rect 191494 199920 199714 203080
rect 200494 199920 208714 203080
rect 209494 199920 217714 203080
rect 218494 199920 226714 203080
rect 227494 199920 235714 203080
rect 236494 199920 244714 203080
rect 245494 199920 253714 203080
rect 254494 199920 262714 203080
rect 263494 199920 271714 203080
rect 272494 199920 280714 203080
rect 281494 199920 289714 203080
rect 290494 199920 298714 203080
rect 299494 199920 307714 203080
rect 308494 199920 316714 203080
rect 317494 199920 325714 203080
rect 326494 199920 334714 203080
rect 335494 199920 343714 203080
rect 344494 199920 352714 203080
rect 353494 199920 361714 203080
rect 362494 199920 370714 203080
rect 371494 199920 379714 203080
rect 380494 199920 388714 203080
rect 389494 199920 397714 203080
rect 398494 199920 406714 203080
rect 407494 199920 415714 203080
rect 416494 199920 424714 203080
rect 425494 199920 433714 203080
rect 434494 199920 442714 203080
rect 443494 199920 451714 203080
rect 452494 199920 460714 203080
rect 461494 199920 469714 203080
rect 470494 199920 478714 203080
rect 479494 199920 487714 203080
rect 488494 199920 496714 203080
rect 497494 199920 505714 203080
rect 506494 199920 514714 203080
rect 515494 199920 523714 203080
rect 524494 199920 532714 203080
rect 533494 199920 541714 203080
rect 542494 199920 545091 203080
rect 19910 176080 545091 199920
rect 20494 172920 28714 176080
rect 29494 172920 37714 176080
rect 38494 172920 46714 176080
rect 47494 172920 55714 176080
rect 56494 172920 64714 176080
rect 65494 172920 73714 176080
rect 74494 172920 82714 176080
rect 83494 172920 91714 176080
rect 92494 172920 100714 176080
rect 101494 172920 109714 176080
rect 110494 172920 118714 176080
rect 119494 172920 127714 176080
rect 128494 172920 136714 176080
rect 137494 172920 145714 176080
rect 146494 172920 154714 176080
rect 155494 172920 163714 176080
rect 164494 172920 172714 176080
rect 173494 172920 181714 176080
rect 182494 172920 190714 176080
rect 191494 172920 199714 176080
rect 200494 172920 208714 176080
rect 209494 172920 217714 176080
rect 218494 172920 226714 176080
rect 227494 172920 235714 176080
rect 236494 172920 244714 176080
rect 245494 172920 253714 176080
rect 254494 172920 262714 176080
rect 263494 172920 271714 176080
rect 272494 172920 280714 176080
rect 281494 172920 289714 176080
rect 290494 172920 298714 176080
rect 299494 172920 307714 176080
rect 308494 172920 316714 176080
rect 317494 172920 325714 176080
rect 326494 172920 334714 176080
rect 335494 172920 343714 176080
rect 344494 172920 352714 176080
rect 353494 172920 361714 176080
rect 362494 172920 370714 176080
rect 371494 172920 379714 176080
rect 380494 172920 388714 176080
rect 389494 172920 397714 176080
rect 398494 172920 406714 176080
rect 407494 172920 415714 176080
rect 416494 172920 424714 176080
rect 425494 172920 433714 176080
rect 434494 172920 442714 176080
rect 443494 172920 451714 176080
rect 452494 172920 460714 176080
rect 461494 172920 469714 176080
rect 470494 172920 478714 176080
rect 479494 172920 487714 176080
rect 488494 172920 496714 176080
rect 497494 172920 505714 176080
rect 506494 172920 514714 176080
rect 515494 172920 523714 176080
rect 524494 172920 532714 176080
rect 533494 172920 541714 176080
rect 542494 172920 545091 176080
rect 19910 149080 545091 172920
rect 20494 145920 28714 149080
rect 29494 145920 37714 149080
rect 38494 145920 46714 149080
rect 47494 145920 55714 149080
rect 56494 145920 64714 149080
rect 65494 145920 73714 149080
rect 74494 145920 82714 149080
rect 83494 145920 91714 149080
rect 92494 145920 100714 149080
rect 101494 145920 109714 149080
rect 110494 145920 118714 149080
rect 119494 145920 127714 149080
rect 128494 145920 136714 149080
rect 137494 145920 145714 149080
rect 146494 145920 154714 149080
rect 155494 145920 163714 149080
rect 164494 145920 172714 149080
rect 173494 145920 181714 149080
rect 182494 145920 190714 149080
rect 191494 145920 199714 149080
rect 200494 145920 208714 149080
rect 209494 145920 217714 149080
rect 218494 145920 226714 149080
rect 227494 145920 235714 149080
rect 236494 145920 244714 149080
rect 245494 145920 253714 149080
rect 254494 145920 262714 149080
rect 263494 145920 271714 149080
rect 272494 145920 280714 149080
rect 281494 145920 289714 149080
rect 290494 145920 298714 149080
rect 299494 145920 307714 149080
rect 308494 145920 316714 149080
rect 317494 145920 325714 149080
rect 326494 145920 334714 149080
rect 335494 145920 343714 149080
rect 344494 145920 352714 149080
rect 353494 145920 361714 149080
rect 362494 145920 370714 149080
rect 371494 145920 379714 149080
rect 380494 145920 388714 149080
rect 389494 145920 397714 149080
rect 398494 145920 406714 149080
rect 407494 145920 415714 149080
rect 416494 145920 424714 149080
rect 425494 145920 433714 149080
rect 434494 145920 442714 149080
rect 443494 145920 451714 149080
rect 452494 145920 460714 149080
rect 461494 145920 469714 149080
rect 470494 145920 478714 149080
rect 479494 145920 487714 149080
rect 488494 145920 496714 149080
rect 497494 145920 505714 149080
rect 506494 145920 514714 149080
rect 515494 145920 523714 149080
rect 524494 145920 532714 149080
rect 533494 145920 541714 149080
rect 542494 145920 545091 149080
rect 19910 122080 545091 145920
rect 20494 118920 28714 122080
rect 29494 118920 37714 122080
rect 38494 118920 46714 122080
rect 47494 118920 55714 122080
rect 56494 118920 64714 122080
rect 65494 118920 73714 122080
rect 74494 118920 82714 122080
rect 83494 118920 91714 122080
rect 92494 118920 100714 122080
rect 101494 118920 109714 122080
rect 110494 118920 118714 122080
rect 119494 118920 127714 122080
rect 128494 118920 136714 122080
rect 137494 118920 145714 122080
rect 146494 118920 154714 122080
rect 155494 118920 163714 122080
rect 164494 118920 172714 122080
rect 173494 118920 181714 122080
rect 182494 118920 190714 122080
rect 191494 118920 199714 122080
rect 200494 118920 208714 122080
rect 209494 118920 217714 122080
rect 218494 118920 226714 122080
rect 227494 118920 235714 122080
rect 236494 118920 244714 122080
rect 245494 118920 253714 122080
rect 254494 118920 262714 122080
rect 263494 118920 271714 122080
rect 272494 118920 280714 122080
rect 281494 118920 289714 122080
rect 290494 118920 298714 122080
rect 299494 118920 307714 122080
rect 308494 118920 316714 122080
rect 317494 118920 325714 122080
rect 326494 118920 334714 122080
rect 335494 118920 343714 122080
rect 344494 118920 352714 122080
rect 353494 118920 361714 122080
rect 362494 118920 370714 122080
rect 371494 118920 379714 122080
rect 380494 118920 388714 122080
rect 389494 118920 397714 122080
rect 398494 118920 406714 122080
rect 407494 118920 415714 122080
rect 416494 118920 424714 122080
rect 425494 118920 433714 122080
rect 434494 118920 442714 122080
rect 443494 118920 451714 122080
rect 452494 118920 460714 122080
rect 461494 118920 469714 122080
rect 470494 118920 478714 122080
rect 479494 118920 487714 122080
rect 488494 118920 496714 122080
rect 497494 118920 505714 122080
rect 506494 118920 514714 122080
rect 515494 118920 523714 122080
rect 524494 118920 532714 122080
rect 533494 118920 541714 122080
rect 542494 118920 545091 122080
rect 19910 95080 545091 118920
rect 20494 91920 28714 95080
rect 29494 91920 37714 95080
rect 38494 91920 46714 95080
rect 47494 91920 55714 95080
rect 56494 91920 64714 95080
rect 65494 91920 73714 95080
rect 74494 91920 82714 95080
rect 83494 91920 91714 95080
rect 92494 91920 100714 95080
rect 101494 91920 109714 95080
rect 110494 91920 118714 95080
rect 119494 91920 127714 95080
rect 128494 91920 136714 95080
rect 137494 91920 145714 95080
rect 146494 91920 154714 95080
rect 155494 91920 163714 95080
rect 164494 91920 172714 95080
rect 173494 91920 181714 95080
rect 182494 91920 190714 95080
rect 191494 91920 199714 95080
rect 200494 91920 208714 95080
rect 209494 91920 217714 95080
rect 218494 91920 226714 95080
rect 227494 91920 235714 95080
rect 236494 91920 244714 95080
rect 245494 91920 253714 95080
rect 254494 91920 262714 95080
rect 263494 91920 271714 95080
rect 272494 91920 280714 95080
rect 281494 91920 289714 95080
rect 290494 91920 298714 95080
rect 299494 91920 307714 95080
rect 308494 91920 316714 95080
rect 317494 91920 325714 95080
rect 326494 91920 334714 95080
rect 335494 91920 343714 95080
rect 344494 91920 352714 95080
rect 353494 91920 361714 95080
rect 362494 91920 370714 95080
rect 371494 91920 379714 95080
rect 380494 91920 388714 95080
rect 389494 91920 397714 95080
rect 398494 91920 406714 95080
rect 407494 91920 415714 95080
rect 416494 91920 424714 95080
rect 425494 91920 433714 95080
rect 434494 91920 442714 95080
rect 443494 91920 451714 95080
rect 452494 91920 460714 95080
rect 461494 91920 469714 95080
rect 470494 91920 478714 95080
rect 479494 91920 487714 95080
rect 488494 91920 496714 95080
rect 497494 91920 505714 95080
rect 506494 91920 514714 95080
rect 515494 91920 523714 95080
rect 524494 91920 532714 95080
rect 533494 91920 541714 95080
rect 542494 91920 545091 95080
rect 19910 68080 545091 91920
rect 20494 64920 28714 68080
rect 29494 64920 37714 68080
rect 38494 64920 46714 68080
rect 47494 64920 55714 68080
rect 56494 64920 64714 68080
rect 65494 64920 73714 68080
rect 74494 64920 82714 68080
rect 83494 64920 91714 68080
rect 92494 64920 100714 68080
rect 101494 64920 109714 68080
rect 110494 64920 118714 68080
rect 119494 64920 127714 68080
rect 128494 64920 136714 68080
rect 137494 64920 145714 68080
rect 146494 64920 154714 68080
rect 155494 64920 163714 68080
rect 164494 64920 172714 68080
rect 173494 64920 181714 68080
rect 182494 64920 190714 68080
rect 191494 64920 199714 68080
rect 200494 64920 208714 68080
rect 209494 64920 217714 68080
rect 218494 64920 226714 68080
rect 227494 64920 235714 68080
rect 236494 64920 244714 68080
rect 245494 64920 253714 68080
rect 254494 64920 262714 68080
rect 263494 64920 271714 68080
rect 272494 64920 280714 68080
rect 281494 64920 289714 68080
rect 290494 64920 298714 68080
rect 299494 64920 307714 68080
rect 308494 64920 316714 68080
rect 317494 64920 325714 68080
rect 326494 64920 334714 68080
rect 335494 64920 343714 68080
rect 344494 64920 352714 68080
rect 353494 64920 361714 68080
rect 362494 64920 370714 68080
rect 371494 64920 379714 68080
rect 380494 64920 388714 68080
rect 389494 64920 397714 68080
rect 398494 64920 406714 68080
rect 407494 64920 415714 68080
rect 416494 64920 424714 68080
rect 425494 64920 433714 68080
rect 434494 64920 442714 68080
rect 443494 64920 451714 68080
rect 452494 64920 460714 68080
rect 461494 64920 469714 68080
rect 470494 64920 478714 68080
rect 479494 64920 487714 68080
rect 488494 64920 496714 68080
rect 497494 64920 505714 68080
rect 506494 64920 514714 68080
rect 515494 64920 523714 68080
rect 524494 64920 532714 68080
rect 533494 64920 541714 68080
rect 542494 64920 545091 68080
rect 19910 41080 545091 64920
rect 20494 37920 28714 41080
rect 29494 37920 37714 41080
rect 38494 37920 46714 41080
rect 47494 37920 55714 41080
rect 56494 37920 64714 41080
rect 19910 18128 64714 37920
rect 65494 37920 73714 41080
rect 74494 37920 82714 41080
rect 83494 37920 91714 41080
rect 92494 37920 100714 41080
rect 101494 37920 109714 41080
rect 110494 37920 118714 41080
rect 119494 37920 127714 41080
rect 128494 37920 136714 41080
rect 137494 37920 145714 41080
rect 146494 37920 154714 41080
rect 155494 37920 163714 41080
rect 164494 37920 172714 41080
rect 173494 37920 181714 41080
rect 182494 37920 190714 41080
rect 191494 37920 199714 41080
rect 200494 37920 208714 41080
rect 209494 37920 217714 41080
rect 218494 37920 226714 41080
rect 227494 37920 235714 41080
rect 236494 37920 244714 41080
rect 245494 37920 253714 41080
rect 254494 37920 262714 41080
rect 263494 37920 271714 41080
rect 272494 37920 280714 41080
rect 281494 37920 289714 41080
rect 290494 37920 298714 41080
rect 299494 37920 307714 41080
rect 308494 37920 316714 41080
rect 317494 37920 325714 41080
rect 326494 37920 334714 41080
rect 335494 37920 343714 41080
rect 344494 37920 352714 41080
rect 353494 37920 361714 41080
rect 362494 37920 370714 41080
rect 371494 37920 379714 41080
rect 380494 37920 388714 41080
rect 389494 37920 397714 41080
rect 398494 37920 406714 41080
rect 407494 37920 415714 41080
rect 416494 37920 424714 41080
rect 425494 37920 433714 41080
rect 434494 37920 442714 41080
rect 443494 37920 451714 41080
rect 452494 37920 460714 41080
rect 461494 37920 469714 41080
rect 470494 37920 478714 41080
rect 479494 37920 487714 41080
rect 488494 37920 496714 41080
rect 497494 37920 505714 41080
rect 506494 37920 514714 41080
rect 515494 37920 523714 41080
rect 524494 37920 532714 41080
rect 533494 37920 541714 41080
rect 542494 37920 545091 41080
rect 65494 18128 545091 37920
<< metal5 >>
rect -2966 705210 586890 705830
rect -2006 704250 585930 704870
rect -2966 695866 586890 696486
rect -2966 686866 586890 687486
rect -2966 677866 586890 678486
rect -2966 668866 586890 669486
rect 19794 660806 542414 661426
rect -2966 659866 586890 660486
rect -2966 650866 586890 651486
rect -2966 641866 586890 642486
rect 28794 633806 551414 634426
rect -2966 632866 586890 633486
rect -2966 623866 586890 624486
rect -2966 614866 586890 615486
rect 19794 606806 542414 607426
rect -2966 605866 586890 606486
rect -2966 596866 586890 597486
rect -2966 587866 586890 588486
rect 28794 579806 551414 580426
rect -2966 578866 586890 579486
rect -2966 569866 586890 570486
rect -2966 560866 586890 561486
rect 19794 552806 542414 553426
rect -2966 551866 586890 552486
rect -2966 542866 586890 543486
rect -2966 533866 586890 534486
rect 28794 525806 551414 526426
rect -2966 524866 586890 525486
rect -2966 515866 586890 516486
rect -2966 506866 586890 507486
rect 19794 498806 542414 499426
rect -2966 497866 586890 498486
rect -2966 488866 586890 489486
rect -2966 479866 586890 480486
rect 28794 471806 551414 472426
rect -2966 470866 586890 471486
rect -2966 461866 586890 462486
rect -2966 452866 586890 453486
rect 19794 444806 542414 445426
rect -2966 443866 586890 444486
rect -2966 434866 586890 435486
rect -2966 425866 586890 426486
rect 28794 417806 551414 418426
rect -2966 416866 586890 417486
rect -2966 407866 586890 408486
rect -2966 398866 586890 399486
rect 19794 390806 542414 391426
rect -2966 389866 586890 390486
rect -2966 380866 586890 381486
rect -2966 371866 586890 372486
rect 28794 363806 551414 364426
rect -2966 362866 586890 363486
rect -2966 353866 586890 354486
rect -2966 344866 586890 345486
rect 19794 336806 542414 337426
rect -2966 335866 586890 336486
rect -2966 326866 586890 327486
rect -2966 317866 586890 318486
rect 28794 309806 551414 310426
rect -2966 308866 586890 309486
rect -2966 299866 586890 300486
rect -2966 290866 586890 291486
rect 19794 282806 542414 283426
rect -2966 281866 586890 282486
rect -2966 272866 586890 273486
rect -2966 263866 586890 264486
rect 28794 255806 551414 256426
rect -2966 254866 586890 255486
rect -2966 245866 586890 246486
rect -2966 236866 586890 237486
rect 19794 228806 542414 229426
rect -2966 227866 586890 228486
rect -2966 218866 586890 219486
rect -2966 209866 586890 210486
rect 28794 201806 551414 202426
rect -2966 200866 586890 201486
rect -2966 191866 586890 192486
rect -2966 182866 586890 183486
rect 19794 174806 542414 175426
rect -2966 173866 586890 174486
rect -2966 164866 586890 165486
rect -2966 155866 586890 156486
rect 28794 147806 551414 148426
rect -2966 146866 586890 147486
rect -2966 137866 586890 138486
rect -2966 128866 586890 129486
rect 19794 120806 542414 121426
rect -2966 119866 586890 120486
rect -2966 110866 586890 111486
rect -2966 101866 586890 102486
rect 28794 93806 551414 94426
rect -2966 92866 586890 93486
rect -2966 83866 586890 84486
rect -2966 74866 586890 75486
rect 19794 66806 542414 67426
rect -2966 65866 586890 66486
rect -2966 56866 586890 57486
rect -2966 47866 586890 48486
rect 28794 39806 551414 40426
rect -2966 38866 586890 39486
rect -2966 29866 586890 30486
rect -2966 20866 586890 21486
rect -2966 11866 586890 12486
rect -2966 2866 586890 3486
rect -2006 -934 585930 -314
rect -2966 -1894 586890 -1274
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 46 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 47 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 48 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 49 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 50 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 51 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 53 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 54 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 55 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 56 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 57 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 58 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 59 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 60 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 122 nsew signal output
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 123 nsew signal output
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 124 nsew signal output
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 125 nsew signal output
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 126 nsew signal output
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 127 nsew signal output
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 129 nsew signal output
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 130 nsew signal output
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 131 nsew signal output
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 132 nsew signal output
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 133 nsew signal output
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 134 nsew signal output
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 135 nsew signal output
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 136 nsew signal output
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 528 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 531 nsew signal output
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 532 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 20866 586890 21486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 56866 586890 57486 6 vccd1
port 532 nsew power input
rlabel metal5 s 19794 66806 542414 67426 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 92866 586890 93486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 532 nsew power input
rlabel metal5 s 19794 120806 542414 121426 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 128866 586890 129486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 164866 586890 165486 6 vccd1
port 532 nsew power input
rlabel metal5 s 19794 174806 542414 175426 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 200866 586890 201486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 532 nsew power input
rlabel metal5 s 19794 228806 542414 229426 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 236866 586890 237486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 272866 586890 273486 6 vccd1
port 532 nsew power input
rlabel metal5 s 19794 282806 542414 283426 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 308866 586890 309486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 532 nsew power input
rlabel metal5 s 19794 336806 542414 337426 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 344866 586890 345486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 380866 586890 381486 6 vccd1
port 532 nsew power input
rlabel metal5 s 19794 390806 542414 391426 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 416866 586890 417486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 532 nsew power input
rlabel metal5 s 19794 444806 542414 445426 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 452866 586890 453486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 488866 586890 489486 6 vccd1
port 532 nsew power input
rlabel metal5 s 19794 498806 542414 499426 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 524866 586890 525486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 532 nsew power input
rlabel metal5 s 19794 552806 542414 553426 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 560866 586890 561486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 596866 586890 597486 6 vccd1
port 532 nsew power input
rlabel metal5 s 19794 606806 542414 607426 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 632866 586890 633486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 532 nsew power input
rlabel metal5 s 19794 660806 542414 661426 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 668866 586890 669486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 532 nsew power input
rlabel metal4 s 19794 -1894 20414 14000 6 vccd1
port 532 nsew power input
rlabel metal4 s 37794 -1894 38414 14000 6 vccd1
port 532 nsew power input
rlabel metal4 s 55794 -1894 56414 14000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 -1894 74414 14000 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 -1894 92414 14000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 -1894 110414 14000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 -1894 128414 14000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 -1894 146414 14000 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 -1894 164414 14000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 -1894 182414 14000 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 -1894 200414 14000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 -1894 218414 14000 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 -1894 236414 14000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 -1894 254414 14000 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 -1894 272414 14000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 -1894 290414 14000 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 -1894 308414 14000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 -1894 326414 14000 6 vccd1
port 532 nsew power input
rlabel metal4 s 343794 -1894 344414 14000 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 -1894 362414 14000 6 vccd1
port 532 nsew power input
rlabel metal4 s 379794 -1894 380414 14000 6 vccd1
port 532 nsew power input
rlabel metal4 s 397794 -1894 398414 14000 6 vccd1
port 532 nsew power input
rlabel metal4 s 415794 -1894 416414 14000 6 vccd1
port 532 nsew power input
rlabel metal4 s 433794 -1894 434414 14000 6 vccd1
port 532 nsew power input
rlabel metal4 s 451794 -1894 452414 14000 6 vccd1
port 532 nsew power input
rlabel metal4 s 469794 -1894 470414 14000 6 vccd1
port 532 nsew power input
rlabel metal4 s 487794 -1894 488414 14000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 -1894 506414 14000 6 vccd1
port 532 nsew power input
rlabel metal4 s 523794 -1894 524414 14000 6 vccd1
port 532 nsew power input
rlabel metal4 s 541794 -1894 542414 14000 6 vccd1
port 532 nsew power input
rlabel metal4 s 19794 38000 20414 41000 6 vccd1
port 532 nsew power input
rlabel metal4 s 37794 38000 38414 41000 6 vccd1
port 532 nsew power input
rlabel metal4 s 55794 38000 56414 41000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 38000 74414 41000 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 38000 92414 41000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 38000 110414 41000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 38000 128414 41000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 38000 146414 41000 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 38000 164414 41000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 38000 182414 41000 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 38000 200414 41000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 38000 218414 41000 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 38000 236414 41000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 38000 254414 41000 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 38000 272414 41000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 38000 290414 41000 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 38000 308414 41000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 38000 326414 41000 6 vccd1
port 532 nsew power input
rlabel metal4 s 343794 38000 344414 41000 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 38000 362414 41000 6 vccd1
port 532 nsew power input
rlabel metal4 s 379794 38000 380414 41000 6 vccd1
port 532 nsew power input
rlabel metal4 s 397794 38000 398414 41000 6 vccd1
port 532 nsew power input
rlabel metal4 s 415794 38000 416414 41000 6 vccd1
port 532 nsew power input
rlabel metal4 s 433794 38000 434414 41000 6 vccd1
port 532 nsew power input
rlabel metal4 s 451794 38000 452414 41000 6 vccd1
port 532 nsew power input
rlabel metal4 s 469794 38000 470414 41000 6 vccd1
port 532 nsew power input
rlabel metal4 s 487794 38000 488414 41000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 38000 506414 41000 6 vccd1
port 532 nsew power input
rlabel metal4 s 523794 38000 524414 41000 6 vccd1
port 532 nsew power input
rlabel metal4 s 541794 38000 542414 41000 6 vccd1
port 532 nsew power input
rlabel metal4 s 19794 65000 20414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 37794 65000 38414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 55794 65000 56414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 65000 74414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 65000 92414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 65000 110414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 65000 128414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 65000 146414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 65000 164414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 65000 182414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 65000 200414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 65000 218414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 65000 236414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 65000 254414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 65000 272414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 65000 290414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 65000 308414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 65000 326414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 343794 65000 344414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 65000 362414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 379794 65000 380414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 397794 65000 398414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 415794 65000 416414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 433794 65000 434414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 451794 65000 452414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 469794 65000 470414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 487794 65000 488414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 65000 506414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 523794 65000 524414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 541794 65000 542414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 19794 92000 20414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 37794 92000 38414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 55794 92000 56414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 92000 74414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 92000 92414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 92000 110414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 92000 128414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 92000 146414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 92000 164414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 92000 182414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 92000 200414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 92000 218414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 92000 236414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 92000 254414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 92000 272414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 92000 290414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 92000 308414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 92000 326414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 343794 92000 344414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 92000 362414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 379794 92000 380414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 397794 92000 398414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 415794 92000 416414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 433794 92000 434414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 451794 92000 452414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 469794 92000 470414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 487794 92000 488414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 92000 506414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 523794 92000 524414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 541794 92000 542414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 19794 119000 20414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 37794 119000 38414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 55794 119000 56414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 119000 74414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 119000 92414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 119000 110414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 119000 128414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 119000 146414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 119000 164414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 119000 182414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 119000 200414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 119000 218414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 119000 236414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 119000 254414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 119000 272414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 119000 290414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 119000 308414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 119000 326414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 343794 119000 344414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 119000 362414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 379794 119000 380414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 397794 119000 398414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 415794 119000 416414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 433794 119000 434414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 451794 119000 452414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 469794 119000 470414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 487794 119000 488414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 119000 506414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 523794 119000 524414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 541794 119000 542414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 19794 146000 20414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 37794 146000 38414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 55794 146000 56414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 146000 74414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 146000 92414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 146000 110414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 146000 128414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 146000 146414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 146000 164414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 146000 182414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 146000 200414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 146000 218414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 146000 236414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 146000 254414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 146000 272414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 146000 290414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 146000 308414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 146000 326414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 343794 146000 344414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 146000 362414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 379794 146000 380414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 397794 146000 398414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 415794 146000 416414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 433794 146000 434414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 451794 146000 452414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 469794 146000 470414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 487794 146000 488414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 146000 506414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 523794 146000 524414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 541794 146000 542414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 19794 173000 20414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 37794 173000 38414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 55794 173000 56414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 173000 74414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 173000 92414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 173000 110414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 173000 128414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 173000 146414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 173000 164414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 173000 182414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 173000 200414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 173000 218414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 173000 236414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 173000 254414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 173000 272414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 173000 290414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 173000 308414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 173000 326414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 343794 173000 344414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 173000 362414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 379794 173000 380414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 397794 173000 398414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 415794 173000 416414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 433794 173000 434414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 451794 173000 452414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 469794 173000 470414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 487794 173000 488414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 173000 506414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 523794 173000 524414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 541794 173000 542414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 19794 200000 20414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 37794 200000 38414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 55794 200000 56414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 200000 74414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 200000 92414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 200000 110414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 200000 128414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 200000 146414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 200000 164414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 200000 182414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 200000 200414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 200000 218414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 200000 236414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 200000 254414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 200000 272414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 200000 290414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 200000 308414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 200000 326414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 343794 200000 344414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 200000 362414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 379794 200000 380414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 397794 200000 398414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 415794 200000 416414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 433794 200000 434414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 451794 200000 452414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 469794 200000 470414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 487794 200000 488414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 200000 506414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 523794 200000 524414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 541794 200000 542414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 19794 227000 20414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 37794 227000 38414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 55794 227000 56414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 227000 74414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 227000 92414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 227000 110414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 227000 128414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 227000 146414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 227000 164414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 227000 182414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 227000 200414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 227000 218414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 227000 236414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 227000 254414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 227000 272414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 227000 290414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 227000 308414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 227000 326414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 343794 227000 344414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 227000 362414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 379794 227000 380414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 397794 227000 398414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 415794 227000 416414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 433794 227000 434414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 451794 227000 452414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 469794 227000 470414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 487794 227000 488414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 227000 506414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 523794 227000 524414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 541794 227000 542414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 19794 254000 20414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 37794 254000 38414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 55794 254000 56414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 254000 74414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 254000 92414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 254000 110414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 254000 128414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 254000 146414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 254000 164414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 254000 182414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 254000 200414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 254000 218414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 254000 236414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 254000 254414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 254000 272414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 254000 290414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 254000 308414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 254000 326414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 343794 254000 344414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 254000 362414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 379794 254000 380414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 397794 254000 398414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 415794 254000 416414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 433794 254000 434414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 451794 254000 452414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 469794 254000 470414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 487794 254000 488414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 254000 506414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 523794 254000 524414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 541794 254000 542414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 19794 281000 20414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 37794 281000 38414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 55794 281000 56414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 281000 74414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 281000 92414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 281000 110414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 281000 128414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 281000 146414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 281000 164414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 281000 182414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 281000 200414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 281000 218414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 281000 236414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 281000 254414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 281000 272414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 281000 290414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 281000 308414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 281000 326414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 343794 281000 344414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 281000 362414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 379794 281000 380414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 397794 281000 398414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 415794 281000 416414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 433794 281000 434414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 451794 281000 452414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 469794 281000 470414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 487794 281000 488414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 281000 506414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 523794 281000 524414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 541794 281000 542414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 19794 308000 20414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 37794 308000 38414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 55794 308000 56414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 308000 74414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 308000 92414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 308000 110414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 308000 128414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 308000 146414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 308000 164414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 308000 182414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 308000 200414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 308000 218414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 308000 236414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 308000 254414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 308000 272414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 308000 290414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 308000 308414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 308000 326414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 343794 308000 344414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 308000 362414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 379794 308000 380414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 397794 308000 398414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 415794 308000 416414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 433794 308000 434414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 451794 308000 452414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 469794 308000 470414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 487794 308000 488414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 308000 506414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 523794 308000 524414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 541794 308000 542414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 19794 335000 20414 338000 6 vccd1
port 532 nsew power input
rlabel metal4 s 37794 335000 38414 338000 6 vccd1
port 532 nsew power input
rlabel metal4 s 55794 335000 56414 338000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 335000 74414 338000 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 335000 92414 338000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 335000 110414 338000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 335000 128414 338000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 335000 146414 338000 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 335000 164414 338000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 335000 182414 338000 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 335000 200414 338000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 335000 218414 338000 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 335000 236414 338000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 335000 254414 338000 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 335000 272414 338000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 335000 290414 338000 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 335000 308414 338000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 335000 326414 338000 6 vccd1
port 532 nsew power input
rlabel metal4 s 343794 335000 344414 338000 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 335000 362414 338000 6 vccd1
port 532 nsew power input
rlabel metal4 s 379794 335000 380414 338000 6 vccd1
port 532 nsew power input
rlabel metal4 s 397794 335000 398414 338000 6 vccd1
port 532 nsew power input
rlabel metal4 s 415794 335000 416414 338000 6 vccd1
port 532 nsew power input
rlabel metal4 s 433794 335000 434414 338000 6 vccd1
port 532 nsew power input
rlabel metal4 s 451794 335000 452414 338000 6 vccd1
port 532 nsew power input
rlabel metal4 s 469794 335000 470414 338000 6 vccd1
port 532 nsew power input
rlabel metal4 s 487794 335000 488414 338000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 335000 506414 338000 6 vccd1
port 532 nsew power input
rlabel metal4 s 523794 335000 524414 338000 6 vccd1
port 532 nsew power input
rlabel metal4 s 541794 335000 542414 338000 6 vccd1
port 532 nsew power input
rlabel metal4 s 19794 362000 20414 365000 6 vccd1
port 532 nsew power input
rlabel metal4 s 37794 362000 38414 365000 6 vccd1
port 532 nsew power input
rlabel metal4 s 55794 362000 56414 365000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 362000 74414 365000 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 362000 92414 365000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 362000 110414 365000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 362000 128414 365000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 362000 146414 365000 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 362000 164414 365000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 362000 182414 365000 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 362000 200414 365000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 362000 218414 365000 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 362000 236414 365000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 362000 254414 365000 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 362000 272414 365000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 362000 290414 365000 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 362000 308414 365000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 362000 326414 365000 6 vccd1
port 532 nsew power input
rlabel metal4 s 343794 362000 344414 365000 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 362000 362414 365000 6 vccd1
port 532 nsew power input
rlabel metal4 s 379794 362000 380414 365000 6 vccd1
port 532 nsew power input
rlabel metal4 s 397794 362000 398414 365000 6 vccd1
port 532 nsew power input
rlabel metal4 s 415794 362000 416414 365000 6 vccd1
port 532 nsew power input
rlabel metal4 s 433794 362000 434414 365000 6 vccd1
port 532 nsew power input
rlabel metal4 s 451794 362000 452414 365000 6 vccd1
port 532 nsew power input
rlabel metal4 s 469794 362000 470414 365000 6 vccd1
port 532 nsew power input
rlabel metal4 s 487794 362000 488414 365000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 362000 506414 365000 6 vccd1
port 532 nsew power input
rlabel metal4 s 523794 362000 524414 365000 6 vccd1
port 532 nsew power input
rlabel metal4 s 541794 362000 542414 365000 6 vccd1
port 532 nsew power input
rlabel metal4 s 19794 389000 20414 392000 6 vccd1
port 532 nsew power input
rlabel metal4 s 37794 389000 38414 392000 6 vccd1
port 532 nsew power input
rlabel metal4 s 55794 389000 56414 392000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 389000 74414 392000 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 389000 92414 392000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 389000 110414 392000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 389000 128414 392000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 389000 146414 392000 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 389000 164414 392000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 389000 182414 392000 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 389000 200414 392000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 389000 218414 392000 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 389000 236414 392000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 389000 254414 392000 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 389000 272414 392000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 389000 290414 392000 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 389000 308414 392000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 389000 326414 392000 6 vccd1
port 532 nsew power input
rlabel metal4 s 343794 389000 344414 392000 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 389000 362414 392000 6 vccd1
port 532 nsew power input
rlabel metal4 s 379794 389000 380414 392000 6 vccd1
port 532 nsew power input
rlabel metal4 s 397794 389000 398414 392000 6 vccd1
port 532 nsew power input
rlabel metal4 s 415794 389000 416414 392000 6 vccd1
port 532 nsew power input
rlabel metal4 s 433794 389000 434414 392000 6 vccd1
port 532 nsew power input
rlabel metal4 s 451794 389000 452414 392000 6 vccd1
port 532 nsew power input
rlabel metal4 s 469794 389000 470414 392000 6 vccd1
port 532 nsew power input
rlabel metal4 s 487794 389000 488414 392000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 389000 506414 392000 6 vccd1
port 532 nsew power input
rlabel metal4 s 523794 389000 524414 392000 6 vccd1
port 532 nsew power input
rlabel metal4 s 541794 389000 542414 392000 6 vccd1
port 532 nsew power input
rlabel metal4 s 19794 416000 20414 419000 6 vccd1
port 532 nsew power input
rlabel metal4 s 37794 416000 38414 419000 6 vccd1
port 532 nsew power input
rlabel metal4 s 55794 416000 56414 419000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 416000 74414 419000 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 416000 92414 419000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 416000 110414 419000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 416000 128414 419000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 416000 146414 419000 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 416000 164414 419000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 416000 182414 419000 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 416000 200414 419000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 416000 218414 419000 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 416000 236414 419000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 416000 254414 419000 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 416000 272414 419000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 416000 290414 419000 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 416000 308414 419000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 416000 326414 419000 6 vccd1
port 532 nsew power input
rlabel metal4 s 343794 416000 344414 419000 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 416000 362414 419000 6 vccd1
port 532 nsew power input
rlabel metal4 s 379794 416000 380414 419000 6 vccd1
port 532 nsew power input
rlabel metal4 s 397794 416000 398414 419000 6 vccd1
port 532 nsew power input
rlabel metal4 s 415794 416000 416414 419000 6 vccd1
port 532 nsew power input
rlabel metal4 s 433794 416000 434414 419000 6 vccd1
port 532 nsew power input
rlabel metal4 s 451794 416000 452414 419000 6 vccd1
port 532 nsew power input
rlabel metal4 s 469794 416000 470414 419000 6 vccd1
port 532 nsew power input
rlabel metal4 s 487794 416000 488414 419000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 416000 506414 419000 6 vccd1
port 532 nsew power input
rlabel metal4 s 523794 416000 524414 419000 6 vccd1
port 532 nsew power input
rlabel metal4 s 541794 416000 542414 419000 6 vccd1
port 532 nsew power input
rlabel metal4 s 19794 443000 20414 446000 6 vccd1
port 532 nsew power input
rlabel metal4 s 37794 443000 38414 446000 6 vccd1
port 532 nsew power input
rlabel metal4 s 55794 443000 56414 446000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 443000 74414 446000 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 443000 92414 446000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 443000 110414 446000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 443000 128414 446000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 443000 146414 446000 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 443000 164414 446000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 443000 182414 446000 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 443000 200414 446000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 443000 218414 446000 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 443000 236414 446000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 443000 254414 446000 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 443000 272414 446000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 443000 290414 446000 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 443000 308414 446000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 443000 326414 446000 6 vccd1
port 532 nsew power input
rlabel metal4 s 343794 443000 344414 446000 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 443000 362414 446000 6 vccd1
port 532 nsew power input
rlabel metal4 s 379794 443000 380414 446000 6 vccd1
port 532 nsew power input
rlabel metal4 s 397794 443000 398414 446000 6 vccd1
port 532 nsew power input
rlabel metal4 s 415794 443000 416414 446000 6 vccd1
port 532 nsew power input
rlabel metal4 s 433794 443000 434414 446000 6 vccd1
port 532 nsew power input
rlabel metal4 s 451794 443000 452414 446000 6 vccd1
port 532 nsew power input
rlabel metal4 s 469794 443000 470414 446000 6 vccd1
port 532 nsew power input
rlabel metal4 s 487794 443000 488414 446000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 443000 506414 446000 6 vccd1
port 532 nsew power input
rlabel metal4 s 523794 443000 524414 446000 6 vccd1
port 532 nsew power input
rlabel metal4 s 541794 443000 542414 446000 6 vccd1
port 532 nsew power input
rlabel metal4 s 19794 470000 20414 473000 6 vccd1
port 532 nsew power input
rlabel metal4 s 37794 470000 38414 473000 6 vccd1
port 532 nsew power input
rlabel metal4 s 55794 470000 56414 473000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 470000 74414 473000 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 470000 92414 473000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 470000 110414 473000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 470000 128414 473000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 470000 146414 473000 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 470000 164414 473000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 470000 182414 473000 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 470000 200414 473000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 470000 218414 473000 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 470000 236414 473000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 470000 254414 473000 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 470000 272414 473000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 470000 290414 473000 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 470000 308414 473000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 470000 326414 473000 6 vccd1
port 532 nsew power input
rlabel metal4 s 343794 470000 344414 473000 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 470000 362414 473000 6 vccd1
port 532 nsew power input
rlabel metal4 s 379794 470000 380414 473000 6 vccd1
port 532 nsew power input
rlabel metal4 s 397794 470000 398414 473000 6 vccd1
port 532 nsew power input
rlabel metal4 s 415794 470000 416414 473000 6 vccd1
port 532 nsew power input
rlabel metal4 s 433794 470000 434414 473000 6 vccd1
port 532 nsew power input
rlabel metal4 s 451794 470000 452414 473000 6 vccd1
port 532 nsew power input
rlabel metal4 s 469794 470000 470414 473000 6 vccd1
port 532 nsew power input
rlabel metal4 s 487794 470000 488414 473000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 470000 506414 473000 6 vccd1
port 532 nsew power input
rlabel metal4 s 523794 470000 524414 473000 6 vccd1
port 532 nsew power input
rlabel metal4 s 541794 470000 542414 473000 6 vccd1
port 532 nsew power input
rlabel metal4 s 19794 497000 20414 500000 6 vccd1
port 532 nsew power input
rlabel metal4 s 37794 497000 38414 500000 6 vccd1
port 532 nsew power input
rlabel metal4 s 55794 497000 56414 500000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 497000 74414 500000 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 497000 92414 500000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 497000 110414 500000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 497000 128414 500000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 497000 146414 500000 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 497000 164414 500000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 497000 182414 500000 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 497000 200414 500000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 497000 218414 500000 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 497000 236414 500000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 497000 254414 500000 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 497000 272414 500000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 497000 290414 500000 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 497000 308414 500000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 497000 326414 500000 6 vccd1
port 532 nsew power input
rlabel metal4 s 343794 497000 344414 500000 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 497000 362414 500000 6 vccd1
port 532 nsew power input
rlabel metal4 s 379794 497000 380414 500000 6 vccd1
port 532 nsew power input
rlabel metal4 s 397794 497000 398414 500000 6 vccd1
port 532 nsew power input
rlabel metal4 s 415794 497000 416414 500000 6 vccd1
port 532 nsew power input
rlabel metal4 s 433794 497000 434414 500000 6 vccd1
port 532 nsew power input
rlabel metal4 s 451794 497000 452414 500000 6 vccd1
port 532 nsew power input
rlabel metal4 s 469794 497000 470414 500000 6 vccd1
port 532 nsew power input
rlabel metal4 s 487794 497000 488414 500000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 497000 506414 500000 6 vccd1
port 532 nsew power input
rlabel metal4 s 523794 497000 524414 500000 6 vccd1
port 532 nsew power input
rlabel metal4 s 541794 497000 542414 500000 6 vccd1
port 532 nsew power input
rlabel metal4 s 19794 524000 20414 527000 6 vccd1
port 532 nsew power input
rlabel metal4 s 37794 524000 38414 527000 6 vccd1
port 532 nsew power input
rlabel metal4 s 55794 524000 56414 527000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 524000 74414 527000 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 524000 92414 527000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 524000 110414 527000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 524000 128414 527000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 524000 146414 527000 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 524000 164414 527000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 524000 182414 527000 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 524000 200414 527000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 524000 218414 527000 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 524000 236414 527000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 524000 254414 527000 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 524000 272414 527000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 524000 290414 527000 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 524000 308414 527000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 524000 326414 527000 6 vccd1
port 532 nsew power input
rlabel metal4 s 343794 524000 344414 527000 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 524000 362414 527000 6 vccd1
port 532 nsew power input
rlabel metal4 s 379794 524000 380414 527000 6 vccd1
port 532 nsew power input
rlabel metal4 s 397794 524000 398414 527000 6 vccd1
port 532 nsew power input
rlabel metal4 s 415794 524000 416414 527000 6 vccd1
port 532 nsew power input
rlabel metal4 s 433794 524000 434414 527000 6 vccd1
port 532 nsew power input
rlabel metal4 s 451794 524000 452414 527000 6 vccd1
port 532 nsew power input
rlabel metal4 s 469794 524000 470414 527000 6 vccd1
port 532 nsew power input
rlabel metal4 s 487794 524000 488414 527000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 524000 506414 527000 6 vccd1
port 532 nsew power input
rlabel metal4 s 523794 524000 524414 527000 6 vccd1
port 532 nsew power input
rlabel metal4 s 541794 524000 542414 527000 6 vccd1
port 532 nsew power input
rlabel metal4 s 19794 551000 20414 554000 6 vccd1
port 532 nsew power input
rlabel metal4 s 37794 551000 38414 554000 6 vccd1
port 532 nsew power input
rlabel metal4 s 55794 551000 56414 554000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 551000 74414 554000 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 551000 92414 554000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 551000 110414 554000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 551000 128414 554000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 551000 146414 554000 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 551000 164414 554000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 551000 182414 554000 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 551000 200414 554000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 551000 218414 554000 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 551000 236414 554000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 551000 254414 554000 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 551000 272414 554000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 551000 290414 554000 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 551000 308414 554000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 551000 326414 554000 6 vccd1
port 532 nsew power input
rlabel metal4 s 343794 551000 344414 554000 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 551000 362414 554000 6 vccd1
port 532 nsew power input
rlabel metal4 s 379794 551000 380414 554000 6 vccd1
port 532 nsew power input
rlabel metal4 s 397794 551000 398414 554000 6 vccd1
port 532 nsew power input
rlabel metal4 s 415794 551000 416414 554000 6 vccd1
port 532 nsew power input
rlabel metal4 s 433794 551000 434414 554000 6 vccd1
port 532 nsew power input
rlabel metal4 s 451794 551000 452414 554000 6 vccd1
port 532 nsew power input
rlabel metal4 s 469794 551000 470414 554000 6 vccd1
port 532 nsew power input
rlabel metal4 s 487794 551000 488414 554000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 551000 506414 554000 6 vccd1
port 532 nsew power input
rlabel metal4 s 523794 551000 524414 554000 6 vccd1
port 532 nsew power input
rlabel metal4 s 541794 551000 542414 554000 6 vccd1
port 532 nsew power input
rlabel metal4 s 19794 578000 20414 581000 6 vccd1
port 532 nsew power input
rlabel metal4 s 37794 578000 38414 581000 6 vccd1
port 532 nsew power input
rlabel metal4 s 55794 578000 56414 581000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 578000 74414 581000 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 578000 92414 581000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 578000 110414 581000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 578000 128414 581000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 578000 146414 581000 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 578000 164414 581000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 578000 182414 581000 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 578000 200414 581000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 578000 218414 581000 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 578000 236414 581000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 578000 254414 581000 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 578000 272414 581000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 578000 290414 581000 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 578000 308414 581000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 578000 326414 581000 6 vccd1
port 532 nsew power input
rlabel metal4 s 343794 578000 344414 581000 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 578000 362414 581000 6 vccd1
port 532 nsew power input
rlabel metal4 s 379794 578000 380414 581000 6 vccd1
port 532 nsew power input
rlabel metal4 s 397794 578000 398414 581000 6 vccd1
port 532 nsew power input
rlabel metal4 s 415794 578000 416414 581000 6 vccd1
port 532 nsew power input
rlabel metal4 s 433794 578000 434414 581000 6 vccd1
port 532 nsew power input
rlabel metal4 s 451794 578000 452414 581000 6 vccd1
port 532 nsew power input
rlabel metal4 s 469794 578000 470414 581000 6 vccd1
port 532 nsew power input
rlabel metal4 s 487794 578000 488414 581000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 578000 506414 581000 6 vccd1
port 532 nsew power input
rlabel metal4 s 523794 578000 524414 581000 6 vccd1
port 532 nsew power input
rlabel metal4 s 541794 578000 542414 581000 6 vccd1
port 532 nsew power input
rlabel metal4 s 19794 605000 20414 608000 6 vccd1
port 532 nsew power input
rlabel metal4 s 37794 605000 38414 608000 6 vccd1
port 532 nsew power input
rlabel metal4 s 55794 605000 56414 608000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 605000 74414 608000 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 605000 92414 608000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 605000 110414 608000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 605000 128414 608000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 605000 146414 608000 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 605000 164414 608000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 605000 182414 608000 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 605000 200414 608000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 605000 218414 608000 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 605000 236414 608000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 605000 254414 608000 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 605000 272414 608000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 605000 290414 608000 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 605000 308414 608000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 605000 326414 608000 6 vccd1
port 532 nsew power input
rlabel metal4 s 343794 605000 344414 608000 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 605000 362414 608000 6 vccd1
port 532 nsew power input
rlabel metal4 s 379794 605000 380414 608000 6 vccd1
port 532 nsew power input
rlabel metal4 s 397794 605000 398414 608000 6 vccd1
port 532 nsew power input
rlabel metal4 s 415794 605000 416414 608000 6 vccd1
port 532 nsew power input
rlabel metal4 s 433794 605000 434414 608000 6 vccd1
port 532 nsew power input
rlabel metal4 s 451794 605000 452414 608000 6 vccd1
port 532 nsew power input
rlabel metal4 s 469794 605000 470414 608000 6 vccd1
port 532 nsew power input
rlabel metal4 s 487794 605000 488414 608000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 605000 506414 608000 6 vccd1
port 532 nsew power input
rlabel metal4 s 523794 605000 524414 608000 6 vccd1
port 532 nsew power input
rlabel metal4 s 541794 605000 542414 608000 6 vccd1
port 532 nsew power input
rlabel metal4 s 19794 632000 20414 635000 6 vccd1
port 532 nsew power input
rlabel metal4 s 37794 632000 38414 635000 6 vccd1
port 532 nsew power input
rlabel metal4 s 55794 632000 56414 635000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 632000 74414 635000 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 632000 92414 635000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 632000 110414 635000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 632000 128414 635000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 632000 146414 635000 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 632000 164414 635000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 632000 182414 635000 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 632000 200414 635000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 632000 218414 635000 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 632000 236414 635000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 632000 254414 635000 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 632000 272414 635000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 632000 290414 635000 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 632000 308414 635000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 632000 326414 635000 6 vccd1
port 532 nsew power input
rlabel metal4 s 343794 632000 344414 635000 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 632000 362414 635000 6 vccd1
port 532 nsew power input
rlabel metal4 s 379794 632000 380414 635000 6 vccd1
port 532 nsew power input
rlabel metal4 s 397794 632000 398414 635000 6 vccd1
port 532 nsew power input
rlabel metal4 s 415794 632000 416414 635000 6 vccd1
port 532 nsew power input
rlabel metal4 s 433794 632000 434414 635000 6 vccd1
port 532 nsew power input
rlabel metal4 s 451794 632000 452414 635000 6 vccd1
port 532 nsew power input
rlabel metal4 s 469794 632000 470414 635000 6 vccd1
port 532 nsew power input
rlabel metal4 s 487794 632000 488414 635000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 632000 506414 635000 6 vccd1
port 532 nsew power input
rlabel metal4 s 523794 632000 524414 635000 6 vccd1
port 532 nsew power input
rlabel metal4 s 541794 632000 542414 635000 6 vccd1
port 532 nsew power input
rlabel metal4 s 19794 659000 20414 662000 6 vccd1
port 532 nsew power input
rlabel metal4 s 37794 659000 38414 662000 6 vccd1
port 532 nsew power input
rlabel metal4 s 55794 659000 56414 662000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 659000 74414 662000 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 659000 92414 662000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 659000 110414 662000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 659000 128414 662000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 659000 146414 662000 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 659000 164414 662000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 659000 182414 662000 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 659000 200414 662000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 659000 218414 662000 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 659000 236414 662000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 659000 254414 662000 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 659000 272414 662000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 659000 290414 662000 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 659000 308414 662000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 659000 326414 662000 6 vccd1
port 532 nsew power input
rlabel metal4 s 343794 659000 344414 662000 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 659000 362414 662000 6 vccd1
port 532 nsew power input
rlabel metal4 s 379794 659000 380414 662000 6 vccd1
port 532 nsew power input
rlabel metal4 s 397794 659000 398414 662000 6 vccd1
port 532 nsew power input
rlabel metal4 s 415794 659000 416414 662000 6 vccd1
port 532 nsew power input
rlabel metal4 s 433794 659000 434414 662000 6 vccd1
port 532 nsew power input
rlabel metal4 s 451794 659000 452414 662000 6 vccd1
port 532 nsew power input
rlabel metal4 s 469794 659000 470414 662000 6 vccd1
port 532 nsew power input
rlabel metal4 s 487794 659000 488414 662000 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 659000 506414 662000 6 vccd1
port 532 nsew power input
rlabel metal4 s 523794 659000 524414 662000 6 vccd1
port 532 nsew power input
rlabel metal4 s 541794 659000 542414 662000 6 vccd1
port 532 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 532 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 532 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 19794 686000 20414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 37794 686000 38414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 55794 686000 56414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 686000 74414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 686000 92414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 686000 110414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 686000 128414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 686000 146414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 686000 164414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 686000 182414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 686000 200414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 686000 218414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 686000 236414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 686000 254414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 686000 272414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 686000 290414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 686000 308414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 686000 326414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 343794 686000 344414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 686000 362414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 379794 686000 380414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 397794 686000 398414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 415794 686000 416414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 433794 686000 434414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 451794 686000 452414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 469794 686000 470414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 487794 686000 488414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 686000 506414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 523794 686000 524414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 541794 686000 542414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 559794 -1894 560414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 11866 586890 12486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 29866 586890 30486 6 vssd1
port 533 nsew ground input
rlabel metal5 s 28794 39806 551414 40426 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 47866 586890 48486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 65866 586890 66486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 83866 586890 84486 6 vssd1
port 533 nsew ground input
rlabel metal5 s 28794 93806 551414 94426 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 101866 586890 102486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 119866 586890 120486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 137866 586890 138486 6 vssd1
port 533 nsew ground input
rlabel metal5 s 28794 147806 551414 148426 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 155866 586890 156486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 173866 586890 174486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 191866 586890 192486 6 vssd1
port 533 nsew ground input
rlabel metal5 s 28794 201806 551414 202426 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 209866 586890 210486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 227866 586890 228486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 245866 586890 246486 6 vssd1
port 533 nsew ground input
rlabel metal5 s 28794 255806 551414 256426 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 263866 586890 264486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 281866 586890 282486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 299866 586890 300486 6 vssd1
port 533 nsew ground input
rlabel metal5 s 28794 309806 551414 310426 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 317866 586890 318486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 335866 586890 336486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 353866 586890 354486 6 vssd1
port 533 nsew ground input
rlabel metal5 s 28794 363806 551414 364426 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 371866 586890 372486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 389866 586890 390486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 407866 586890 408486 6 vssd1
port 533 nsew ground input
rlabel metal5 s 28794 417806 551414 418426 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 425866 586890 426486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 443866 586890 444486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 461866 586890 462486 6 vssd1
port 533 nsew ground input
rlabel metal5 s 28794 471806 551414 472426 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 479866 586890 480486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 497866 586890 498486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 515866 586890 516486 6 vssd1
port 533 nsew ground input
rlabel metal5 s 28794 525806 551414 526426 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 533866 586890 534486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 551866 586890 552486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 569866 586890 570486 6 vssd1
port 533 nsew ground input
rlabel metal5 s 28794 579806 551414 580426 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 587866 586890 588486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 605866 586890 606486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 623866 586890 624486 6 vssd1
port 533 nsew ground input
rlabel metal5 s 28794 633806 551414 634426 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 641866 586890 642486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 659866 586890 660486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 677866 586890 678486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 695866 586890 696486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 28794 -1894 29414 14000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 46794 -1894 47414 14000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 -1894 83414 14000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 -1894 101414 14000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 -1894 119414 14000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 -1894 137414 14000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 -1894 155414 14000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 -1894 173414 14000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 -1894 191414 14000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 -1894 209414 14000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 -1894 227414 14000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 -1894 245414 14000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 -1894 263414 14000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 -1894 281414 14000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 -1894 299414 14000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 -1894 317414 14000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 -1894 335414 14000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 352794 -1894 353414 14000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 370794 -1894 371414 14000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 388794 -1894 389414 14000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 406794 -1894 407414 14000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 424794 -1894 425414 14000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 442794 -1894 443414 14000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 460794 -1894 461414 14000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 478794 -1894 479414 14000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 496794 -1894 497414 14000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 514794 -1894 515414 14000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 532794 -1894 533414 14000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 550794 -1894 551414 14000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 28794 38000 29414 41000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 46794 38000 47414 41000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 64794 -1894 65414 41000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 38000 83414 41000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 38000 101414 41000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 38000 119414 41000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 38000 137414 41000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 38000 155414 41000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 38000 173414 41000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 38000 191414 41000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 38000 209414 41000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 38000 227414 41000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 38000 245414 41000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 38000 263414 41000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 38000 281414 41000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 38000 299414 41000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 38000 317414 41000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 38000 335414 41000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 352794 38000 353414 41000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 370794 38000 371414 41000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 388794 38000 389414 41000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 406794 38000 407414 41000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 424794 38000 425414 41000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 442794 38000 443414 41000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 460794 38000 461414 41000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 478794 38000 479414 41000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 496794 38000 497414 41000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 514794 38000 515414 41000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 532794 38000 533414 41000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 550794 38000 551414 41000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 28794 65000 29414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 46794 65000 47414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 64794 65000 65414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 65000 83414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 65000 101414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 65000 119414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 65000 137414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 65000 155414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 65000 173414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 65000 191414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 65000 209414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 65000 227414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 65000 245414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 65000 263414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 65000 281414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 65000 299414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 65000 317414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 65000 335414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 352794 65000 353414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 370794 65000 371414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 388794 65000 389414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 406794 65000 407414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 424794 65000 425414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 442794 65000 443414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 460794 65000 461414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 478794 65000 479414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 496794 65000 497414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 514794 65000 515414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 532794 65000 533414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 550794 65000 551414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 28794 92000 29414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 46794 92000 47414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 64794 92000 65414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 92000 83414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 92000 101414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 92000 119414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 92000 137414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 92000 155414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 92000 173414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 92000 191414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 92000 209414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 92000 227414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 92000 245414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 92000 263414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 92000 281414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 92000 299414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 92000 317414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 92000 335414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 352794 92000 353414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 370794 92000 371414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 388794 92000 389414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 406794 92000 407414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 424794 92000 425414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 442794 92000 443414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 460794 92000 461414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 478794 92000 479414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 496794 92000 497414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 514794 92000 515414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 532794 92000 533414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 550794 92000 551414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 28794 119000 29414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 46794 119000 47414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 64794 119000 65414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 119000 83414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 119000 101414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 119000 119414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 119000 137414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 119000 155414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 119000 173414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 119000 191414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 119000 209414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 119000 227414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 119000 245414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 119000 263414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 119000 281414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 119000 299414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 119000 317414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 119000 335414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 352794 119000 353414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 370794 119000 371414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 388794 119000 389414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 406794 119000 407414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 424794 119000 425414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 442794 119000 443414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 460794 119000 461414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 478794 119000 479414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 496794 119000 497414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 514794 119000 515414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 532794 119000 533414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 550794 119000 551414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 28794 146000 29414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 46794 146000 47414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 64794 146000 65414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 146000 83414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 146000 101414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 146000 119414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 146000 137414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 146000 155414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 146000 173414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 146000 191414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 146000 209414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 146000 227414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 146000 245414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 146000 263414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 146000 281414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 146000 299414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 146000 317414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 146000 335414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 352794 146000 353414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 370794 146000 371414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 388794 146000 389414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 406794 146000 407414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 424794 146000 425414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 442794 146000 443414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 460794 146000 461414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 478794 146000 479414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 496794 146000 497414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 514794 146000 515414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 532794 146000 533414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 550794 146000 551414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 28794 173000 29414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 46794 173000 47414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 64794 173000 65414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 173000 83414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 173000 101414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 173000 119414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 173000 137414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 173000 155414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 173000 173414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 173000 191414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 173000 209414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 173000 227414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 173000 245414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 173000 263414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 173000 281414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 173000 299414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 173000 317414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 173000 335414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 352794 173000 353414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 370794 173000 371414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 388794 173000 389414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 406794 173000 407414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 424794 173000 425414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 442794 173000 443414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 460794 173000 461414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 478794 173000 479414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 496794 173000 497414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 514794 173000 515414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 532794 173000 533414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 550794 173000 551414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 28794 200000 29414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 46794 200000 47414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 64794 200000 65414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 200000 83414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 200000 101414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 200000 119414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 200000 137414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 200000 155414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 200000 173414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 200000 191414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 200000 209414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 200000 227414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 200000 245414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 200000 263414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 200000 281414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 200000 299414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 200000 317414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 200000 335414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 352794 200000 353414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 370794 200000 371414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 388794 200000 389414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 406794 200000 407414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 424794 200000 425414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 442794 200000 443414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 460794 200000 461414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 478794 200000 479414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 496794 200000 497414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 514794 200000 515414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 532794 200000 533414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 550794 200000 551414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 28794 227000 29414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 46794 227000 47414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 64794 227000 65414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 227000 83414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 227000 101414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 227000 119414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 227000 137414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 227000 155414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 227000 173414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 227000 191414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 227000 209414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 227000 227414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 227000 245414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 227000 263414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 227000 281414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 227000 299414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 227000 317414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 227000 335414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 352794 227000 353414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 370794 227000 371414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 388794 227000 389414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 406794 227000 407414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 424794 227000 425414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 442794 227000 443414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 460794 227000 461414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 478794 227000 479414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 496794 227000 497414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 514794 227000 515414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 532794 227000 533414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 550794 227000 551414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 28794 254000 29414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 46794 254000 47414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 64794 254000 65414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 254000 83414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 254000 101414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 254000 119414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 254000 137414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 254000 155414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 254000 173414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 254000 191414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 254000 209414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 254000 227414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 254000 245414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 254000 263414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 254000 281414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 254000 299414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 254000 317414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 254000 335414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 352794 254000 353414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 370794 254000 371414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 388794 254000 389414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 406794 254000 407414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 424794 254000 425414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 442794 254000 443414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 460794 254000 461414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 478794 254000 479414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 496794 254000 497414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 514794 254000 515414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 532794 254000 533414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 550794 254000 551414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 28794 281000 29414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 46794 281000 47414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 64794 281000 65414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 281000 83414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 281000 101414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 281000 119414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 281000 137414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 281000 155414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 281000 173414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 281000 191414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 281000 209414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 281000 227414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 281000 245414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 281000 263414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 281000 281414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 281000 299414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 281000 317414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 281000 335414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 352794 281000 353414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 370794 281000 371414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 388794 281000 389414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 406794 281000 407414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 424794 281000 425414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 442794 281000 443414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 460794 281000 461414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 478794 281000 479414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 496794 281000 497414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 514794 281000 515414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 532794 281000 533414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 550794 281000 551414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 28794 308000 29414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 46794 308000 47414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 64794 308000 65414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 308000 83414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 308000 101414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 308000 119414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 308000 137414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 308000 155414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 308000 173414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 308000 191414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 308000 209414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 308000 227414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 308000 245414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 308000 263414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 308000 281414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 308000 299414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 308000 317414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 308000 335414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 352794 308000 353414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 370794 308000 371414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 388794 308000 389414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 406794 308000 407414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 424794 308000 425414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 442794 308000 443414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 460794 308000 461414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 478794 308000 479414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 496794 308000 497414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 514794 308000 515414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 532794 308000 533414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 550794 308000 551414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 28794 335000 29414 338000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 46794 335000 47414 338000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 64794 335000 65414 338000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 335000 83414 338000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 335000 101414 338000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 335000 119414 338000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 335000 137414 338000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 335000 155414 338000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 335000 173414 338000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 335000 191414 338000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 335000 209414 338000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 335000 227414 338000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 335000 245414 338000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 335000 263414 338000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 335000 281414 338000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 335000 299414 338000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 335000 317414 338000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 335000 335414 338000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 352794 335000 353414 338000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 370794 335000 371414 338000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 388794 335000 389414 338000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 406794 335000 407414 338000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 424794 335000 425414 338000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 442794 335000 443414 338000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 460794 335000 461414 338000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 478794 335000 479414 338000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 496794 335000 497414 338000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 514794 335000 515414 338000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 532794 335000 533414 338000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 550794 335000 551414 338000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 28794 362000 29414 365000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 46794 362000 47414 365000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 64794 362000 65414 365000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 362000 83414 365000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 362000 101414 365000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 362000 119414 365000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 362000 137414 365000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 362000 155414 365000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 362000 173414 365000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 362000 191414 365000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 362000 209414 365000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 362000 227414 365000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 362000 245414 365000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 362000 263414 365000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 362000 281414 365000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 362000 299414 365000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 362000 317414 365000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 362000 335414 365000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 352794 362000 353414 365000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 370794 362000 371414 365000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 388794 362000 389414 365000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 406794 362000 407414 365000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 424794 362000 425414 365000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 442794 362000 443414 365000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 460794 362000 461414 365000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 478794 362000 479414 365000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 496794 362000 497414 365000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 514794 362000 515414 365000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 532794 362000 533414 365000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 550794 362000 551414 365000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 28794 389000 29414 392000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 46794 389000 47414 392000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 64794 389000 65414 392000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 389000 83414 392000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 389000 101414 392000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 389000 119414 392000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 389000 137414 392000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 389000 155414 392000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 389000 173414 392000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 389000 191414 392000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 389000 209414 392000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 389000 227414 392000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 389000 245414 392000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 389000 263414 392000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 389000 281414 392000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 389000 299414 392000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 389000 317414 392000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 389000 335414 392000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 352794 389000 353414 392000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 370794 389000 371414 392000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 388794 389000 389414 392000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 406794 389000 407414 392000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 424794 389000 425414 392000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 442794 389000 443414 392000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 460794 389000 461414 392000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 478794 389000 479414 392000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 496794 389000 497414 392000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 514794 389000 515414 392000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 532794 389000 533414 392000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 550794 389000 551414 392000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 28794 416000 29414 419000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 46794 416000 47414 419000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 64794 416000 65414 419000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 416000 83414 419000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 416000 101414 419000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 416000 119414 419000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 416000 137414 419000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 416000 155414 419000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 416000 173414 419000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 416000 191414 419000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 416000 209414 419000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 416000 227414 419000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 416000 245414 419000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 416000 263414 419000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 416000 281414 419000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 416000 299414 419000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 416000 317414 419000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 416000 335414 419000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 352794 416000 353414 419000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 370794 416000 371414 419000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 388794 416000 389414 419000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 406794 416000 407414 419000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 424794 416000 425414 419000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 442794 416000 443414 419000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 460794 416000 461414 419000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 478794 416000 479414 419000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 496794 416000 497414 419000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 514794 416000 515414 419000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 532794 416000 533414 419000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 550794 416000 551414 419000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 28794 443000 29414 446000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 46794 443000 47414 446000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 64794 443000 65414 446000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 443000 83414 446000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 443000 101414 446000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 443000 119414 446000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 443000 137414 446000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 443000 155414 446000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 443000 173414 446000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 443000 191414 446000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 443000 209414 446000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 443000 227414 446000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 443000 245414 446000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 443000 263414 446000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 443000 281414 446000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 443000 299414 446000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 443000 317414 446000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 443000 335414 446000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 352794 443000 353414 446000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 370794 443000 371414 446000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 388794 443000 389414 446000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 406794 443000 407414 446000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 424794 443000 425414 446000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 442794 443000 443414 446000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 460794 443000 461414 446000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 478794 443000 479414 446000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 496794 443000 497414 446000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 514794 443000 515414 446000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 532794 443000 533414 446000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 550794 443000 551414 446000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 28794 470000 29414 473000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 46794 470000 47414 473000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 64794 470000 65414 473000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 470000 83414 473000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 470000 101414 473000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 470000 119414 473000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 470000 137414 473000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 470000 155414 473000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 470000 173414 473000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 470000 191414 473000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 470000 209414 473000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 470000 227414 473000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 470000 245414 473000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 470000 263414 473000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 470000 281414 473000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 470000 299414 473000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 470000 317414 473000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 470000 335414 473000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 352794 470000 353414 473000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 370794 470000 371414 473000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 388794 470000 389414 473000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 406794 470000 407414 473000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 424794 470000 425414 473000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 442794 470000 443414 473000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 460794 470000 461414 473000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 478794 470000 479414 473000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 496794 470000 497414 473000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 514794 470000 515414 473000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 532794 470000 533414 473000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 550794 470000 551414 473000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 28794 497000 29414 500000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 46794 497000 47414 500000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 64794 497000 65414 500000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 497000 83414 500000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 497000 101414 500000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 497000 119414 500000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 497000 137414 500000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 497000 155414 500000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 497000 173414 500000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 497000 191414 500000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 497000 209414 500000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 497000 227414 500000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 497000 245414 500000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 497000 263414 500000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 497000 281414 500000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 497000 299414 500000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 497000 317414 500000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 497000 335414 500000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 352794 497000 353414 500000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 370794 497000 371414 500000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 388794 497000 389414 500000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 406794 497000 407414 500000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 424794 497000 425414 500000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 442794 497000 443414 500000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 460794 497000 461414 500000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 478794 497000 479414 500000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 496794 497000 497414 500000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 514794 497000 515414 500000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 532794 497000 533414 500000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 550794 497000 551414 500000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 28794 524000 29414 527000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 46794 524000 47414 527000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 64794 524000 65414 527000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 524000 83414 527000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 524000 101414 527000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 524000 119414 527000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 524000 137414 527000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 524000 155414 527000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 524000 173414 527000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 524000 191414 527000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 524000 209414 527000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 524000 227414 527000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 524000 245414 527000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 524000 263414 527000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 524000 281414 527000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 524000 299414 527000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 524000 317414 527000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 524000 335414 527000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 352794 524000 353414 527000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 370794 524000 371414 527000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 388794 524000 389414 527000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 406794 524000 407414 527000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 424794 524000 425414 527000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 442794 524000 443414 527000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 460794 524000 461414 527000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 478794 524000 479414 527000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 496794 524000 497414 527000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 514794 524000 515414 527000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 532794 524000 533414 527000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 550794 524000 551414 527000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 28794 551000 29414 554000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 46794 551000 47414 554000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 64794 551000 65414 554000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 551000 83414 554000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 551000 101414 554000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 551000 119414 554000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 551000 137414 554000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 551000 155414 554000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 551000 173414 554000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 551000 191414 554000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 551000 209414 554000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 551000 227414 554000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 551000 245414 554000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 551000 263414 554000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 551000 281414 554000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 551000 299414 554000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 551000 317414 554000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 551000 335414 554000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 352794 551000 353414 554000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 370794 551000 371414 554000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 388794 551000 389414 554000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 406794 551000 407414 554000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 424794 551000 425414 554000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 442794 551000 443414 554000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 460794 551000 461414 554000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 478794 551000 479414 554000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 496794 551000 497414 554000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 514794 551000 515414 554000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 532794 551000 533414 554000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 550794 551000 551414 554000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 28794 578000 29414 581000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 46794 578000 47414 581000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 64794 578000 65414 581000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 578000 83414 581000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 578000 101414 581000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 578000 119414 581000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 578000 137414 581000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 578000 155414 581000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 578000 173414 581000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 578000 191414 581000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 578000 209414 581000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 578000 227414 581000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 578000 245414 581000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 578000 263414 581000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 578000 281414 581000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 578000 299414 581000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 578000 317414 581000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 578000 335414 581000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 352794 578000 353414 581000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 370794 578000 371414 581000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 388794 578000 389414 581000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 406794 578000 407414 581000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 424794 578000 425414 581000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 442794 578000 443414 581000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 460794 578000 461414 581000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 478794 578000 479414 581000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 496794 578000 497414 581000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 514794 578000 515414 581000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 532794 578000 533414 581000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 550794 578000 551414 581000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 28794 605000 29414 608000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 46794 605000 47414 608000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 64794 605000 65414 608000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 605000 83414 608000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 605000 101414 608000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 605000 119414 608000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 605000 137414 608000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 605000 155414 608000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 605000 173414 608000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 605000 191414 608000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 605000 209414 608000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 605000 227414 608000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 605000 245414 608000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 605000 263414 608000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 605000 281414 608000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 605000 299414 608000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 605000 317414 608000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 605000 335414 608000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 352794 605000 353414 608000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 370794 605000 371414 608000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 388794 605000 389414 608000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 406794 605000 407414 608000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 424794 605000 425414 608000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 442794 605000 443414 608000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 460794 605000 461414 608000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 478794 605000 479414 608000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 496794 605000 497414 608000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 514794 605000 515414 608000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 532794 605000 533414 608000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 550794 605000 551414 608000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 28794 632000 29414 635000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 46794 632000 47414 635000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 64794 632000 65414 635000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 632000 83414 635000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 632000 101414 635000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 632000 119414 635000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 632000 137414 635000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 632000 155414 635000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 632000 173414 635000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 632000 191414 635000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 632000 209414 635000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 632000 227414 635000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 632000 245414 635000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 632000 263414 635000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 632000 281414 635000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 632000 299414 635000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 632000 317414 635000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 632000 335414 635000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 352794 632000 353414 635000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 370794 632000 371414 635000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 388794 632000 389414 635000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 406794 632000 407414 635000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 424794 632000 425414 635000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 442794 632000 443414 635000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 460794 632000 461414 635000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 478794 632000 479414 635000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 496794 632000 497414 635000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 514794 632000 515414 635000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 532794 632000 533414 635000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 550794 632000 551414 635000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 28794 659000 29414 662000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 46794 659000 47414 662000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 64794 659000 65414 662000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 659000 83414 662000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 659000 101414 662000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 659000 119414 662000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 659000 137414 662000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 659000 155414 662000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 659000 173414 662000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 659000 191414 662000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 659000 209414 662000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 659000 227414 662000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 659000 245414 662000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 659000 263414 662000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 659000 281414 662000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 659000 299414 662000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 659000 317414 662000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 659000 335414 662000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 352794 659000 353414 662000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 370794 659000 371414 662000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 388794 659000 389414 662000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 406794 659000 407414 662000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 424794 659000 425414 662000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 442794 659000 443414 662000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 460794 659000 461414 662000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 478794 659000 479414 662000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 496794 659000 497414 662000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 514794 659000 515414 662000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 532794 659000 533414 662000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 550794 659000 551414 662000 6 vssd1
port 533 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 533 nsew ground input
rlabel metal4 s 10794 -1894 11414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 28794 686000 29414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 46794 686000 47414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 64794 686000 65414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 686000 83414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 686000 101414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 686000 119414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 686000 137414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 686000 155414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 686000 173414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 686000 191414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 686000 209414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 686000 227414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 686000 245414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 686000 263414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 686000 281414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 686000 299414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 686000 317414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 686000 335414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 352794 686000 353414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 370794 686000 371414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 388794 686000 389414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 406794 686000 407414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 424794 686000 425414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 442794 686000 443414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 460794 686000 461414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 478794 686000 479414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 496794 686000 497414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 514794 686000 515414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 532794 686000 533414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 550794 686000 551414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 568794 -1894 569414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 533 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 534 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 535 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 536 nsew signal output
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 537 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 538 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 539 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 540 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 541 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 542 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 543 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 544 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 545 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 546 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 547 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 548 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 549 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 550 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 551 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 552 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 553 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 554 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 555 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 556 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 557 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 558 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 559 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 560 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 561 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 562 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 563 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 564 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 565 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 566 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 567 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 568 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 569 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 570 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 571 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 572 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 573 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 574 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 575 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 576 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 577 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 578 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 579 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 580 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 581 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 582 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 583 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 584 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 585 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 586 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 587 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 588 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 589 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 590 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 591 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 592 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 593 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 594 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 595 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 596 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 597 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 598 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 599 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 600 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 601 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 602 nsew signal output
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 603 nsew signal output
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 604 nsew signal output
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 605 nsew signal output
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 606 nsew signal output
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 607 nsew signal output
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 608 nsew signal output
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 609 nsew signal output
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 610 nsew signal output
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 611 nsew signal output
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 612 nsew signal output
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 613 nsew signal output
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 614 nsew signal output
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 615 nsew signal output
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 616 nsew signal output
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 617 nsew signal output
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 618 nsew signal output
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 619 nsew signal output
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 620 nsew signal output
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 621 nsew signal output
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 622 nsew signal output
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 623 nsew signal output
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 624 nsew signal output
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 625 nsew signal output
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 626 nsew signal output
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 627 nsew signal output
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 628 nsew signal output
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 629 nsew signal output
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 630 nsew signal output
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 631 nsew signal output
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 632 nsew signal output
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 633 nsew signal output
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 634 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 635 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 636 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 637 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 638 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 639 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 5371550
string GDS_FILE /home/matt/work/asic-workshop/shuttle6/tapeout_100/openlane/user_project_wrapper/runs/user_project_wrapper/results/finishing/user_project_wrapper.magic.gds
string GDS_START 1457838
<< end >>

