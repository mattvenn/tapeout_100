* NGSPICE file created from user_project_wrapper.ext - technology: sky130A

* Black-box entry subcircuit for scan_wrapper_lesson_1 abstract view
.subckt scan_wrapper_lesson_1 clk_in clk_out data_in data_out latch_enable_in latch_enable_out
+ scan_select_in scan_select_out vccd1 vssd1
.ends

.subckt user_project_wrapper analog_io[0] analog_io[10] analog_io[11] analog_io[12]
+ analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18]
+ analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23]
+ analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[2]
+ analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7] analog_io[8] analog_io[9]
+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36]
+ io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100]
+ la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105]
+ la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110]
+ la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115]
+ la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120]
+ la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125]
+ la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64]
+ la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6]
+ la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75]
+ la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80]
+ la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86]
+ la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91]
+ la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97]
+ la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101]
+ la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106]
+ la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110]
+ la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115]
+ la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11]
+ la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124]
+ la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33]
+ la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43]
+ la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48]
+ la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63]
+ la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68]
+ la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73]
+ la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78]
+ la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83]
+ la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88]
+ la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93]
+ la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98]
+ la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102]
+ la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109]
+ la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115]
+ la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121]
+ la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12]
+ la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19]
+ la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25]
+ la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31]
+ la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38]
+ la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44]
+ la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50]
+ la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57]
+ la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63]
+ la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6]
+ la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76]
+ la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82]
+ la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89]
+ la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95]
+ la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0]
+ user_irq[1] user_irq[2] vccd1 vssd1 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10]
+ wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16]
+ wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21]
+ wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27]
+ wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3]
+ wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i
+ wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
Xinstance_90 instance_90/clk_in instance_91/clk_in instance_90/data_in instance_91/data_in
+ instance_90/latch_enable_in instance_91/latch_enable_in instance_90/scan_select_in
+ instance_91/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_80 instance_80/clk_in instance_81/clk_in instance_80/data_in instance_81/data_in
+ instance_80/latch_enable_in instance_81/latch_enable_in instance_80/scan_select_in
+ instance_81/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_91 instance_91/clk_in instance_92/clk_in instance_91/data_in instance_92/data_in
+ instance_91/latch_enable_in instance_92/latch_enable_in instance_91/scan_select_in
+ instance_92/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_70 instance_70/clk_in instance_71/clk_in instance_70/data_in instance_71/data_in
+ instance_70/latch_enable_in instance_71/latch_enable_in instance_70/scan_select_in
+ instance_71/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_81 instance_81/clk_in instance_82/clk_in instance_81/data_in instance_82/data_in
+ instance_81/latch_enable_in instance_82/latch_enable_in instance_81/scan_select_in
+ instance_82/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_92 instance_92/clk_in instance_93/clk_in instance_92/data_in instance_93/data_in
+ instance_92/latch_enable_in instance_93/latch_enable_in instance_92/scan_select_in
+ instance_93/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_0 io_in[8] instance_1/clk_in io_in[9] instance_1/data_in io_in[11] instance_1/latch_enable_in
+ io_in[10] instance_1/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_60 instance_60/clk_in instance_61/clk_in instance_60/data_in instance_61/data_in
+ instance_60/latch_enable_in instance_61/latch_enable_in instance_60/scan_select_in
+ instance_61/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_71 instance_71/clk_in instance_72/clk_in instance_71/data_in instance_72/data_in
+ instance_71/latch_enable_in instance_72/latch_enable_in instance_71/scan_select_in
+ instance_72/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_82 instance_82/clk_in instance_83/clk_in instance_82/data_in instance_83/data_in
+ instance_82/latch_enable_in instance_83/latch_enable_in instance_82/scan_select_in
+ instance_83/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_93 instance_93/clk_in instance_94/clk_in instance_93/data_in instance_94/data_in
+ instance_93/latch_enable_in instance_94/latch_enable_in instance_93/scan_select_in
+ instance_94/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_1 instance_1/clk_in instance_2/clk_in instance_1/data_in instance_2/data_in
+ instance_1/latch_enable_in instance_2/latch_enable_in instance_1/scan_select_in
+ instance_2/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_50 instance_50/clk_in instance_51/clk_in instance_50/data_in instance_51/data_in
+ instance_50/latch_enable_in instance_51/latch_enable_in instance_50/scan_select_in
+ instance_51/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_61 instance_61/clk_in instance_62/clk_in instance_61/data_in instance_62/data_in
+ instance_61/latch_enable_in instance_62/latch_enable_in instance_61/scan_select_in
+ instance_62/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_72 instance_72/clk_in instance_73/clk_in instance_72/data_in instance_73/data_in
+ instance_72/latch_enable_in instance_73/latch_enable_in instance_72/scan_select_in
+ instance_73/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_83 instance_83/clk_in instance_84/clk_in instance_83/data_in instance_84/data_in
+ instance_83/latch_enable_in instance_84/latch_enable_in instance_83/scan_select_in
+ instance_84/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_94 instance_94/clk_in instance_95/clk_in instance_94/data_in instance_95/data_in
+ instance_94/latch_enable_in instance_95/latch_enable_in instance_94/scan_select_in
+ instance_95/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_2 instance_2/clk_in instance_3/clk_in instance_2/data_in instance_3/data_in
+ instance_2/latch_enable_in instance_3/latch_enable_in instance_2/scan_select_in
+ instance_3/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_40 instance_40/clk_in instance_41/clk_in instance_40/data_in instance_41/data_in
+ instance_40/latch_enable_in instance_41/latch_enable_in instance_40/scan_select_in
+ instance_41/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_51 instance_51/clk_in instance_52/clk_in instance_51/data_in instance_52/data_in
+ instance_51/latch_enable_in instance_52/latch_enable_in instance_51/scan_select_in
+ instance_52/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_62 instance_62/clk_in instance_63/clk_in instance_62/data_in instance_63/data_in
+ instance_62/latch_enable_in instance_63/latch_enable_in instance_62/scan_select_in
+ instance_63/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_73 instance_73/clk_in instance_74/clk_in instance_73/data_in instance_74/data_in
+ instance_73/latch_enable_in instance_74/latch_enable_in instance_73/scan_select_in
+ instance_74/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_84 instance_84/clk_in instance_85/clk_in instance_84/data_in instance_85/data_in
+ instance_84/latch_enable_in instance_85/latch_enable_in instance_84/scan_select_in
+ instance_85/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_95 instance_95/clk_in instance_96/clk_in instance_95/data_in instance_96/data_in
+ instance_95/latch_enable_in instance_96/latch_enable_in instance_95/scan_select_in
+ instance_96/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_3 instance_3/clk_in instance_4/clk_in instance_3/data_in instance_4/data_in
+ instance_3/latch_enable_in instance_4/latch_enable_in instance_3/scan_select_in
+ instance_4/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_96 instance_96/clk_in instance_97/clk_in instance_96/data_in instance_97/data_in
+ instance_96/latch_enable_in instance_97/latch_enable_in instance_96/scan_select_in
+ instance_97/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_30 instance_30/clk_in instance_31/clk_in instance_30/data_in instance_31/data_in
+ instance_30/latch_enable_in instance_31/latch_enable_in instance_30/scan_select_in
+ instance_31/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_41 instance_41/clk_in instance_42/clk_in instance_41/data_in instance_42/data_in
+ instance_41/latch_enable_in instance_42/latch_enable_in instance_41/scan_select_in
+ instance_42/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_52 instance_52/clk_in instance_53/clk_in instance_52/data_in instance_53/data_in
+ instance_52/latch_enable_in instance_53/latch_enable_in instance_52/scan_select_in
+ instance_53/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_63 instance_63/clk_in instance_64/clk_in instance_63/data_in instance_64/data_in
+ instance_63/latch_enable_in instance_64/latch_enable_in instance_63/scan_select_in
+ instance_64/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_74 instance_74/clk_in instance_75/clk_in instance_74/data_in instance_75/data_in
+ instance_74/latch_enable_in instance_75/latch_enable_in instance_74/scan_select_in
+ instance_75/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_85 instance_85/clk_in instance_86/clk_in instance_85/data_in instance_86/data_in
+ instance_85/latch_enable_in instance_86/latch_enable_in instance_85/scan_select_in
+ instance_86/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_4 instance_4/clk_in instance_5/clk_in instance_4/data_in instance_5/data_in
+ instance_4/latch_enable_in instance_5/latch_enable_in instance_4/scan_select_in
+ instance_5/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_97 instance_97/clk_in instance_98/clk_in instance_97/data_in instance_98/data_in
+ instance_97/latch_enable_in instance_98/latch_enable_in instance_97/scan_select_in
+ instance_98/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_20 instance_20/clk_in instance_21/clk_in instance_20/data_in instance_21/data_in
+ instance_20/latch_enable_in instance_21/latch_enable_in instance_20/scan_select_in
+ instance_21/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_31 instance_31/clk_in instance_32/clk_in instance_31/data_in instance_32/data_in
+ instance_31/latch_enable_in instance_32/latch_enable_in instance_31/scan_select_in
+ instance_32/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_42 instance_42/clk_in instance_43/clk_in instance_42/data_in instance_43/data_in
+ instance_42/latch_enable_in instance_43/latch_enable_in instance_42/scan_select_in
+ instance_43/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_53 instance_53/clk_in instance_54/clk_in instance_53/data_in instance_54/data_in
+ instance_53/latch_enable_in instance_54/latch_enable_in instance_53/scan_select_in
+ instance_54/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_64 instance_64/clk_in instance_65/clk_in instance_64/data_in instance_65/data_in
+ instance_64/latch_enable_in instance_65/latch_enable_in instance_64/scan_select_in
+ instance_65/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_75 instance_75/clk_in instance_76/clk_in instance_75/data_in instance_76/data_in
+ instance_75/latch_enable_in instance_76/latch_enable_in instance_75/scan_select_in
+ instance_76/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_86 instance_86/clk_in instance_87/clk_in instance_86/data_in instance_87/data_in
+ instance_86/latch_enable_in instance_87/latch_enable_in instance_86/scan_select_in
+ instance_87/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_5 instance_5/clk_in instance_6/clk_in instance_5/data_in instance_6/data_in
+ instance_5/latch_enable_in instance_6/latch_enable_in instance_5/scan_select_in
+ instance_6/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_98 instance_98/clk_in instance_99/clk_in instance_98/data_in instance_99/data_in
+ instance_98/latch_enable_in instance_99/latch_enable_in instance_98/scan_select_in
+ instance_99/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_10 instance_9/clk_out instance_11/clk_in instance_9/data_out instance_11/data_in
+ instance_9/latch_enable_out instance_11/latch_enable_in instance_9/scan_select_out
+ instance_11/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_21 instance_21/clk_in instance_22/clk_in instance_21/data_in instance_22/data_in
+ instance_21/latch_enable_in instance_22/latch_enable_in instance_21/scan_select_in
+ instance_22/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_32 instance_32/clk_in instance_33/clk_in instance_32/data_in instance_33/data_in
+ instance_32/latch_enable_in instance_33/latch_enable_in instance_32/scan_select_in
+ instance_33/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_43 instance_43/clk_in instance_44/clk_in instance_43/data_in instance_44/data_in
+ instance_43/latch_enable_in instance_44/latch_enable_in instance_43/scan_select_in
+ instance_44/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_54 instance_54/clk_in instance_55/clk_in instance_54/data_in instance_55/data_in
+ instance_54/latch_enable_in instance_55/latch_enable_in instance_54/scan_select_in
+ instance_55/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_65 instance_65/clk_in instance_66/clk_in instance_65/data_in instance_66/data_in
+ instance_65/latch_enable_in instance_66/latch_enable_in instance_65/scan_select_in
+ instance_66/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_76 instance_76/clk_in instance_77/clk_in instance_76/data_in instance_77/data_in
+ instance_76/latch_enable_in instance_77/latch_enable_in instance_76/scan_select_in
+ instance_77/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_87 instance_87/clk_in instance_88/clk_in instance_87/data_in instance_88/data_in
+ instance_87/latch_enable_in instance_88/latch_enable_in instance_87/scan_select_in
+ instance_88/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_6 instance_6/clk_in instance_7/clk_in instance_6/data_in instance_7/data_in
+ instance_6/latch_enable_in instance_7/latch_enable_in instance_6/scan_select_in
+ instance_7/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_99 instance_99/clk_in instance_99/clk_out instance_99/data_in io_out[11]
+ instance_99/latch_enable_in instance_99/latch_enable_out instance_99/scan_select_in
+ instance_99/scan_select_out vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_11 instance_11/clk_in instance_12/clk_in instance_11/data_in instance_12/data_in
+ instance_11/latch_enable_in instance_12/latch_enable_in instance_11/scan_select_in
+ instance_12/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_22 instance_22/clk_in instance_23/clk_in instance_22/data_in instance_23/data_in
+ instance_22/latch_enable_in instance_23/latch_enable_in instance_22/scan_select_in
+ instance_23/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_33 instance_33/clk_in instance_34/clk_in instance_33/data_in instance_34/data_in
+ instance_33/latch_enable_in instance_34/latch_enable_in instance_33/scan_select_in
+ instance_34/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_44 instance_44/clk_in instance_45/clk_in instance_44/data_in instance_45/data_in
+ instance_44/latch_enable_in instance_45/latch_enable_in instance_44/scan_select_in
+ instance_45/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_55 instance_55/clk_in instance_56/clk_in instance_55/data_in instance_56/data_in
+ instance_55/latch_enable_in instance_56/latch_enable_in instance_55/scan_select_in
+ instance_56/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_66 instance_66/clk_in instance_67/clk_in instance_66/data_in instance_67/data_in
+ instance_66/latch_enable_in instance_67/latch_enable_in instance_66/scan_select_in
+ instance_67/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_77 instance_77/clk_in instance_78/clk_in instance_77/data_in instance_78/data_in
+ instance_77/latch_enable_in instance_78/latch_enable_in instance_77/scan_select_in
+ instance_78/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_88 instance_88/clk_in instance_89/clk_in instance_88/data_in instance_89/data_in
+ instance_88/latch_enable_in instance_89/latch_enable_in instance_88/scan_select_in
+ instance_89/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_7 instance_7/clk_in instance_8/clk_in instance_7/data_in instance_8/data_in
+ instance_7/latch_enable_in instance_8/latch_enable_in instance_7/scan_select_in
+ instance_8/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_12 instance_12/clk_in instance_13/clk_in instance_12/data_in instance_13/data_in
+ instance_12/latch_enable_in instance_13/latch_enable_in instance_12/scan_select_in
+ instance_13/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_23 instance_23/clk_in instance_24/clk_in instance_23/data_in instance_24/data_in
+ instance_23/latch_enable_in instance_24/latch_enable_in instance_23/scan_select_in
+ instance_24/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_34 instance_34/clk_in instance_35/clk_in instance_34/data_in instance_35/data_in
+ instance_34/latch_enable_in instance_35/latch_enable_in instance_34/scan_select_in
+ instance_35/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_45 instance_45/clk_in instance_46/clk_in instance_45/data_in instance_46/data_in
+ instance_45/latch_enable_in instance_46/latch_enable_in instance_45/scan_select_in
+ instance_46/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_56 instance_56/clk_in instance_57/clk_in instance_56/data_in instance_57/data_in
+ instance_56/latch_enable_in instance_57/latch_enable_in instance_56/scan_select_in
+ instance_57/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_67 instance_67/clk_in instance_68/clk_in instance_67/data_in instance_68/data_in
+ instance_67/latch_enable_in instance_68/latch_enable_in instance_67/scan_select_in
+ instance_68/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_78 instance_78/clk_in instance_79/clk_in instance_78/data_in instance_79/data_in
+ instance_78/latch_enable_in instance_79/latch_enable_in instance_78/scan_select_in
+ instance_79/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_89 instance_89/clk_in instance_90/clk_in instance_89/data_in instance_90/data_in
+ instance_89/latch_enable_in instance_90/latch_enable_in instance_89/scan_select_in
+ instance_90/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_8 instance_8/clk_in instance_9/clk_in instance_8/data_in instance_9/data_in
+ instance_8/latch_enable_in instance_9/latch_enable_in instance_8/scan_select_in
+ instance_9/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_13 instance_13/clk_in instance_14/clk_in instance_13/data_in instance_14/data_in
+ instance_13/latch_enable_in instance_14/latch_enable_in instance_13/scan_select_in
+ instance_14/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_24 instance_24/clk_in instance_25/clk_in instance_24/data_in instance_25/data_in
+ instance_24/latch_enable_in instance_25/latch_enable_in instance_24/scan_select_in
+ instance_25/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_35 instance_35/clk_in instance_36/clk_in instance_35/data_in instance_36/data_in
+ instance_35/latch_enable_in instance_36/latch_enable_in instance_35/scan_select_in
+ instance_36/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_46 instance_46/clk_in instance_47/clk_in instance_46/data_in instance_47/data_in
+ instance_46/latch_enable_in instance_47/latch_enable_in instance_46/scan_select_in
+ instance_47/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_57 instance_57/clk_in instance_58/clk_in instance_57/data_in instance_58/data_in
+ instance_57/latch_enable_in instance_58/latch_enable_in instance_57/scan_select_in
+ instance_58/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_68 instance_68/clk_in instance_69/clk_in instance_68/data_in instance_69/data_in
+ instance_68/latch_enable_in instance_69/latch_enable_in instance_68/scan_select_in
+ instance_69/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_79 instance_79/clk_in instance_80/clk_in instance_79/data_in instance_80/data_in
+ instance_79/latch_enable_in instance_80/latch_enable_in instance_79/scan_select_in
+ instance_80/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_9 instance_9/clk_in instance_9/clk_out instance_9/data_in instance_9/data_out
+ instance_9/latch_enable_in instance_9/latch_enable_out instance_9/scan_select_in
+ instance_9/scan_select_out vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_14 instance_14/clk_in instance_15/clk_in instance_14/data_in instance_15/data_in
+ instance_14/latch_enable_in instance_15/latch_enable_in instance_14/scan_select_in
+ instance_15/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_25 instance_25/clk_in instance_26/clk_in instance_25/data_in instance_26/data_in
+ instance_25/latch_enable_in instance_26/latch_enable_in instance_25/scan_select_in
+ instance_26/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_36 instance_36/clk_in instance_37/clk_in instance_36/data_in instance_37/data_in
+ instance_36/latch_enable_in instance_37/latch_enable_in instance_36/scan_select_in
+ instance_37/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_47 instance_47/clk_in instance_48/clk_in instance_47/data_in instance_48/data_in
+ instance_47/latch_enable_in instance_48/latch_enable_in instance_47/scan_select_in
+ instance_48/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_58 instance_58/clk_in instance_59/clk_in instance_58/data_in instance_59/data_in
+ instance_58/latch_enable_in instance_59/latch_enable_in instance_58/scan_select_in
+ instance_59/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_69 instance_69/clk_in instance_70/clk_in instance_69/data_in instance_70/data_in
+ instance_69/latch_enable_in instance_70/latch_enable_in instance_69/scan_select_in
+ instance_70/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_15 instance_15/clk_in instance_16/clk_in instance_15/data_in instance_16/data_in
+ instance_15/latch_enable_in instance_16/latch_enable_in instance_15/scan_select_in
+ instance_16/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_26 instance_26/clk_in instance_27/clk_in instance_26/data_in instance_27/data_in
+ instance_26/latch_enable_in instance_27/latch_enable_in instance_26/scan_select_in
+ instance_27/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_37 instance_37/clk_in instance_38/clk_in instance_37/data_in instance_38/data_in
+ instance_37/latch_enable_in instance_38/latch_enable_in instance_37/scan_select_in
+ instance_38/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_48 instance_48/clk_in instance_49/clk_in instance_48/data_in instance_49/data_in
+ instance_48/latch_enable_in instance_49/latch_enable_in instance_48/scan_select_in
+ instance_49/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_59 instance_59/clk_in instance_60/clk_in instance_59/data_in instance_60/data_in
+ instance_59/latch_enable_in instance_60/latch_enable_in instance_59/scan_select_in
+ instance_60/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_16 instance_16/clk_in instance_17/clk_in instance_16/data_in instance_17/data_in
+ instance_16/latch_enable_in instance_17/latch_enable_in instance_16/scan_select_in
+ instance_17/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_27 instance_27/clk_in instance_28/clk_in instance_27/data_in instance_28/data_in
+ instance_27/latch_enable_in instance_28/latch_enable_in instance_27/scan_select_in
+ instance_28/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_38 instance_38/clk_in instance_39/clk_in instance_38/data_in instance_39/data_in
+ instance_38/latch_enable_in instance_39/latch_enable_in instance_38/scan_select_in
+ instance_39/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_49 instance_49/clk_in instance_50/clk_in instance_49/data_in instance_50/data_in
+ instance_49/latch_enable_in instance_50/latch_enable_in instance_49/scan_select_in
+ instance_50/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_17 instance_17/clk_in instance_18/clk_in instance_17/data_in instance_18/data_in
+ instance_17/latch_enable_in instance_18/latch_enable_in instance_17/scan_select_in
+ instance_18/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_28 instance_28/clk_in instance_29/clk_in instance_28/data_in instance_29/data_in
+ instance_28/latch_enable_in instance_29/latch_enable_in instance_28/scan_select_in
+ instance_29/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_39 instance_39/clk_in instance_40/clk_in instance_39/data_in instance_40/data_in
+ instance_39/latch_enable_in instance_40/latch_enable_in instance_39/scan_select_in
+ instance_40/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_18 instance_18/clk_in instance_19/clk_in instance_18/data_in instance_19/data_in
+ instance_18/latch_enable_in instance_19/latch_enable_in instance_18/scan_select_in
+ instance_19/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_29 instance_29/clk_in instance_30/clk_in instance_29/data_in instance_30/data_in
+ instance_29/latch_enable_in instance_30/latch_enable_in instance_29/scan_select_in
+ instance_30/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_19 instance_19/clk_in instance_20/clk_in instance_19/data_in instance_20/data_in
+ instance_19/latch_enable_in instance_20/latch_enable_in instance_19/scan_select_in
+ instance_20/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
.ends

