VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO scan_wrapper_lesson_1
  CLASS BLOCK ;
  FOREIGN scan_wrapper_lesson_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 70.000 BY 70.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.540 4.000 58.740 ;
    END
  END clk
  PIN data_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -0.050 0.000 0.510 4.000 ;
    END
  END data_in
  PIN data_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 66.000 40.540 70.000 41.740 ;
    END
  END data_out
  PIN latch_enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.810 66.000 42.370 70.000 ;
    END
  END latch_enable
  PIN scan_select
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.690 0.000 55.250 4.000 ;
    END
  END scan_select
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 14.550 10.640 16.150 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 34.200 10.640 35.800 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 53.855 10.640 55.455 57.360 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.370 10.640 25.970 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 44.025 10.640 45.625 57.360 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 64.400 57.205 ;
      LAYER met1 ;
        RECT 0.070 10.640 64.400 57.360 ;
      LAYER met2 ;
        RECT 0.100 65.720 41.530 66.000 ;
        RECT 42.650 65.720 61.080 66.000 ;
        RECT 0.100 4.280 61.080 65.720 ;
        RECT 0.790 4.000 54.410 4.280 ;
        RECT 55.530 4.000 61.080 4.280 ;
      LAYER met3 ;
        RECT 4.400 57.140 66.000 58.305 ;
        RECT 4.000 42.140 66.000 57.140 ;
        RECT 4.000 40.140 65.600 42.140 ;
        RECT 4.000 10.715 66.000 40.140 ;
      LAYER met4 ;
        RECT 16.550 10.640 23.970 57.360 ;
        RECT 26.370 10.640 33.800 57.360 ;
        RECT 36.200 10.640 43.625 57.360 ;
        RECT 46.025 10.640 53.455 57.360 ;
  END
END scan_wrapper_lesson_1
END LIBRARY

