* NGSPICE file created from user_project_wrapper.ext - technology: sky130A

* Black-box entry subcircuit for scan_wrapper_lesson_1 abstract view
.subckt scan_wrapper_lesson_1 clk_in clk_out data_in data_out latch_enable_in latch_enable_out
+ scan_select_in scan_select_out vccd1 vssd1
.ends

.subckt user_project_wrapper analog_io[0] analog_io[10] analog_io[11] analog_io[12]
+ analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18]
+ analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23]
+ analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[2]
+ analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7] analog_io[8] analog_io[9]
+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36]
+ io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100]
+ la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105]
+ la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110]
+ la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115]
+ la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120]
+ la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125]
+ la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64]
+ la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6]
+ la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75]
+ la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80]
+ la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86]
+ la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91]
+ la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97]
+ la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101]
+ la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106]
+ la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110]
+ la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115]
+ la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11]
+ la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124]
+ la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33]
+ la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43]
+ la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48]
+ la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63]
+ la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68]
+ la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73]
+ la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78]
+ la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83]
+ la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88]
+ la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93]
+ la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98]
+ la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102]
+ la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109]
+ la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115]
+ la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121]
+ la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12]
+ la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19]
+ la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25]
+ la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31]
+ la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38]
+ la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44]
+ la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50]
+ la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57]
+ la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63]
+ la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6]
+ la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76]
+ la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82]
+ la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89]
+ la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95]
+ la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0]
+ user_irq[1] user_irq[2] vccd1 vssd1 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10]
+ wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16]
+ wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21]
+ wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27]
+ wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3]
+ wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i
+ wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
Xinstance_389 instance_389/clk_in instance_390/clk_in instance_389/data_in instance_390/data_in
+ instance_389/latch_enable_in instance_390/latch_enable_in instance_389/scan_select_in
+ instance_390/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_301 instance_301/clk_in instance_302/clk_in instance_301/data_in instance_302/data_in
+ instance_301/latch_enable_in instance_302/latch_enable_in instance_301/scan_select_in
+ instance_302/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_312 instance_312/clk_in instance_313/clk_in instance_312/data_in instance_313/data_in
+ instance_312/latch_enable_in instance_313/latch_enable_in instance_312/scan_select_in
+ instance_313/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_323 instance_323/clk_in instance_324/clk_in instance_323/data_in instance_324/data_in
+ instance_323/latch_enable_in instance_324/latch_enable_in instance_323/scan_select_in
+ instance_324/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_334 instance_334/clk_in instance_335/clk_in instance_334/data_in instance_335/data_in
+ instance_334/latch_enable_in instance_335/latch_enable_in instance_334/scan_select_in
+ instance_335/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_345 instance_345/clk_in instance_346/clk_in instance_345/data_in instance_346/data_in
+ instance_345/latch_enable_in instance_346/latch_enable_in instance_345/scan_select_in
+ instance_346/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_356 instance_356/clk_in instance_357/clk_in instance_356/data_in instance_357/data_in
+ instance_356/latch_enable_in instance_357/latch_enable_in instance_356/scan_select_in
+ instance_357/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_367 instance_367/clk_in instance_368/clk_in instance_367/data_in instance_368/data_in
+ instance_367/latch_enable_in instance_368/latch_enable_in instance_367/scan_select_in
+ instance_368/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_378 instance_378/clk_in instance_379/clk_in instance_378/data_in instance_379/data_in
+ instance_378/latch_enable_in instance_379/latch_enable_in instance_378/scan_select_in
+ instance_379/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_120 instance_120/clk_in instance_121/clk_in instance_120/data_in instance_121/data_in
+ instance_120/latch_enable_in instance_121/latch_enable_in instance_120/scan_select_in
+ instance_121/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_131 instance_131/clk_in instance_132/clk_in instance_131/data_in instance_132/data_in
+ instance_131/latch_enable_in instance_132/latch_enable_in instance_131/scan_select_in
+ instance_132/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_142 instance_142/clk_in instance_143/clk_in instance_142/data_in instance_143/data_in
+ instance_142/latch_enable_in instance_143/latch_enable_in instance_142/scan_select_in
+ instance_143/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_153 instance_153/clk_in instance_154/clk_in instance_153/data_in instance_154/data_in
+ instance_153/latch_enable_in instance_154/latch_enable_in instance_153/scan_select_in
+ instance_154/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_164 instance_164/clk_in instance_165/clk_in instance_164/data_in instance_165/data_in
+ instance_164/latch_enable_in instance_165/latch_enable_in instance_164/scan_select_in
+ instance_165/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_175 instance_175/clk_in instance_176/clk_in instance_175/data_in instance_176/data_in
+ instance_175/latch_enable_in instance_176/latch_enable_in instance_175/scan_select_in
+ instance_176/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_186 instance_186/clk_in instance_187/clk_in instance_186/data_in instance_187/data_in
+ instance_186/latch_enable_in instance_187/latch_enable_in instance_186/scan_select_in
+ instance_187/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_197 instance_197/clk_in instance_198/clk_in instance_197/data_in instance_198/data_in
+ instance_197/latch_enable_in instance_198/latch_enable_in instance_197/scan_select_in
+ instance_198/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_302 instance_302/clk_in instance_303/clk_in instance_302/data_in instance_303/data_in
+ instance_302/latch_enable_in instance_303/latch_enable_in instance_302/scan_select_in
+ instance_303/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_313 instance_313/clk_in instance_314/clk_in instance_313/data_in instance_314/data_in
+ instance_313/latch_enable_in instance_314/latch_enable_in instance_313/scan_select_in
+ instance_314/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_324 instance_324/clk_in instance_325/clk_in instance_324/data_in instance_325/data_in
+ instance_324/latch_enable_in instance_325/latch_enable_in instance_324/scan_select_in
+ instance_325/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_335 instance_335/clk_in instance_336/clk_in instance_335/data_in instance_336/data_in
+ instance_335/latch_enable_in instance_336/latch_enable_in instance_335/scan_select_in
+ instance_336/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_346 instance_346/clk_in instance_347/clk_in instance_346/data_in instance_347/data_in
+ instance_346/latch_enable_in instance_347/latch_enable_in instance_346/scan_select_in
+ instance_347/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_357 instance_357/clk_in instance_358/clk_in instance_357/data_in instance_358/data_in
+ instance_357/latch_enable_in instance_358/latch_enable_in instance_357/scan_select_in
+ instance_358/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_368 instance_368/clk_in instance_369/clk_in instance_368/data_in instance_369/data_in
+ instance_368/latch_enable_in instance_369/latch_enable_in instance_368/scan_select_in
+ instance_369/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_379 instance_379/clk_in instance_380/clk_in instance_379/data_in instance_380/data_in
+ instance_379/latch_enable_in instance_380/latch_enable_in instance_379/scan_select_in
+ instance_380/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_110 instance_110/clk_in instance_111/clk_in instance_110/data_in instance_111/data_in
+ instance_110/latch_enable_in instance_111/latch_enable_in instance_110/scan_select_in
+ instance_111/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_121 instance_121/clk_in instance_122/clk_in instance_121/data_in instance_122/data_in
+ instance_121/latch_enable_in instance_122/latch_enable_in instance_121/scan_select_in
+ instance_122/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_132 instance_132/clk_in instance_133/clk_in instance_132/data_in instance_133/data_in
+ instance_132/latch_enable_in instance_133/latch_enable_in instance_132/scan_select_in
+ instance_133/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_143 instance_143/clk_in instance_144/clk_in instance_143/data_in instance_144/data_in
+ instance_143/latch_enable_in instance_144/latch_enable_in instance_143/scan_select_in
+ instance_144/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_154 instance_154/clk_in instance_155/clk_in instance_154/data_in instance_155/data_in
+ instance_154/latch_enable_in instance_155/latch_enable_in instance_154/scan_select_in
+ instance_155/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_165 instance_165/clk_in instance_166/clk_in instance_165/data_in instance_166/data_in
+ instance_165/latch_enable_in instance_166/latch_enable_in instance_165/scan_select_in
+ instance_166/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_176 instance_176/clk_in instance_177/clk_in instance_176/data_in instance_177/data_in
+ instance_176/latch_enable_in instance_177/latch_enable_in instance_176/scan_select_in
+ instance_177/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_187 instance_187/clk_in instance_188/clk_in instance_187/data_in instance_188/data_in
+ instance_187/latch_enable_in instance_188/latch_enable_in instance_187/scan_select_in
+ instance_188/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_198 instance_198/clk_in instance_199/clk_in instance_198/data_in instance_199/data_in
+ instance_198/latch_enable_in instance_199/latch_enable_in instance_198/scan_select_in
+ instance_199/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_303 instance_303/clk_in instance_304/clk_in instance_303/data_in instance_304/data_in
+ instance_303/latch_enable_in instance_304/latch_enable_in instance_303/scan_select_in
+ instance_304/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_314 instance_314/clk_in instance_315/clk_in instance_314/data_in instance_315/data_in
+ instance_314/latch_enable_in instance_315/latch_enable_in instance_314/scan_select_in
+ instance_315/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_325 instance_325/clk_in instance_326/clk_in instance_325/data_in instance_326/data_in
+ instance_325/latch_enable_in instance_326/latch_enable_in instance_325/scan_select_in
+ instance_326/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_336 instance_336/clk_in instance_337/clk_in instance_336/data_in instance_337/data_in
+ instance_336/latch_enable_in instance_337/latch_enable_in instance_336/scan_select_in
+ instance_337/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_347 instance_347/clk_in instance_348/clk_in instance_347/data_in instance_348/data_in
+ instance_347/latch_enable_in instance_348/latch_enable_in instance_347/scan_select_in
+ instance_348/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_358 instance_358/clk_in instance_359/clk_in instance_358/data_in instance_359/data_in
+ instance_358/latch_enable_in instance_359/latch_enable_in instance_358/scan_select_in
+ instance_359/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_369 instance_369/clk_in instance_370/clk_in instance_369/data_in instance_370/data_in
+ instance_369/latch_enable_in instance_370/latch_enable_in instance_369/scan_select_in
+ instance_370/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_100 instance_99/clk_out instance_101/clk_in instance_99/data_out instance_101/data_in
+ instance_99/latch_enable_out instance_101/latch_enable_in instance_99/scan_select_out
+ instance_101/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_111 instance_111/clk_in instance_112/clk_in instance_111/data_in instance_112/data_in
+ instance_111/latch_enable_in instance_112/latch_enable_in instance_111/scan_select_in
+ instance_112/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_122 instance_122/clk_in instance_123/clk_in instance_122/data_in instance_123/data_in
+ instance_122/latch_enable_in instance_123/latch_enable_in instance_122/scan_select_in
+ instance_123/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_133 instance_133/clk_in instance_134/clk_in instance_133/data_in instance_134/data_in
+ instance_133/latch_enable_in instance_134/latch_enable_in instance_133/scan_select_in
+ instance_134/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_144 instance_144/clk_in instance_145/clk_in instance_144/data_in instance_145/data_in
+ instance_144/latch_enable_in instance_145/latch_enable_in instance_144/scan_select_in
+ instance_145/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_155 instance_155/clk_in instance_156/clk_in instance_155/data_in instance_156/data_in
+ instance_155/latch_enable_in instance_156/latch_enable_in instance_155/scan_select_in
+ instance_156/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_166 instance_166/clk_in instance_167/clk_in instance_166/data_in instance_167/data_in
+ instance_166/latch_enable_in instance_167/latch_enable_in instance_166/scan_select_in
+ instance_167/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_177 instance_177/clk_in instance_178/clk_in instance_177/data_in instance_178/data_in
+ instance_177/latch_enable_in instance_178/latch_enable_in instance_177/scan_select_in
+ instance_178/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_188 instance_188/clk_in instance_189/clk_in instance_188/data_in instance_189/data_in
+ instance_188/latch_enable_in instance_189/latch_enable_in instance_188/scan_select_in
+ instance_189/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_199 instance_199/clk_in instance_200/clk_in instance_199/data_in instance_200/data_in
+ instance_199/latch_enable_in instance_200/latch_enable_in instance_199/scan_select_in
+ instance_200/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_304 instance_304/clk_in instance_305/clk_in instance_304/data_in instance_305/data_in
+ instance_304/latch_enable_in instance_305/latch_enable_in instance_304/scan_select_in
+ instance_305/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_315 instance_315/clk_in instance_316/clk_in instance_315/data_in instance_316/data_in
+ instance_315/latch_enable_in instance_316/latch_enable_in instance_315/scan_select_in
+ instance_316/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_326 instance_326/clk_in instance_327/clk_in instance_326/data_in instance_327/data_in
+ instance_326/latch_enable_in instance_327/latch_enable_in instance_326/scan_select_in
+ instance_327/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_337 instance_337/clk_in instance_338/clk_in instance_337/data_in instance_338/data_in
+ instance_337/latch_enable_in instance_338/latch_enable_in instance_337/scan_select_in
+ instance_338/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_348 instance_348/clk_in instance_349/clk_in instance_348/data_in instance_349/data_in
+ instance_348/latch_enable_in instance_349/latch_enable_in instance_348/scan_select_in
+ instance_349/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_359 instance_359/clk_in instance_360/clk_in instance_359/data_in instance_360/data_in
+ instance_359/latch_enable_in instance_360/latch_enable_in instance_359/scan_select_in
+ instance_360/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_101 instance_101/clk_in instance_102/clk_in instance_101/data_in instance_102/data_in
+ instance_101/latch_enable_in instance_102/latch_enable_in instance_101/scan_select_in
+ instance_102/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_112 instance_112/clk_in instance_113/clk_in instance_112/data_in instance_113/data_in
+ instance_112/latch_enable_in instance_113/latch_enable_in instance_112/scan_select_in
+ instance_113/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_123 instance_123/clk_in instance_124/clk_in instance_123/data_in instance_124/data_in
+ instance_123/latch_enable_in instance_124/latch_enable_in instance_123/scan_select_in
+ instance_124/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_134 instance_134/clk_in instance_135/clk_in instance_134/data_in instance_135/data_in
+ instance_134/latch_enable_in instance_135/latch_enable_in instance_134/scan_select_in
+ instance_135/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_145 instance_145/clk_in instance_146/clk_in instance_145/data_in instance_146/data_in
+ instance_145/latch_enable_in instance_146/latch_enable_in instance_145/scan_select_in
+ instance_146/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_156 instance_156/clk_in instance_157/clk_in instance_156/data_in instance_157/data_in
+ instance_156/latch_enable_in instance_157/latch_enable_in instance_156/scan_select_in
+ instance_157/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_167 instance_167/clk_in instance_168/clk_in instance_167/data_in instance_168/data_in
+ instance_167/latch_enable_in instance_168/latch_enable_in instance_167/scan_select_in
+ instance_168/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_178 instance_178/clk_in instance_179/clk_in instance_178/data_in instance_179/data_in
+ instance_178/latch_enable_in instance_179/latch_enable_in instance_178/scan_select_in
+ instance_179/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_189 instance_189/clk_in instance_190/clk_in instance_189/data_in instance_190/data_in
+ instance_189/latch_enable_in instance_190/latch_enable_in instance_189/scan_select_in
+ instance_190/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_305 instance_305/clk_in instance_306/clk_in instance_305/data_in instance_306/data_in
+ instance_305/latch_enable_in instance_306/latch_enable_in instance_305/scan_select_in
+ instance_306/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_316 instance_316/clk_in instance_317/clk_in instance_316/data_in instance_317/data_in
+ instance_316/latch_enable_in instance_317/latch_enable_in instance_316/scan_select_in
+ instance_317/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_327 instance_327/clk_in instance_328/clk_in instance_327/data_in instance_328/data_in
+ instance_327/latch_enable_in instance_328/latch_enable_in instance_327/scan_select_in
+ instance_328/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_338 instance_338/clk_in instance_339/clk_in instance_338/data_in instance_339/data_in
+ instance_338/latch_enable_in instance_339/latch_enable_in instance_338/scan_select_in
+ instance_339/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_349 instance_349/clk_in instance_350/clk_in instance_349/data_in instance_350/data_in
+ instance_349/latch_enable_in instance_350/latch_enable_in instance_349/scan_select_in
+ instance_350/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_102 instance_102/clk_in instance_103/clk_in instance_102/data_in instance_103/data_in
+ instance_102/latch_enable_in instance_103/latch_enable_in instance_102/scan_select_in
+ instance_103/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_113 instance_113/clk_in instance_114/clk_in instance_113/data_in instance_114/data_in
+ instance_113/latch_enable_in instance_114/latch_enable_in instance_113/scan_select_in
+ instance_114/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_124 instance_124/clk_in instance_125/clk_in instance_124/data_in instance_125/data_in
+ instance_124/latch_enable_in instance_125/latch_enable_in instance_124/scan_select_in
+ instance_125/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_135 instance_135/clk_in instance_136/clk_in instance_135/data_in instance_136/data_in
+ instance_135/latch_enable_in instance_136/latch_enable_in instance_135/scan_select_in
+ instance_136/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_146 instance_146/clk_in instance_147/clk_in instance_146/data_in instance_147/data_in
+ instance_146/latch_enable_in instance_147/latch_enable_in instance_146/scan_select_in
+ instance_147/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_157 instance_157/clk_in instance_158/clk_in instance_157/data_in instance_158/data_in
+ instance_157/latch_enable_in instance_158/latch_enable_in instance_157/scan_select_in
+ instance_158/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_168 instance_168/clk_in instance_169/clk_in instance_168/data_in instance_169/data_in
+ instance_168/latch_enable_in instance_169/latch_enable_in instance_168/scan_select_in
+ instance_169/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_179 instance_179/clk_in instance_180/clk_in instance_179/data_in instance_180/data_in
+ instance_179/latch_enable_in instance_180/latch_enable_in instance_179/scan_select_in
+ instance_180/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_306 instance_306/clk_in instance_307/clk_in instance_306/data_in instance_307/data_in
+ instance_306/latch_enable_in instance_307/latch_enable_in instance_306/scan_select_in
+ instance_307/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_317 instance_317/clk_in instance_318/clk_in instance_317/data_in instance_318/data_in
+ instance_317/latch_enable_in instance_318/latch_enable_in instance_317/scan_select_in
+ instance_318/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_328 instance_328/clk_in instance_329/clk_in instance_328/data_in instance_329/data_in
+ instance_328/latch_enable_in instance_329/latch_enable_in instance_328/scan_select_in
+ instance_329/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_339 instance_339/clk_in instance_340/clk_in instance_339/data_in instance_340/data_in
+ instance_339/latch_enable_in instance_340/latch_enable_in instance_339/scan_select_in
+ instance_340/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_103 instance_103/clk_in instance_104/clk_in instance_103/data_in instance_104/data_in
+ instance_103/latch_enable_in instance_104/latch_enable_in instance_103/scan_select_in
+ instance_104/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_114 instance_114/clk_in instance_115/clk_in instance_114/data_in instance_115/data_in
+ instance_114/latch_enable_in instance_115/latch_enable_in instance_114/scan_select_in
+ instance_115/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_125 instance_125/clk_in instance_126/clk_in instance_125/data_in instance_126/data_in
+ instance_125/latch_enable_in instance_126/latch_enable_in instance_125/scan_select_in
+ instance_126/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_136 instance_136/clk_in instance_137/clk_in instance_136/data_in instance_137/data_in
+ instance_136/latch_enable_in instance_137/latch_enable_in instance_136/scan_select_in
+ instance_137/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_147 instance_147/clk_in instance_148/clk_in instance_147/data_in instance_148/data_in
+ instance_147/latch_enable_in instance_148/latch_enable_in instance_147/scan_select_in
+ instance_148/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_158 instance_158/clk_in instance_159/clk_in instance_158/data_in instance_159/data_in
+ instance_158/latch_enable_in instance_159/latch_enable_in instance_158/scan_select_in
+ instance_159/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_169 instance_169/clk_in instance_170/clk_in instance_169/data_in instance_170/data_in
+ instance_169/latch_enable_in instance_170/latch_enable_in instance_169/scan_select_in
+ instance_170/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_307 instance_307/clk_in instance_308/clk_in instance_307/data_in instance_308/data_in
+ instance_307/latch_enable_in instance_308/latch_enable_in instance_307/scan_select_in
+ instance_308/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_318 instance_318/clk_in instance_319/clk_in instance_318/data_in instance_319/data_in
+ instance_318/latch_enable_in instance_319/latch_enable_in instance_318/scan_select_in
+ instance_319/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_329 instance_329/clk_in instance_330/clk_in instance_329/data_in instance_330/data_in
+ instance_329/latch_enable_in instance_330/latch_enable_in instance_329/scan_select_in
+ instance_330/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_104 instance_104/clk_in instance_105/clk_in instance_104/data_in instance_105/data_in
+ instance_104/latch_enable_in instance_105/latch_enable_in instance_104/scan_select_in
+ instance_105/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_115 instance_115/clk_in instance_116/clk_in instance_115/data_in instance_116/data_in
+ instance_115/latch_enable_in instance_116/latch_enable_in instance_115/scan_select_in
+ instance_116/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_126 instance_126/clk_in instance_127/clk_in instance_126/data_in instance_127/data_in
+ instance_126/latch_enable_in instance_127/latch_enable_in instance_126/scan_select_in
+ instance_127/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_137 instance_137/clk_in instance_138/clk_in instance_137/data_in instance_138/data_in
+ instance_137/latch_enable_in instance_138/latch_enable_in instance_137/scan_select_in
+ instance_138/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_148 instance_148/clk_in instance_149/clk_in instance_148/data_in instance_149/data_in
+ instance_148/latch_enable_in instance_149/latch_enable_in instance_148/scan_select_in
+ instance_149/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_159 instance_159/clk_in instance_160/clk_in instance_159/data_in instance_160/data_in
+ instance_159/latch_enable_in instance_160/latch_enable_in instance_159/scan_select_in
+ instance_160/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_308 instance_308/clk_in instance_309/clk_in instance_308/data_in instance_309/data_in
+ instance_308/latch_enable_in instance_309/latch_enable_in instance_308/scan_select_in
+ instance_309/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_319 instance_319/clk_in instance_320/clk_in instance_319/data_in instance_320/data_in
+ instance_319/latch_enable_in instance_320/latch_enable_in instance_319/scan_select_in
+ instance_320/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_105 instance_105/clk_in instance_106/clk_in instance_105/data_in instance_106/data_in
+ instance_105/latch_enable_in instance_106/latch_enable_in instance_105/scan_select_in
+ instance_106/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_116 instance_116/clk_in instance_117/clk_in instance_116/data_in instance_117/data_in
+ instance_116/latch_enable_in instance_117/latch_enable_in instance_116/scan_select_in
+ instance_117/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_127 instance_127/clk_in instance_128/clk_in instance_127/data_in instance_128/data_in
+ instance_127/latch_enable_in instance_128/latch_enable_in instance_127/scan_select_in
+ instance_128/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_138 instance_138/clk_in instance_139/clk_in instance_138/data_in instance_139/data_in
+ instance_138/latch_enable_in instance_139/latch_enable_in instance_138/scan_select_in
+ instance_139/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_149 instance_149/clk_in instance_150/clk_in instance_149/data_in instance_150/data_in
+ instance_149/latch_enable_in instance_150/latch_enable_in instance_149/scan_select_in
+ instance_150/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_309 instance_309/clk_in instance_310/clk_in instance_309/data_in instance_310/data_in
+ instance_309/latch_enable_in instance_310/latch_enable_in instance_309/scan_select_in
+ instance_310/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_106 instance_106/clk_in instance_107/clk_in instance_106/data_in instance_107/data_in
+ instance_106/latch_enable_in instance_107/latch_enable_in instance_106/scan_select_in
+ instance_107/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_117 instance_117/clk_in instance_118/clk_in instance_117/data_in instance_118/data_in
+ instance_117/latch_enable_in instance_118/latch_enable_in instance_117/scan_select_in
+ instance_118/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_128 instance_128/clk_in instance_129/clk_in instance_128/data_in instance_129/data_in
+ instance_128/latch_enable_in instance_129/latch_enable_in instance_128/scan_select_in
+ instance_129/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_139 instance_139/clk_in instance_140/clk_in instance_139/data_in instance_140/data_in
+ instance_139/latch_enable_in instance_140/latch_enable_in instance_139/scan_select_in
+ instance_140/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_107 instance_107/clk_in instance_108/clk_in instance_107/data_in instance_108/data_in
+ instance_107/latch_enable_in instance_108/latch_enable_in instance_107/scan_select_in
+ instance_108/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_118 instance_118/clk_in instance_119/clk_in instance_118/data_in instance_119/data_in
+ instance_118/latch_enable_in instance_119/latch_enable_in instance_118/scan_select_in
+ instance_119/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_129 instance_129/clk_in instance_130/clk_in instance_129/data_in instance_130/data_in
+ instance_129/latch_enable_in instance_130/latch_enable_in instance_129/scan_select_in
+ instance_130/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_290 instance_290/clk_in instance_291/clk_in instance_290/data_in instance_291/data_in
+ instance_290/latch_enable_in instance_291/latch_enable_in instance_290/scan_select_in
+ instance_291/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_108 instance_108/clk_in instance_109/clk_in instance_108/data_in instance_109/data_in
+ instance_108/latch_enable_in instance_109/latch_enable_in instance_108/scan_select_in
+ instance_109/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_119 instance_119/clk_in instance_120/clk_in instance_119/data_in instance_120/data_in
+ instance_119/latch_enable_in instance_120/latch_enable_in instance_119/scan_select_in
+ instance_120/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_280 instance_280/clk_in instance_281/clk_in instance_280/data_in instance_281/data_in
+ instance_280/latch_enable_in instance_281/latch_enable_in instance_280/scan_select_in
+ instance_281/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_291 instance_291/clk_in instance_292/clk_in instance_291/data_in instance_292/data_in
+ instance_291/latch_enable_in instance_292/latch_enable_in instance_291/scan_select_in
+ instance_292/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_109 instance_109/clk_in instance_110/clk_in instance_109/data_in instance_110/data_in
+ instance_109/latch_enable_in instance_110/latch_enable_in instance_109/scan_select_in
+ instance_110/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_270 instance_270/clk_in instance_271/clk_in instance_270/data_in instance_271/data_in
+ instance_270/latch_enable_in instance_271/latch_enable_in instance_270/scan_select_in
+ instance_271/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_281 instance_281/clk_in instance_282/clk_in instance_281/data_in instance_282/data_in
+ instance_281/latch_enable_in instance_282/latch_enable_in instance_281/scan_select_in
+ instance_282/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_292 instance_292/clk_in instance_293/clk_in instance_292/data_in instance_293/data_in
+ instance_292/latch_enable_in instance_293/latch_enable_in instance_292/scan_select_in
+ instance_293/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_260 instance_260/clk_in instance_261/clk_in instance_260/data_in instance_261/data_in
+ instance_260/latch_enable_in instance_261/latch_enable_in instance_260/scan_select_in
+ instance_261/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_271 instance_271/clk_in instance_272/clk_in instance_271/data_in instance_272/data_in
+ instance_271/latch_enable_in instance_272/latch_enable_in instance_271/scan_select_in
+ instance_272/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_282 instance_282/clk_in instance_283/clk_in instance_282/data_in instance_283/data_in
+ instance_282/latch_enable_in instance_283/latch_enable_in instance_282/scan_select_in
+ instance_283/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_293 instance_293/clk_in instance_294/clk_in instance_293/data_in instance_294/data_in
+ instance_293/latch_enable_in instance_294/latch_enable_in instance_293/scan_select_in
+ instance_294/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_250 instance_250/clk_in instance_251/clk_in instance_250/data_in instance_251/data_in
+ instance_250/latch_enable_in instance_251/latch_enable_in instance_250/scan_select_in
+ instance_251/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_261 instance_261/clk_in instance_262/clk_in instance_261/data_in instance_262/data_in
+ instance_261/latch_enable_in instance_262/latch_enable_in instance_261/scan_select_in
+ instance_262/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_272 instance_272/clk_in instance_273/clk_in instance_272/data_in instance_273/data_in
+ instance_272/latch_enable_in instance_273/latch_enable_in instance_272/scan_select_in
+ instance_273/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_283 instance_283/clk_in instance_284/clk_in instance_283/data_in instance_284/data_in
+ instance_283/latch_enable_in instance_284/latch_enable_in instance_283/scan_select_in
+ instance_284/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_294 instance_294/clk_in instance_295/clk_in instance_294/data_in instance_295/data_in
+ instance_294/latch_enable_in instance_295/latch_enable_in instance_294/scan_select_in
+ instance_295/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_90 instance_90/clk_in instance_91/clk_in instance_90/data_in instance_91/data_in
+ instance_90/latch_enable_in instance_91/latch_enable_in instance_90/scan_select_in
+ instance_91/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_240 instance_240/clk_in instance_241/clk_in instance_240/data_in instance_241/data_in
+ instance_240/latch_enable_in instance_241/latch_enable_in instance_240/scan_select_in
+ instance_241/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_251 instance_251/clk_in instance_252/clk_in instance_251/data_in instance_252/data_in
+ instance_251/latch_enable_in instance_252/latch_enable_in instance_251/scan_select_in
+ instance_252/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_262 instance_262/clk_in instance_263/clk_in instance_262/data_in instance_263/data_in
+ instance_262/latch_enable_in instance_263/latch_enable_in instance_262/scan_select_in
+ instance_263/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_273 instance_273/clk_in instance_274/clk_in instance_273/data_in instance_274/data_in
+ instance_273/latch_enable_in instance_274/latch_enable_in instance_273/scan_select_in
+ instance_274/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_284 instance_284/clk_in instance_285/clk_in instance_284/data_in instance_285/data_in
+ instance_284/latch_enable_in instance_285/latch_enable_in instance_284/scan_select_in
+ instance_285/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_295 instance_295/clk_in instance_296/clk_in instance_295/data_in instance_296/data_in
+ instance_295/latch_enable_in instance_296/latch_enable_in instance_295/scan_select_in
+ instance_296/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_91 instance_91/clk_in instance_92/clk_in instance_91/data_in instance_92/data_in
+ instance_91/latch_enable_in instance_92/latch_enable_in instance_91/scan_select_in
+ instance_92/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_80 instance_80/clk_in instance_81/clk_in instance_80/data_in instance_81/data_in
+ instance_80/latch_enable_in instance_81/latch_enable_in instance_80/scan_select_in
+ instance_81/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_230 instance_230/clk_in instance_231/clk_in instance_230/data_in instance_231/data_in
+ instance_230/latch_enable_in instance_231/latch_enable_in instance_230/scan_select_in
+ instance_231/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_241 instance_241/clk_in instance_242/clk_in instance_241/data_in instance_242/data_in
+ instance_241/latch_enable_in instance_242/latch_enable_in instance_241/scan_select_in
+ instance_242/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_252 instance_252/clk_in instance_253/clk_in instance_252/data_in instance_253/data_in
+ instance_252/latch_enable_in instance_253/latch_enable_in instance_252/scan_select_in
+ instance_253/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_263 instance_263/clk_in instance_264/clk_in instance_263/data_in instance_264/data_in
+ instance_263/latch_enable_in instance_264/latch_enable_in instance_263/scan_select_in
+ instance_264/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_274 instance_274/clk_in instance_275/clk_in instance_274/data_in instance_275/data_in
+ instance_274/latch_enable_in instance_275/latch_enable_in instance_274/scan_select_in
+ instance_275/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_285 instance_285/clk_in instance_286/clk_in instance_285/data_in instance_286/data_in
+ instance_285/latch_enable_in instance_286/latch_enable_in instance_285/scan_select_in
+ instance_286/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_296 instance_296/clk_in instance_297/clk_in instance_296/data_in instance_297/data_in
+ instance_296/latch_enable_in instance_297/latch_enable_in instance_296/scan_select_in
+ instance_297/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_92 instance_92/clk_in instance_93/clk_in instance_92/data_in instance_93/data_in
+ instance_92/latch_enable_in instance_93/latch_enable_in instance_92/scan_select_in
+ instance_93/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_81 instance_81/clk_in instance_82/clk_in instance_81/data_in instance_82/data_in
+ instance_81/latch_enable_in instance_82/latch_enable_in instance_81/scan_select_in
+ instance_82/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_70 instance_70/clk_in instance_71/clk_in instance_70/data_in instance_71/data_in
+ instance_70/latch_enable_in instance_71/latch_enable_in instance_70/scan_select_in
+ instance_71/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_220 instance_220/clk_in instance_221/clk_in instance_220/data_in instance_221/data_in
+ instance_220/latch_enable_in instance_221/latch_enable_in instance_220/scan_select_in
+ instance_221/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_231 instance_231/clk_in instance_232/clk_in instance_231/data_in instance_232/data_in
+ instance_231/latch_enable_in instance_232/latch_enable_in instance_231/scan_select_in
+ instance_232/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_242 instance_242/clk_in instance_243/clk_in instance_242/data_in instance_243/data_in
+ instance_242/latch_enable_in instance_243/latch_enable_in instance_242/scan_select_in
+ instance_243/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_253 instance_253/clk_in instance_254/clk_in instance_253/data_in instance_254/data_in
+ instance_253/latch_enable_in instance_254/latch_enable_in instance_253/scan_select_in
+ instance_254/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_264 instance_264/clk_in instance_265/clk_in instance_264/data_in instance_265/data_in
+ instance_264/latch_enable_in instance_265/latch_enable_in instance_264/scan_select_in
+ instance_265/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_275 instance_275/clk_in instance_276/clk_in instance_275/data_in instance_276/data_in
+ instance_275/latch_enable_in instance_276/latch_enable_in instance_275/scan_select_in
+ instance_276/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_286 instance_286/clk_in instance_287/clk_in instance_286/data_in instance_287/data_in
+ instance_286/latch_enable_in instance_287/latch_enable_in instance_286/scan_select_in
+ instance_287/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_297 instance_297/clk_in instance_298/clk_in instance_297/data_in instance_298/data_in
+ instance_297/latch_enable_in instance_298/latch_enable_in instance_297/scan_select_in
+ instance_298/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_0 io_in[8] instance_1/clk_in io_in[9] instance_1/data_in io_in[11] instance_1/latch_enable_in
+ io_in[10] instance_1/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_93 instance_93/clk_in instance_94/clk_in instance_93/data_in instance_94/data_in
+ instance_93/latch_enable_in instance_94/latch_enable_in instance_93/scan_select_in
+ instance_94/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_82 instance_82/clk_in instance_83/clk_in instance_82/data_in instance_83/data_in
+ instance_82/latch_enable_in instance_83/latch_enable_in instance_82/scan_select_in
+ instance_83/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_71 instance_71/clk_in instance_72/clk_in instance_71/data_in instance_72/data_in
+ instance_71/latch_enable_in instance_72/latch_enable_in instance_71/scan_select_in
+ instance_72/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_60 instance_60/clk_in instance_61/clk_in instance_60/data_in instance_61/data_in
+ instance_60/latch_enable_in instance_61/latch_enable_in instance_60/scan_select_in
+ instance_61/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_210 instance_210/clk_in instance_211/clk_in instance_210/data_in instance_211/data_in
+ instance_210/latch_enable_in instance_211/latch_enable_in instance_210/scan_select_in
+ instance_211/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_221 instance_221/clk_in instance_222/clk_in instance_221/data_in instance_222/data_in
+ instance_221/latch_enable_in instance_222/latch_enable_in instance_221/scan_select_in
+ instance_222/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_232 instance_232/clk_in instance_233/clk_in instance_232/data_in instance_233/data_in
+ instance_232/latch_enable_in instance_233/latch_enable_in instance_232/scan_select_in
+ instance_233/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_243 instance_243/clk_in instance_244/clk_in instance_243/data_in instance_244/data_in
+ instance_243/latch_enable_in instance_244/latch_enable_in instance_243/scan_select_in
+ instance_244/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_254 instance_254/clk_in instance_255/clk_in instance_254/data_in instance_255/data_in
+ instance_254/latch_enable_in instance_255/latch_enable_in instance_254/scan_select_in
+ instance_255/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_265 instance_265/clk_in instance_266/clk_in instance_265/data_in instance_266/data_in
+ instance_265/latch_enable_in instance_266/latch_enable_in instance_265/scan_select_in
+ instance_266/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_276 instance_276/clk_in instance_277/clk_in instance_276/data_in instance_277/data_in
+ instance_276/latch_enable_in instance_277/latch_enable_in instance_276/scan_select_in
+ instance_277/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_287 instance_287/clk_in instance_288/clk_in instance_287/data_in instance_288/data_in
+ instance_287/latch_enable_in instance_288/latch_enable_in instance_287/scan_select_in
+ instance_288/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_298 instance_298/clk_in instance_299/clk_in instance_298/data_in instance_299/data_in
+ instance_298/latch_enable_in instance_299/latch_enable_in instance_298/scan_select_in
+ instance_299/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_1 instance_1/clk_in instance_2/clk_in instance_1/data_in instance_2/data_in
+ instance_1/latch_enable_in instance_2/latch_enable_in instance_1/scan_select_in
+ instance_2/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_94 instance_94/clk_in instance_95/clk_in instance_94/data_in instance_95/data_in
+ instance_94/latch_enable_in instance_95/latch_enable_in instance_94/scan_select_in
+ instance_95/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_83 instance_83/clk_in instance_84/clk_in instance_83/data_in instance_84/data_in
+ instance_83/latch_enable_in instance_84/latch_enable_in instance_83/scan_select_in
+ instance_84/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_72 instance_72/clk_in instance_73/clk_in instance_72/data_in instance_73/data_in
+ instance_72/latch_enable_in instance_73/latch_enable_in instance_72/scan_select_in
+ instance_73/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_61 instance_61/clk_in instance_62/clk_in instance_61/data_in instance_62/data_in
+ instance_61/latch_enable_in instance_62/latch_enable_in instance_61/scan_select_in
+ instance_62/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_50 instance_50/clk_in instance_51/clk_in instance_50/data_in instance_51/data_in
+ instance_50/latch_enable_in instance_51/latch_enable_in instance_50/scan_select_in
+ instance_51/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_200 instance_200/clk_in instance_201/clk_in instance_200/data_in instance_201/data_in
+ instance_200/latch_enable_in instance_201/latch_enable_in instance_200/scan_select_in
+ instance_201/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_211 instance_211/clk_in instance_212/clk_in instance_211/data_in instance_212/data_in
+ instance_211/latch_enable_in instance_212/latch_enable_in instance_211/scan_select_in
+ instance_212/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_222 instance_222/clk_in instance_223/clk_in instance_222/data_in instance_223/data_in
+ instance_222/latch_enable_in instance_223/latch_enable_in instance_222/scan_select_in
+ instance_223/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_233 instance_233/clk_in instance_234/clk_in instance_233/data_in instance_234/data_in
+ instance_233/latch_enable_in instance_234/latch_enable_in instance_233/scan_select_in
+ instance_234/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_244 instance_244/clk_in instance_245/clk_in instance_244/data_in instance_245/data_in
+ instance_244/latch_enable_in instance_245/latch_enable_in instance_244/scan_select_in
+ instance_245/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_255 instance_255/clk_in instance_256/clk_in instance_255/data_in instance_256/data_in
+ instance_255/latch_enable_in instance_256/latch_enable_in instance_255/scan_select_in
+ instance_256/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_266 instance_266/clk_in instance_267/clk_in instance_266/data_in instance_267/data_in
+ instance_266/latch_enable_in instance_267/latch_enable_in instance_266/scan_select_in
+ instance_267/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_277 instance_277/clk_in instance_278/clk_in instance_277/data_in instance_278/data_in
+ instance_277/latch_enable_in instance_278/latch_enable_in instance_277/scan_select_in
+ instance_278/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_288 instance_288/clk_in instance_289/clk_in instance_288/data_in instance_289/data_in
+ instance_288/latch_enable_in instance_289/latch_enable_in instance_288/scan_select_in
+ instance_289/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_299 instance_299/clk_in instance_300/clk_in instance_299/data_in instance_300/data_in
+ instance_299/latch_enable_in instance_300/latch_enable_in instance_299/scan_select_in
+ instance_300/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_2 instance_2/clk_in instance_3/clk_in instance_2/data_in instance_3/data_in
+ instance_2/latch_enable_in instance_3/latch_enable_in instance_2/scan_select_in
+ instance_3/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_95 instance_95/clk_in instance_96/clk_in instance_95/data_in instance_96/data_in
+ instance_95/latch_enable_in instance_96/latch_enable_in instance_95/scan_select_in
+ instance_96/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_84 instance_84/clk_in instance_85/clk_in instance_84/data_in instance_85/data_in
+ instance_84/latch_enable_in instance_85/latch_enable_in instance_84/scan_select_in
+ instance_85/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_73 instance_73/clk_in instance_74/clk_in instance_73/data_in instance_74/data_in
+ instance_73/latch_enable_in instance_74/latch_enable_in instance_73/scan_select_in
+ instance_74/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_62 instance_62/clk_in instance_63/clk_in instance_62/data_in instance_63/data_in
+ instance_62/latch_enable_in instance_63/latch_enable_in instance_62/scan_select_in
+ instance_63/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_51 instance_51/clk_in instance_52/clk_in instance_51/data_in instance_52/data_in
+ instance_51/latch_enable_in instance_52/latch_enable_in instance_51/scan_select_in
+ instance_52/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_40 instance_40/clk_in instance_41/clk_in instance_40/data_in instance_41/data_in
+ instance_40/latch_enable_in instance_41/latch_enable_in instance_40/scan_select_in
+ instance_41/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_201 instance_201/clk_in instance_202/clk_in instance_201/data_in instance_202/data_in
+ instance_201/latch_enable_in instance_202/latch_enable_in instance_201/scan_select_in
+ instance_202/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_212 instance_212/clk_in instance_213/clk_in instance_212/data_in instance_213/data_in
+ instance_212/latch_enable_in instance_213/latch_enable_in instance_212/scan_select_in
+ instance_213/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_223 instance_223/clk_in instance_224/clk_in instance_223/data_in instance_224/data_in
+ instance_223/latch_enable_in instance_224/latch_enable_in instance_223/scan_select_in
+ instance_224/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_234 instance_234/clk_in instance_235/clk_in instance_234/data_in instance_235/data_in
+ instance_234/latch_enable_in instance_235/latch_enable_in instance_234/scan_select_in
+ instance_235/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_245 instance_245/clk_in instance_246/clk_in instance_245/data_in instance_246/data_in
+ instance_245/latch_enable_in instance_246/latch_enable_in instance_245/scan_select_in
+ instance_246/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_256 instance_256/clk_in instance_257/clk_in instance_256/data_in instance_257/data_in
+ instance_256/latch_enable_in instance_257/latch_enable_in instance_256/scan_select_in
+ instance_257/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_267 instance_267/clk_in instance_268/clk_in instance_267/data_in instance_268/data_in
+ instance_267/latch_enable_in instance_268/latch_enable_in instance_267/scan_select_in
+ instance_268/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_278 instance_278/clk_in instance_279/clk_in instance_278/data_in instance_279/data_in
+ instance_278/latch_enable_in instance_279/latch_enable_in instance_278/scan_select_in
+ instance_279/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_289 instance_289/clk_in instance_290/clk_in instance_289/data_in instance_290/data_in
+ instance_289/latch_enable_in instance_290/latch_enable_in instance_289/scan_select_in
+ instance_290/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_3 instance_3/clk_in instance_4/clk_in instance_3/data_in instance_4/data_in
+ instance_3/latch_enable_in instance_4/latch_enable_in instance_3/scan_select_in
+ instance_4/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_85 instance_85/clk_in instance_86/clk_in instance_85/data_in instance_86/data_in
+ instance_85/latch_enable_in instance_86/latch_enable_in instance_85/scan_select_in
+ instance_86/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_74 instance_74/clk_in instance_75/clk_in instance_74/data_in instance_75/data_in
+ instance_74/latch_enable_in instance_75/latch_enable_in instance_74/scan_select_in
+ instance_75/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_63 instance_63/clk_in instance_64/clk_in instance_63/data_in instance_64/data_in
+ instance_63/latch_enable_in instance_64/latch_enable_in instance_63/scan_select_in
+ instance_64/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_52 instance_52/clk_in instance_53/clk_in instance_52/data_in instance_53/data_in
+ instance_52/latch_enable_in instance_53/latch_enable_in instance_52/scan_select_in
+ instance_53/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_41 instance_41/clk_in instance_42/clk_in instance_41/data_in instance_42/data_in
+ instance_41/latch_enable_in instance_42/latch_enable_in instance_41/scan_select_in
+ instance_42/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_30 instance_30/clk_in instance_31/clk_in instance_30/data_in instance_31/data_in
+ instance_30/latch_enable_in instance_31/latch_enable_in instance_30/scan_select_in
+ instance_31/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_96 instance_96/clk_in instance_97/clk_in instance_96/data_in instance_97/data_in
+ instance_96/latch_enable_in instance_97/latch_enable_in instance_96/scan_select_in
+ instance_97/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_202 instance_202/clk_in instance_203/clk_in instance_202/data_in instance_203/data_in
+ instance_202/latch_enable_in instance_203/latch_enable_in instance_202/scan_select_in
+ instance_203/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_213 instance_213/clk_in instance_214/clk_in instance_213/data_in instance_214/data_in
+ instance_213/latch_enable_in instance_214/latch_enable_in instance_213/scan_select_in
+ instance_214/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_224 instance_224/clk_in instance_225/clk_in instance_224/data_in instance_225/data_in
+ instance_224/latch_enable_in instance_225/latch_enable_in instance_224/scan_select_in
+ instance_225/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_235 instance_235/clk_in instance_236/clk_in instance_235/data_in instance_236/data_in
+ instance_235/latch_enable_in instance_236/latch_enable_in instance_235/scan_select_in
+ instance_236/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_246 instance_246/clk_in instance_247/clk_in instance_246/data_in instance_247/data_in
+ instance_246/latch_enable_in instance_247/latch_enable_in instance_246/scan_select_in
+ instance_247/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_257 instance_257/clk_in instance_258/clk_in instance_257/data_in instance_258/data_in
+ instance_257/latch_enable_in instance_258/latch_enable_in instance_257/scan_select_in
+ instance_258/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_268 instance_268/clk_in instance_269/clk_in instance_268/data_in instance_269/data_in
+ instance_268/latch_enable_in instance_269/latch_enable_in instance_268/scan_select_in
+ instance_269/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_279 instance_279/clk_in instance_280/clk_in instance_279/data_in instance_280/data_in
+ instance_279/latch_enable_in instance_280/latch_enable_in instance_279/scan_select_in
+ instance_280/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_4 instance_4/clk_in instance_5/clk_in instance_4/data_in instance_5/data_in
+ instance_4/latch_enable_in instance_5/latch_enable_in instance_4/scan_select_in
+ instance_5/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_86 instance_86/clk_in instance_87/clk_in instance_86/data_in instance_87/data_in
+ instance_86/latch_enable_in instance_87/latch_enable_in instance_86/scan_select_in
+ instance_87/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_75 instance_75/clk_in instance_76/clk_in instance_75/data_in instance_76/data_in
+ instance_75/latch_enable_in instance_76/latch_enable_in instance_75/scan_select_in
+ instance_76/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_64 instance_64/clk_in instance_65/clk_in instance_64/data_in instance_65/data_in
+ instance_64/latch_enable_in instance_65/latch_enable_in instance_64/scan_select_in
+ instance_65/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_53 instance_53/clk_in instance_54/clk_in instance_53/data_in instance_54/data_in
+ instance_53/latch_enable_in instance_54/latch_enable_in instance_53/scan_select_in
+ instance_54/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_42 instance_42/clk_in instance_43/clk_in instance_42/data_in instance_43/data_in
+ instance_42/latch_enable_in instance_43/latch_enable_in instance_42/scan_select_in
+ instance_43/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_31 instance_31/clk_in instance_32/clk_in instance_31/data_in instance_32/data_in
+ instance_31/latch_enable_in instance_32/latch_enable_in instance_31/scan_select_in
+ instance_32/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_20 instance_20/clk_in instance_21/clk_in instance_20/data_in instance_21/data_in
+ instance_20/latch_enable_in instance_21/latch_enable_in instance_20/scan_select_in
+ instance_21/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_97 instance_97/clk_in instance_98/clk_in instance_97/data_in instance_98/data_in
+ instance_97/latch_enable_in instance_98/latch_enable_in instance_97/scan_select_in
+ instance_98/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_203 instance_203/clk_in instance_204/clk_in instance_203/data_in instance_204/data_in
+ instance_203/latch_enable_in instance_204/latch_enable_in instance_203/scan_select_in
+ instance_204/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_214 instance_214/clk_in instance_215/clk_in instance_214/data_in instance_215/data_in
+ instance_214/latch_enable_in instance_215/latch_enable_in instance_214/scan_select_in
+ instance_215/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_225 instance_225/clk_in instance_226/clk_in instance_225/data_in instance_226/data_in
+ instance_225/latch_enable_in instance_226/latch_enable_in instance_225/scan_select_in
+ instance_226/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_236 instance_236/clk_in instance_237/clk_in instance_236/data_in instance_237/data_in
+ instance_236/latch_enable_in instance_237/latch_enable_in instance_236/scan_select_in
+ instance_237/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_247 instance_247/clk_in instance_248/clk_in instance_247/data_in instance_248/data_in
+ instance_247/latch_enable_in instance_248/latch_enable_in instance_247/scan_select_in
+ instance_248/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_258 instance_258/clk_in instance_259/clk_in instance_258/data_in instance_259/data_in
+ instance_258/latch_enable_in instance_259/latch_enable_in instance_258/scan_select_in
+ instance_259/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_269 instance_269/clk_in instance_270/clk_in instance_269/data_in instance_270/data_in
+ instance_269/latch_enable_in instance_270/latch_enable_in instance_269/scan_select_in
+ instance_270/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_5 instance_5/clk_in instance_6/clk_in instance_5/data_in instance_6/data_in
+ instance_5/latch_enable_in instance_6/latch_enable_in instance_5/scan_select_in
+ instance_6/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_87 instance_87/clk_in instance_88/clk_in instance_87/data_in instance_88/data_in
+ instance_87/latch_enable_in instance_88/latch_enable_in instance_87/scan_select_in
+ instance_88/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_76 instance_76/clk_in instance_77/clk_in instance_76/data_in instance_77/data_in
+ instance_76/latch_enable_in instance_77/latch_enable_in instance_76/scan_select_in
+ instance_77/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_65 instance_65/clk_in instance_66/clk_in instance_65/data_in instance_66/data_in
+ instance_65/latch_enable_in instance_66/latch_enable_in instance_65/scan_select_in
+ instance_66/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_54 instance_54/clk_in instance_55/clk_in instance_54/data_in instance_55/data_in
+ instance_54/latch_enable_in instance_55/latch_enable_in instance_54/scan_select_in
+ instance_55/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_43 instance_43/clk_in instance_44/clk_in instance_43/data_in instance_44/data_in
+ instance_43/latch_enable_in instance_44/latch_enable_in instance_43/scan_select_in
+ instance_44/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_32 instance_32/clk_in instance_33/clk_in instance_32/data_in instance_33/data_in
+ instance_32/latch_enable_in instance_33/latch_enable_in instance_32/scan_select_in
+ instance_33/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_21 instance_21/clk_in instance_22/clk_in instance_21/data_in instance_22/data_in
+ instance_21/latch_enable_in instance_22/latch_enable_in instance_21/scan_select_in
+ instance_22/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_10 instance_9/clk_out instance_11/clk_in instance_9/data_out instance_11/data_in
+ instance_9/latch_enable_out instance_11/latch_enable_in instance_9/scan_select_out
+ instance_11/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_98 instance_98/clk_in instance_99/clk_in instance_98/data_in instance_99/data_in
+ instance_98/latch_enable_in instance_99/latch_enable_in instance_98/scan_select_in
+ instance_99/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_204 instance_204/clk_in instance_205/clk_in instance_204/data_in instance_205/data_in
+ instance_204/latch_enable_in instance_205/latch_enable_in instance_204/scan_select_in
+ instance_205/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_215 instance_215/clk_in instance_216/clk_in instance_215/data_in instance_216/data_in
+ instance_215/latch_enable_in instance_216/latch_enable_in instance_215/scan_select_in
+ instance_216/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_226 instance_226/clk_in instance_227/clk_in instance_226/data_in instance_227/data_in
+ instance_226/latch_enable_in instance_227/latch_enable_in instance_226/scan_select_in
+ instance_227/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_237 instance_237/clk_in instance_238/clk_in instance_237/data_in instance_238/data_in
+ instance_237/latch_enable_in instance_238/latch_enable_in instance_237/scan_select_in
+ instance_238/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_248 instance_248/clk_in instance_249/clk_in instance_248/data_in instance_249/data_in
+ instance_248/latch_enable_in instance_249/latch_enable_in instance_248/scan_select_in
+ instance_249/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_259 instance_259/clk_in instance_260/clk_in instance_259/data_in instance_260/data_in
+ instance_259/latch_enable_in instance_260/latch_enable_in instance_259/scan_select_in
+ instance_260/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_6 instance_6/clk_in instance_7/clk_in instance_6/data_in instance_7/data_in
+ instance_6/latch_enable_in instance_7/latch_enable_in instance_6/scan_select_in
+ instance_7/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_88 instance_88/clk_in instance_89/clk_in instance_88/data_in instance_89/data_in
+ instance_88/latch_enable_in instance_89/latch_enable_in instance_88/scan_select_in
+ instance_89/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_77 instance_77/clk_in instance_78/clk_in instance_77/data_in instance_78/data_in
+ instance_77/latch_enable_in instance_78/latch_enable_in instance_77/scan_select_in
+ instance_78/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_66 instance_66/clk_in instance_67/clk_in instance_66/data_in instance_67/data_in
+ instance_66/latch_enable_in instance_67/latch_enable_in instance_66/scan_select_in
+ instance_67/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_55 instance_55/clk_in instance_56/clk_in instance_55/data_in instance_56/data_in
+ instance_55/latch_enable_in instance_56/latch_enable_in instance_55/scan_select_in
+ instance_56/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_44 instance_44/clk_in instance_45/clk_in instance_44/data_in instance_45/data_in
+ instance_44/latch_enable_in instance_45/latch_enable_in instance_44/scan_select_in
+ instance_45/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_33 instance_33/clk_in instance_34/clk_in instance_33/data_in instance_34/data_in
+ instance_33/latch_enable_in instance_34/latch_enable_in instance_33/scan_select_in
+ instance_34/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_22 instance_22/clk_in instance_23/clk_in instance_22/data_in instance_23/data_in
+ instance_22/latch_enable_in instance_23/latch_enable_in instance_22/scan_select_in
+ instance_23/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_11 instance_11/clk_in instance_12/clk_in instance_11/data_in instance_12/data_in
+ instance_11/latch_enable_in instance_12/latch_enable_in instance_11/scan_select_in
+ instance_12/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_99 instance_99/clk_in instance_99/clk_out instance_99/data_in instance_99/data_out
+ instance_99/latch_enable_in instance_99/latch_enable_out instance_99/scan_select_in
+ instance_99/scan_select_out vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_205 instance_205/clk_in instance_206/clk_in instance_205/data_in instance_206/data_in
+ instance_205/latch_enable_in instance_206/latch_enable_in instance_205/scan_select_in
+ instance_206/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_216 instance_216/clk_in instance_217/clk_in instance_216/data_in instance_217/data_in
+ instance_216/latch_enable_in instance_217/latch_enable_in instance_216/scan_select_in
+ instance_217/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_227 instance_227/clk_in instance_228/clk_in instance_227/data_in instance_228/data_in
+ instance_227/latch_enable_in instance_228/latch_enable_in instance_227/scan_select_in
+ instance_228/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_238 instance_238/clk_in instance_239/clk_in instance_238/data_in instance_239/data_in
+ instance_238/latch_enable_in instance_239/latch_enable_in instance_238/scan_select_in
+ instance_239/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_249 instance_249/clk_in instance_250/clk_in instance_249/data_in instance_250/data_in
+ instance_249/latch_enable_in instance_250/latch_enable_in instance_249/scan_select_in
+ instance_250/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_7 instance_7/clk_in instance_8/clk_in instance_7/data_in instance_8/data_in
+ instance_7/latch_enable_in instance_8/latch_enable_in instance_7/scan_select_in
+ instance_8/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_89 instance_89/clk_in instance_90/clk_in instance_89/data_in instance_90/data_in
+ instance_89/latch_enable_in instance_90/latch_enable_in instance_89/scan_select_in
+ instance_90/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_78 instance_78/clk_in instance_79/clk_in instance_78/data_in instance_79/data_in
+ instance_78/latch_enable_in instance_79/latch_enable_in instance_78/scan_select_in
+ instance_79/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_67 instance_67/clk_in instance_68/clk_in instance_67/data_in instance_68/data_in
+ instance_67/latch_enable_in instance_68/latch_enable_in instance_67/scan_select_in
+ instance_68/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_56 instance_56/clk_in instance_57/clk_in instance_56/data_in instance_57/data_in
+ instance_56/latch_enable_in instance_57/latch_enable_in instance_56/scan_select_in
+ instance_57/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_45 instance_45/clk_in instance_46/clk_in instance_45/data_in instance_46/data_in
+ instance_45/latch_enable_in instance_46/latch_enable_in instance_45/scan_select_in
+ instance_46/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_34 instance_34/clk_in instance_35/clk_in instance_34/data_in instance_35/data_in
+ instance_34/latch_enable_in instance_35/latch_enable_in instance_34/scan_select_in
+ instance_35/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_23 instance_23/clk_in instance_24/clk_in instance_23/data_in instance_24/data_in
+ instance_23/latch_enable_in instance_24/latch_enable_in instance_23/scan_select_in
+ instance_24/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_12 instance_12/clk_in instance_13/clk_in instance_12/data_in instance_13/data_in
+ instance_12/latch_enable_in instance_13/latch_enable_in instance_12/scan_select_in
+ instance_13/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_206 instance_206/clk_in instance_207/clk_in instance_206/data_in instance_207/data_in
+ instance_206/latch_enable_in instance_207/latch_enable_in instance_206/scan_select_in
+ instance_207/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_217 instance_217/clk_in instance_218/clk_in instance_217/data_in instance_218/data_in
+ instance_217/latch_enable_in instance_218/latch_enable_in instance_217/scan_select_in
+ instance_218/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_228 instance_228/clk_in instance_229/clk_in instance_228/data_in instance_229/data_in
+ instance_228/latch_enable_in instance_229/latch_enable_in instance_228/scan_select_in
+ instance_229/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_239 instance_239/clk_in instance_240/clk_in instance_239/data_in instance_240/data_in
+ instance_239/latch_enable_in instance_240/latch_enable_in instance_239/scan_select_in
+ instance_240/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_8 instance_8/clk_in instance_9/clk_in instance_8/data_in instance_9/data_in
+ instance_8/latch_enable_in instance_9/latch_enable_in instance_8/scan_select_in
+ instance_9/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_79 instance_79/clk_in instance_80/clk_in instance_79/data_in instance_80/data_in
+ instance_79/latch_enable_in instance_80/latch_enable_in instance_79/scan_select_in
+ instance_80/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_68 instance_68/clk_in instance_69/clk_in instance_68/data_in instance_69/data_in
+ instance_68/latch_enable_in instance_69/latch_enable_in instance_68/scan_select_in
+ instance_69/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_57 instance_57/clk_in instance_58/clk_in instance_57/data_in instance_58/data_in
+ instance_57/latch_enable_in instance_58/latch_enable_in instance_57/scan_select_in
+ instance_58/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_46 instance_46/clk_in instance_47/clk_in instance_46/data_in instance_47/data_in
+ instance_46/latch_enable_in instance_47/latch_enable_in instance_46/scan_select_in
+ instance_47/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_35 instance_35/clk_in instance_36/clk_in instance_35/data_in instance_36/data_in
+ instance_35/latch_enable_in instance_36/latch_enable_in instance_35/scan_select_in
+ instance_36/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_24 instance_24/clk_in instance_25/clk_in instance_24/data_in instance_25/data_in
+ instance_24/latch_enable_in instance_25/latch_enable_in instance_24/scan_select_in
+ instance_25/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_13 instance_13/clk_in instance_14/clk_in instance_13/data_in instance_14/data_in
+ instance_13/latch_enable_in instance_14/latch_enable_in instance_13/scan_select_in
+ instance_14/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_207 instance_207/clk_in instance_208/clk_in instance_207/data_in instance_208/data_in
+ instance_207/latch_enable_in instance_208/latch_enable_in instance_207/scan_select_in
+ instance_208/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_218 instance_218/clk_in instance_219/clk_in instance_218/data_in instance_219/data_in
+ instance_218/latch_enable_in instance_219/latch_enable_in instance_218/scan_select_in
+ instance_219/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_229 instance_229/clk_in instance_230/clk_in instance_229/data_in instance_230/data_in
+ instance_229/latch_enable_in instance_230/latch_enable_in instance_229/scan_select_in
+ instance_230/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_390 instance_390/clk_in instance_390/clk_out instance_390/data_in io_out[11]
+ instance_390/latch_enable_in instance_390/latch_enable_out instance_390/scan_select_in
+ instance_390/scan_select_out vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_9 instance_9/clk_in instance_9/clk_out instance_9/data_in instance_9/data_out
+ instance_9/latch_enable_in instance_9/latch_enable_out instance_9/scan_select_in
+ instance_9/scan_select_out vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_69 instance_69/clk_in instance_70/clk_in instance_69/data_in instance_70/data_in
+ instance_69/latch_enable_in instance_70/latch_enable_in instance_69/scan_select_in
+ instance_70/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_58 instance_58/clk_in instance_59/clk_in instance_58/data_in instance_59/data_in
+ instance_58/latch_enable_in instance_59/latch_enable_in instance_58/scan_select_in
+ instance_59/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_47 instance_47/clk_in instance_48/clk_in instance_47/data_in instance_48/data_in
+ instance_47/latch_enable_in instance_48/latch_enable_in instance_47/scan_select_in
+ instance_48/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_36 instance_36/clk_in instance_37/clk_in instance_36/data_in instance_37/data_in
+ instance_36/latch_enable_in instance_37/latch_enable_in instance_36/scan_select_in
+ instance_37/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_25 instance_25/clk_in instance_26/clk_in instance_25/data_in instance_26/data_in
+ instance_25/latch_enable_in instance_26/latch_enable_in instance_25/scan_select_in
+ instance_26/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_14 instance_14/clk_in instance_15/clk_in instance_14/data_in instance_15/data_in
+ instance_14/latch_enable_in instance_15/latch_enable_in instance_14/scan_select_in
+ instance_15/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_208 instance_208/clk_in instance_209/clk_in instance_208/data_in instance_209/data_in
+ instance_208/latch_enable_in instance_209/latch_enable_in instance_208/scan_select_in
+ instance_209/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_219 instance_219/clk_in instance_220/clk_in instance_219/data_in instance_220/data_in
+ instance_219/latch_enable_in instance_220/latch_enable_in instance_219/scan_select_in
+ instance_220/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_380 instance_380/clk_in instance_381/clk_in instance_380/data_in instance_381/data_in
+ instance_380/latch_enable_in instance_381/latch_enable_in instance_380/scan_select_in
+ instance_381/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_59 instance_59/clk_in instance_60/clk_in instance_59/data_in instance_60/data_in
+ instance_59/latch_enable_in instance_60/latch_enable_in instance_59/scan_select_in
+ instance_60/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_48 instance_48/clk_in instance_49/clk_in instance_48/data_in instance_49/data_in
+ instance_48/latch_enable_in instance_49/latch_enable_in instance_48/scan_select_in
+ instance_49/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_37 instance_37/clk_in instance_38/clk_in instance_37/data_in instance_38/data_in
+ instance_37/latch_enable_in instance_38/latch_enable_in instance_37/scan_select_in
+ instance_38/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_26 instance_26/clk_in instance_27/clk_in instance_26/data_in instance_27/data_in
+ instance_26/latch_enable_in instance_27/latch_enable_in instance_26/scan_select_in
+ instance_27/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_15 instance_15/clk_in instance_16/clk_in instance_15/data_in instance_16/data_in
+ instance_15/latch_enable_in instance_16/latch_enable_in instance_15/scan_select_in
+ instance_16/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_209 instance_209/clk_in instance_210/clk_in instance_209/data_in instance_210/data_in
+ instance_209/latch_enable_in instance_210/latch_enable_in instance_209/scan_select_in
+ instance_210/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_370 instance_370/clk_in instance_371/clk_in instance_370/data_in instance_371/data_in
+ instance_370/latch_enable_in instance_371/latch_enable_in instance_370/scan_select_in
+ instance_371/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_381 instance_381/clk_in instance_382/clk_in instance_381/data_in instance_382/data_in
+ instance_381/latch_enable_in instance_382/latch_enable_in instance_381/scan_select_in
+ instance_382/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_16 instance_16/clk_in instance_17/clk_in instance_16/data_in instance_17/data_in
+ instance_16/latch_enable_in instance_17/latch_enable_in instance_16/scan_select_in
+ instance_17/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_49 instance_49/clk_in instance_50/clk_in instance_49/data_in instance_50/data_in
+ instance_49/latch_enable_in instance_50/latch_enable_in instance_49/scan_select_in
+ instance_50/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_38 instance_38/clk_in instance_39/clk_in instance_38/data_in instance_39/data_in
+ instance_38/latch_enable_in instance_39/latch_enable_in instance_38/scan_select_in
+ instance_39/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_27 instance_27/clk_in instance_28/clk_in instance_27/data_in instance_28/data_in
+ instance_27/latch_enable_in instance_28/latch_enable_in instance_27/scan_select_in
+ instance_28/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_360 instance_360/clk_in instance_361/clk_in instance_360/data_in instance_361/data_in
+ instance_360/latch_enable_in instance_361/latch_enable_in instance_360/scan_select_in
+ instance_361/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_371 instance_371/clk_in instance_372/clk_in instance_371/data_in instance_372/data_in
+ instance_371/latch_enable_in instance_372/latch_enable_in instance_371/scan_select_in
+ instance_372/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_382 instance_382/clk_in instance_383/clk_in instance_382/data_in instance_383/data_in
+ instance_382/latch_enable_in instance_383/latch_enable_in instance_382/scan_select_in
+ instance_383/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_190 instance_190/clk_in instance_191/clk_in instance_190/data_in instance_191/data_in
+ instance_190/latch_enable_in instance_191/latch_enable_in instance_190/scan_select_in
+ instance_191/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_39 instance_39/clk_in instance_40/clk_in instance_39/data_in instance_40/data_in
+ instance_39/latch_enable_in instance_40/latch_enable_in instance_39/scan_select_in
+ instance_40/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_28 instance_28/clk_in instance_29/clk_in instance_28/data_in instance_29/data_in
+ instance_28/latch_enable_in instance_29/latch_enable_in instance_28/scan_select_in
+ instance_29/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_17 instance_17/clk_in instance_18/clk_in instance_17/data_in instance_18/data_in
+ instance_17/latch_enable_in instance_18/latch_enable_in instance_17/scan_select_in
+ instance_18/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_350 instance_350/clk_in instance_351/clk_in instance_350/data_in instance_351/data_in
+ instance_350/latch_enable_in instance_351/latch_enable_in instance_350/scan_select_in
+ instance_351/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_361 instance_361/clk_in instance_362/clk_in instance_361/data_in instance_362/data_in
+ instance_361/latch_enable_in instance_362/latch_enable_in instance_361/scan_select_in
+ instance_362/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_372 instance_372/clk_in instance_373/clk_in instance_372/data_in instance_373/data_in
+ instance_372/latch_enable_in instance_373/latch_enable_in instance_372/scan_select_in
+ instance_373/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_383 instance_383/clk_in instance_384/clk_in instance_383/data_in instance_384/data_in
+ instance_383/latch_enable_in instance_384/latch_enable_in instance_383/scan_select_in
+ instance_384/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_180 instance_180/clk_in instance_181/clk_in instance_180/data_in instance_181/data_in
+ instance_180/latch_enable_in instance_181/latch_enable_in instance_180/scan_select_in
+ instance_181/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_191 instance_191/clk_in instance_192/clk_in instance_191/data_in instance_192/data_in
+ instance_191/latch_enable_in instance_192/latch_enable_in instance_191/scan_select_in
+ instance_192/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_29 instance_29/clk_in instance_30/clk_in instance_29/data_in instance_30/data_in
+ instance_29/latch_enable_in instance_30/latch_enable_in instance_29/scan_select_in
+ instance_30/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_18 instance_18/clk_in instance_19/clk_in instance_18/data_in instance_19/data_in
+ instance_18/latch_enable_in instance_19/latch_enable_in instance_18/scan_select_in
+ instance_19/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_340 instance_340/clk_in instance_341/clk_in instance_340/data_in instance_341/data_in
+ instance_340/latch_enable_in instance_341/latch_enable_in instance_340/scan_select_in
+ instance_341/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_351 instance_351/clk_in instance_352/clk_in instance_351/data_in instance_352/data_in
+ instance_351/latch_enable_in instance_352/latch_enable_in instance_351/scan_select_in
+ instance_352/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_362 instance_362/clk_in instance_363/clk_in instance_362/data_in instance_363/data_in
+ instance_362/latch_enable_in instance_363/latch_enable_in instance_362/scan_select_in
+ instance_363/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_373 instance_373/clk_in instance_374/clk_in instance_373/data_in instance_374/data_in
+ instance_373/latch_enable_in instance_374/latch_enable_in instance_373/scan_select_in
+ instance_374/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_384 instance_384/clk_in instance_385/clk_in instance_384/data_in instance_385/data_in
+ instance_384/latch_enable_in instance_385/latch_enable_in instance_384/scan_select_in
+ instance_385/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_170 instance_170/clk_in instance_171/clk_in instance_170/data_in instance_171/data_in
+ instance_170/latch_enable_in instance_171/latch_enable_in instance_170/scan_select_in
+ instance_171/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_181 instance_181/clk_in instance_182/clk_in instance_181/data_in instance_182/data_in
+ instance_181/latch_enable_in instance_182/latch_enable_in instance_181/scan_select_in
+ instance_182/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_192 instance_192/clk_in instance_193/clk_in instance_192/data_in instance_193/data_in
+ instance_192/latch_enable_in instance_193/latch_enable_in instance_192/scan_select_in
+ instance_193/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_19 instance_19/clk_in instance_20/clk_in instance_19/data_in instance_20/data_in
+ instance_19/latch_enable_in instance_20/latch_enable_in instance_19/scan_select_in
+ instance_20/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_385 instance_385/clk_in instance_386/clk_in instance_385/data_in instance_386/data_in
+ instance_385/latch_enable_in instance_386/latch_enable_in instance_385/scan_select_in
+ instance_386/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_330 instance_330/clk_in instance_331/clk_in instance_330/data_in instance_331/data_in
+ instance_330/latch_enable_in instance_331/latch_enable_in instance_330/scan_select_in
+ instance_331/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_341 instance_341/clk_in instance_342/clk_in instance_341/data_in instance_342/data_in
+ instance_341/latch_enable_in instance_342/latch_enable_in instance_341/scan_select_in
+ instance_342/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_352 instance_352/clk_in instance_353/clk_in instance_352/data_in instance_353/data_in
+ instance_352/latch_enable_in instance_353/latch_enable_in instance_352/scan_select_in
+ instance_353/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_363 instance_363/clk_in instance_364/clk_in instance_363/data_in instance_364/data_in
+ instance_363/latch_enable_in instance_364/latch_enable_in instance_363/scan_select_in
+ instance_364/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_374 instance_374/clk_in instance_375/clk_in instance_374/data_in instance_375/data_in
+ instance_374/latch_enable_in instance_375/latch_enable_in instance_374/scan_select_in
+ instance_375/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_160 instance_160/clk_in instance_161/clk_in instance_160/data_in instance_161/data_in
+ instance_160/latch_enable_in instance_161/latch_enable_in instance_160/scan_select_in
+ instance_161/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_171 instance_171/clk_in instance_172/clk_in instance_171/data_in instance_172/data_in
+ instance_171/latch_enable_in instance_172/latch_enable_in instance_171/scan_select_in
+ instance_172/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_182 instance_182/clk_in instance_183/clk_in instance_182/data_in instance_183/data_in
+ instance_182/latch_enable_in instance_183/latch_enable_in instance_182/scan_select_in
+ instance_183/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_193 instance_193/clk_in instance_194/clk_in instance_193/data_in instance_194/data_in
+ instance_193/latch_enable_in instance_194/latch_enable_in instance_193/scan_select_in
+ instance_194/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_386 instance_386/clk_in instance_387/clk_in instance_386/data_in instance_387/data_in
+ instance_386/latch_enable_in instance_387/latch_enable_in instance_386/scan_select_in
+ instance_387/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_320 instance_320/clk_in instance_321/clk_in instance_320/data_in instance_321/data_in
+ instance_320/latch_enable_in instance_321/latch_enable_in instance_320/scan_select_in
+ instance_321/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_331 instance_331/clk_in instance_332/clk_in instance_331/data_in instance_332/data_in
+ instance_331/latch_enable_in instance_332/latch_enable_in instance_331/scan_select_in
+ instance_332/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_342 instance_342/clk_in instance_343/clk_in instance_342/data_in instance_343/data_in
+ instance_342/latch_enable_in instance_343/latch_enable_in instance_342/scan_select_in
+ instance_343/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_353 instance_353/clk_in instance_354/clk_in instance_353/data_in instance_354/data_in
+ instance_353/latch_enable_in instance_354/latch_enable_in instance_353/scan_select_in
+ instance_354/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_364 instance_364/clk_in instance_365/clk_in instance_364/data_in instance_365/data_in
+ instance_364/latch_enable_in instance_365/latch_enable_in instance_364/scan_select_in
+ instance_365/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_375 instance_375/clk_in instance_376/clk_in instance_375/data_in instance_376/data_in
+ instance_375/latch_enable_in instance_376/latch_enable_in instance_375/scan_select_in
+ instance_376/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_150 instance_150/clk_in instance_151/clk_in instance_150/data_in instance_151/data_in
+ instance_150/latch_enable_in instance_151/latch_enable_in instance_150/scan_select_in
+ instance_151/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_161 instance_161/clk_in instance_162/clk_in instance_161/data_in instance_162/data_in
+ instance_161/latch_enable_in instance_162/latch_enable_in instance_161/scan_select_in
+ instance_162/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_172 instance_172/clk_in instance_173/clk_in instance_172/data_in instance_173/data_in
+ instance_172/latch_enable_in instance_173/latch_enable_in instance_172/scan_select_in
+ instance_173/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_183 instance_183/clk_in instance_184/clk_in instance_183/data_in instance_184/data_in
+ instance_183/latch_enable_in instance_184/latch_enable_in instance_183/scan_select_in
+ instance_184/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_194 instance_194/clk_in instance_195/clk_in instance_194/data_in instance_195/data_in
+ instance_194/latch_enable_in instance_195/latch_enable_in instance_194/scan_select_in
+ instance_195/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_387 instance_387/clk_in instance_388/clk_in instance_387/data_in instance_388/data_in
+ instance_387/latch_enable_in instance_388/latch_enable_in instance_387/scan_select_in
+ instance_388/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_310 instance_310/clk_in instance_311/clk_in instance_310/data_in instance_311/data_in
+ instance_310/latch_enable_in instance_311/latch_enable_in instance_310/scan_select_in
+ instance_311/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_321 instance_321/clk_in instance_322/clk_in instance_321/data_in instance_322/data_in
+ instance_321/latch_enable_in instance_322/latch_enable_in instance_321/scan_select_in
+ instance_322/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_332 instance_332/clk_in instance_333/clk_in instance_332/data_in instance_333/data_in
+ instance_332/latch_enable_in instance_333/latch_enable_in instance_332/scan_select_in
+ instance_333/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_343 instance_343/clk_in instance_344/clk_in instance_343/data_in instance_344/data_in
+ instance_343/latch_enable_in instance_344/latch_enable_in instance_343/scan_select_in
+ instance_344/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_354 instance_354/clk_in instance_355/clk_in instance_354/data_in instance_355/data_in
+ instance_354/latch_enable_in instance_355/latch_enable_in instance_354/scan_select_in
+ instance_355/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_365 instance_365/clk_in instance_366/clk_in instance_365/data_in instance_366/data_in
+ instance_365/latch_enable_in instance_366/latch_enable_in instance_365/scan_select_in
+ instance_366/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_376 instance_376/clk_in instance_377/clk_in instance_376/data_in instance_377/data_in
+ instance_376/latch_enable_in instance_377/latch_enable_in instance_376/scan_select_in
+ instance_377/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_140 instance_140/clk_in instance_141/clk_in instance_140/data_in instance_141/data_in
+ instance_140/latch_enable_in instance_141/latch_enable_in instance_140/scan_select_in
+ instance_141/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_151 instance_151/clk_in instance_152/clk_in instance_151/data_in instance_152/data_in
+ instance_151/latch_enable_in instance_152/latch_enable_in instance_151/scan_select_in
+ instance_152/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_162 instance_162/clk_in instance_163/clk_in instance_162/data_in instance_163/data_in
+ instance_162/latch_enable_in instance_163/latch_enable_in instance_162/scan_select_in
+ instance_163/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_173 instance_173/clk_in instance_174/clk_in instance_173/data_in instance_174/data_in
+ instance_173/latch_enable_in instance_174/latch_enable_in instance_173/scan_select_in
+ instance_174/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_184 instance_184/clk_in instance_185/clk_in instance_184/data_in instance_185/data_in
+ instance_184/latch_enable_in instance_185/latch_enable_in instance_184/scan_select_in
+ instance_185/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_195 instance_195/clk_in instance_196/clk_in instance_195/data_in instance_196/data_in
+ instance_195/latch_enable_in instance_196/latch_enable_in instance_195/scan_select_in
+ instance_196/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_388 instance_388/clk_in instance_389/clk_in instance_388/data_in instance_389/data_in
+ instance_388/latch_enable_in instance_389/latch_enable_in instance_388/scan_select_in
+ instance_389/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_300 instance_300/clk_in instance_301/clk_in instance_300/data_in instance_301/data_in
+ instance_300/latch_enable_in instance_301/latch_enable_in instance_300/scan_select_in
+ instance_301/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_311 instance_311/clk_in instance_312/clk_in instance_311/data_in instance_312/data_in
+ instance_311/latch_enable_in instance_312/latch_enable_in instance_311/scan_select_in
+ instance_312/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_322 instance_322/clk_in instance_323/clk_in instance_322/data_in instance_323/data_in
+ instance_322/latch_enable_in instance_323/latch_enable_in instance_322/scan_select_in
+ instance_323/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_333 instance_333/clk_in instance_334/clk_in instance_333/data_in instance_334/data_in
+ instance_333/latch_enable_in instance_334/latch_enable_in instance_333/scan_select_in
+ instance_334/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_344 instance_344/clk_in instance_345/clk_in instance_344/data_in instance_345/data_in
+ instance_344/latch_enable_in instance_345/latch_enable_in instance_344/scan_select_in
+ instance_345/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_355 instance_355/clk_in instance_356/clk_in instance_355/data_in instance_356/data_in
+ instance_355/latch_enable_in instance_356/latch_enable_in instance_355/scan_select_in
+ instance_356/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_366 instance_366/clk_in instance_367/clk_in instance_366/data_in instance_367/data_in
+ instance_366/latch_enable_in instance_367/latch_enable_in instance_366/scan_select_in
+ instance_367/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_377 instance_377/clk_in instance_378/clk_in instance_377/data_in instance_378/data_in
+ instance_377/latch_enable_in instance_378/latch_enable_in instance_377/scan_select_in
+ instance_378/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_130 instance_130/clk_in instance_131/clk_in instance_130/data_in instance_131/data_in
+ instance_130/latch_enable_in instance_131/latch_enable_in instance_130/scan_select_in
+ instance_131/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_141 instance_141/clk_in instance_142/clk_in instance_141/data_in instance_142/data_in
+ instance_141/latch_enable_in instance_142/latch_enable_in instance_141/scan_select_in
+ instance_142/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_152 instance_152/clk_in instance_153/clk_in instance_152/data_in instance_153/data_in
+ instance_152/latch_enable_in instance_153/latch_enable_in instance_152/scan_select_in
+ instance_153/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_163 instance_163/clk_in instance_164/clk_in instance_163/data_in instance_164/data_in
+ instance_163/latch_enable_in instance_164/latch_enable_in instance_163/scan_select_in
+ instance_164/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_174 instance_174/clk_in instance_175/clk_in instance_174/data_in instance_175/data_in
+ instance_174/latch_enable_in instance_175/latch_enable_in instance_174/scan_select_in
+ instance_175/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_185 instance_185/clk_in instance_186/clk_in instance_185/data_in instance_186/data_in
+ instance_185/latch_enable_in instance_186/latch_enable_in instance_185/scan_select_in
+ instance_186/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
Xinstance_196 instance_196/clk_in instance_197/clk_in instance_196/data_in instance_197/data_in
+ instance_196/latch_enable_in instance_197/latch_enable_in instance_196/scan_select_in
+ instance_197/scan_select_in vccd1 vssd1 scan_wrapper_lesson_1
.ends

