magic
tech sky130A
magscale 1 2
timestamp 1656501016
<< obsli1 >>
rect 71104 72159 331860 330425
<< obsm1 >>
rect 68922 68620 580322 524476
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< obsm2 >>
rect 68926 68614 580318 524521
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 583520 298604 584960 298844
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 583520 6476 584960 6716
<< obsm3 >>
rect 68921 524284 583440 524517
rect 68921 511492 583520 524284
rect 68921 511092 583440 511492
rect 68921 498164 583520 511092
rect 68921 497764 583440 498164
rect 68921 484836 583520 497764
rect 68921 484436 583440 484836
rect 68921 471644 583520 484436
rect 68921 471244 583440 471644
rect 68921 458316 583520 471244
rect 68921 457916 583440 458316
rect 68921 444988 583520 457916
rect 68921 444588 583440 444988
rect 68921 431796 583520 444588
rect 68921 431396 583440 431796
rect 68921 418468 583520 431396
rect 68921 418068 583440 418468
rect 68921 405140 583520 418068
rect 68921 404740 583440 405140
rect 68921 391948 583520 404740
rect 68921 391548 583440 391948
rect 68921 378620 583520 391548
rect 68921 378220 583440 378620
rect 68921 365292 583520 378220
rect 68921 364892 583440 365292
rect 68921 352100 583520 364892
rect 68921 351700 583440 352100
rect 68921 338772 583520 351700
rect 68921 338372 583440 338772
rect 68921 325444 583520 338372
rect 68921 325044 583440 325444
rect 68921 312252 583520 325044
rect 68921 311852 583440 312252
rect 68921 298924 583520 311852
rect 68921 298524 583440 298924
rect 68921 285596 583520 298524
rect 68921 285196 583440 285596
rect 68921 272404 583520 285196
rect 68921 272004 583440 272404
rect 68921 259076 583520 272004
rect 68921 258676 583440 259076
rect 68921 245748 583520 258676
rect 68921 245348 583440 245748
rect 68921 232556 583520 245348
rect 68921 232156 583440 232556
rect 68921 219228 583520 232156
rect 68921 218828 583440 219228
rect 68921 205900 583520 218828
rect 68921 205500 583440 205900
rect 68921 192708 583520 205500
rect 68921 192308 583440 192708
rect 68921 179380 583520 192308
rect 68921 178980 583440 179380
rect 68921 166052 583520 178980
rect 68921 165652 583440 166052
rect 68921 152860 583520 165652
rect 68921 152460 583440 152860
rect 68921 139532 583520 152460
rect 68921 139132 583440 139532
rect 68921 126204 583520 139132
rect 68921 125804 583440 126204
rect 68921 113012 583520 125804
rect 68921 112612 583440 113012
rect 68921 99684 583520 112612
rect 68921 99284 583440 99684
rect 68921 86356 583520 99284
rect 68921 85956 583440 86356
rect 68921 73164 583520 85956
rect 68921 72764 583440 73164
rect 68921 72143 583520 72764
<< metal4 >>
rect -2966 -1894 -2346 705830
rect -2006 -934 -1386 704870
rect 1794 -1894 2414 705830
rect 10794 -1894 11414 705830
rect 19794 -1894 20414 705830
rect 28794 -1894 29414 705830
rect 37794 -1894 38414 705830
rect 46794 -1894 47414 705830
rect 55794 -1894 56414 705830
rect 64794 -1894 65414 705830
rect 73794 335000 74414 705830
rect 82794 335000 83414 705830
rect 91794 335000 92414 705830
rect 100794 335000 101414 705830
rect 109794 335000 110414 705830
rect 118794 335000 119414 705830
rect 127794 335000 128414 705830
rect 136794 335000 137414 705830
rect 145794 335000 146414 705830
rect 154794 335000 155414 705830
rect 163794 335000 164414 705830
rect 172794 335000 173414 705830
rect 181794 335000 182414 705830
rect 190794 335000 191414 705830
rect 199794 335000 200414 705830
rect 208794 335000 209414 705830
rect 217794 335000 218414 705830
rect 226794 335000 227414 705830
rect 235794 335000 236414 705830
rect 244794 335000 245414 705830
rect 253794 335000 254414 705830
rect 262794 335000 263414 705830
rect 271794 335000 272414 705830
rect 280794 335000 281414 705830
rect 289794 335000 290414 705830
rect 298794 335000 299414 705830
rect 307794 335000 308414 705830
rect 316794 335000 317414 705830
rect 325794 335000 326414 705830
rect 334794 335000 335414 705830
rect 73794 308000 74414 311000
rect 82794 308000 83414 311000
rect 91794 308000 92414 311000
rect 100794 308000 101414 311000
rect 109794 308000 110414 311000
rect 118794 308000 119414 311000
rect 127794 308000 128414 311000
rect 136794 308000 137414 311000
rect 145794 308000 146414 311000
rect 154794 308000 155414 311000
rect 163794 308000 164414 311000
rect 172794 308000 173414 311000
rect 181794 308000 182414 311000
rect 190794 308000 191414 311000
rect 199794 308000 200414 311000
rect 208794 308000 209414 311000
rect 217794 308000 218414 311000
rect 226794 308000 227414 311000
rect 235794 308000 236414 311000
rect 244794 308000 245414 311000
rect 253794 308000 254414 311000
rect 262794 308000 263414 311000
rect 271794 308000 272414 311000
rect 280794 308000 281414 311000
rect 289794 308000 290414 311000
rect 298794 308000 299414 311000
rect 307794 308000 308414 311000
rect 316794 308000 317414 311000
rect 325794 308000 326414 311000
rect 334794 308000 335414 311000
rect 73794 281000 74414 284000
rect 82794 281000 83414 284000
rect 91794 281000 92414 284000
rect 100794 281000 101414 284000
rect 109794 281000 110414 284000
rect 118794 281000 119414 284000
rect 127794 281000 128414 284000
rect 136794 281000 137414 284000
rect 145794 281000 146414 284000
rect 154794 281000 155414 284000
rect 163794 281000 164414 284000
rect 172794 281000 173414 284000
rect 181794 281000 182414 284000
rect 190794 281000 191414 284000
rect 199794 281000 200414 284000
rect 208794 281000 209414 284000
rect 217794 281000 218414 284000
rect 226794 281000 227414 284000
rect 235794 281000 236414 284000
rect 244794 281000 245414 284000
rect 253794 281000 254414 284000
rect 262794 281000 263414 284000
rect 271794 281000 272414 284000
rect 280794 281000 281414 284000
rect 289794 281000 290414 284000
rect 298794 281000 299414 284000
rect 307794 281000 308414 284000
rect 316794 281000 317414 284000
rect 325794 281000 326414 284000
rect 334794 281000 335414 284000
rect 73794 254000 74414 257000
rect 82794 254000 83414 257000
rect 91794 254000 92414 257000
rect 100794 254000 101414 257000
rect 109794 254000 110414 257000
rect 118794 254000 119414 257000
rect 127794 254000 128414 257000
rect 136794 254000 137414 257000
rect 145794 254000 146414 257000
rect 154794 254000 155414 257000
rect 163794 254000 164414 257000
rect 172794 254000 173414 257000
rect 181794 254000 182414 257000
rect 190794 254000 191414 257000
rect 199794 254000 200414 257000
rect 208794 254000 209414 257000
rect 217794 254000 218414 257000
rect 226794 254000 227414 257000
rect 235794 254000 236414 257000
rect 244794 254000 245414 257000
rect 253794 254000 254414 257000
rect 262794 254000 263414 257000
rect 271794 254000 272414 257000
rect 280794 254000 281414 257000
rect 289794 254000 290414 257000
rect 298794 254000 299414 257000
rect 307794 254000 308414 257000
rect 316794 254000 317414 257000
rect 325794 254000 326414 257000
rect 334794 254000 335414 257000
rect 73794 227000 74414 230000
rect 82794 227000 83414 230000
rect 91794 227000 92414 230000
rect 100794 227000 101414 230000
rect 109794 227000 110414 230000
rect 118794 227000 119414 230000
rect 127794 227000 128414 230000
rect 136794 227000 137414 230000
rect 145794 227000 146414 230000
rect 154794 227000 155414 230000
rect 163794 227000 164414 230000
rect 172794 227000 173414 230000
rect 181794 227000 182414 230000
rect 190794 227000 191414 230000
rect 199794 227000 200414 230000
rect 208794 227000 209414 230000
rect 217794 227000 218414 230000
rect 226794 227000 227414 230000
rect 235794 227000 236414 230000
rect 244794 227000 245414 230000
rect 253794 227000 254414 230000
rect 262794 227000 263414 230000
rect 271794 227000 272414 230000
rect 280794 227000 281414 230000
rect 289794 227000 290414 230000
rect 298794 227000 299414 230000
rect 307794 227000 308414 230000
rect 316794 227000 317414 230000
rect 325794 227000 326414 230000
rect 334794 227000 335414 230000
rect 73794 200000 74414 203000
rect 82794 200000 83414 203000
rect 91794 200000 92414 203000
rect 100794 200000 101414 203000
rect 109794 200000 110414 203000
rect 118794 200000 119414 203000
rect 127794 200000 128414 203000
rect 136794 200000 137414 203000
rect 145794 200000 146414 203000
rect 154794 200000 155414 203000
rect 163794 200000 164414 203000
rect 172794 200000 173414 203000
rect 181794 200000 182414 203000
rect 190794 200000 191414 203000
rect 199794 200000 200414 203000
rect 208794 200000 209414 203000
rect 217794 200000 218414 203000
rect 226794 200000 227414 203000
rect 235794 200000 236414 203000
rect 244794 200000 245414 203000
rect 253794 200000 254414 203000
rect 262794 200000 263414 203000
rect 271794 200000 272414 203000
rect 280794 200000 281414 203000
rect 289794 200000 290414 203000
rect 298794 200000 299414 203000
rect 307794 200000 308414 203000
rect 316794 200000 317414 203000
rect 325794 200000 326414 203000
rect 334794 200000 335414 203000
rect 73794 173000 74414 176000
rect 82794 173000 83414 176000
rect 91794 173000 92414 176000
rect 100794 173000 101414 176000
rect 109794 173000 110414 176000
rect 118794 173000 119414 176000
rect 127794 173000 128414 176000
rect 136794 173000 137414 176000
rect 145794 173000 146414 176000
rect 154794 173000 155414 176000
rect 163794 173000 164414 176000
rect 172794 173000 173414 176000
rect 181794 173000 182414 176000
rect 190794 173000 191414 176000
rect 199794 173000 200414 176000
rect 208794 173000 209414 176000
rect 217794 173000 218414 176000
rect 226794 173000 227414 176000
rect 235794 173000 236414 176000
rect 244794 173000 245414 176000
rect 253794 173000 254414 176000
rect 262794 173000 263414 176000
rect 271794 173000 272414 176000
rect 280794 173000 281414 176000
rect 289794 173000 290414 176000
rect 298794 173000 299414 176000
rect 307794 173000 308414 176000
rect 316794 173000 317414 176000
rect 325794 173000 326414 176000
rect 334794 173000 335414 176000
rect 73794 146000 74414 149000
rect 82794 146000 83414 149000
rect 91794 146000 92414 149000
rect 100794 146000 101414 149000
rect 109794 146000 110414 149000
rect 118794 146000 119414 149000
rect 127794 146000 128414 149000
rect 136794 146000 137414 149000
rect 145794 146000 146414 149000
rect 154794 146000 155414 149000
rect 163794 146000 164414 149000
rect 172794 146000 173414 149000
rect 181794 146000 182414 149000
rect 190794 146000 191414 149000
rect 199794 146000 200414 149000
rect 208794 146000 209414 149000
rect 217794 146000 218414 149000
rect 226794 146000 227414 149000
rect 235794 146000 236414 149000
rect 244794 146000 245414 149000
rect 253794 146000 254414 149000
rect 262794 146000 263414 149000
rect 271794 146000 272414 149000
rect 280794 146000 281414 149000
rect 289794 146000 290414 149000
rect 298794 146000 299414 149000
rect 307794 146000 308414 149000
rect 316794 146000 317414 149000
rect 325794 146000 326414 149000
rect 334794 146000 335414 149000
rect 73794 119000 74414 122000
rect 82794 119000 83414 122000
rect 91794 119000 92414 122000
rect 100794 119000 101414 122000
rect 109794 119000 110414 122000
rect 118794 119000 119414 122000
rect 127794 119000 128414 122000
rect 136794 119000 137414 122000
rect 145794 119000 146414 122000
rect 154794 119000 155414 122000
rect 163794 119000 164414 122000
rect 172794 119000 173414 122000
rect 181794 119000 182414 122000
rect 190794 119000 191414 122000
rect 199794 119000 200414 122000
rect 208794 119000 209414 122000
rect 217794 119000 218414 122000
rect 226794 119000 227414 122000
rect 235794 119000 236414 122000
rect 244794 119000 245414 122000
rect 253794 119000 254414 122000
rect 262794 119000 263414 122000
rect 271794 119000 272414 122000
rect 280794 119000 281414 122000
rect 289794 119000 290414 122000
rect 298794 119000 299414 122000
rect 307794 119000 308414 122000
rect 316794 119000 317414 122000
rect 325794 119000 326414 122000
rect 334794 119000 335414 122000
rect 73794 92000 74414 95000
rect 82794 92000 83414 95000
rect 91794 92000 92414 95000
rect 100794 92000 101414 95000
rect 109794 92000 110414 95000
rect 118794 92000 119414 95000
rect 127794 92000 128414 95000
rect 136794 92000 137414 95000
rect 145794 92000 146414 95000
rect 154794 92000 155414 95000
rect 163794 92000 164414 95000
rect 172794 92000 173414 95000
rect 181794 92000 182414 95000
rect 190794 92000 191414 95000
rect 199794 92000 200414 95000
rect 208794 92000 209414 95000
rect 217794 92000 218414 95000
rect 226794 92000 227414 95000
rect 235794 92000 236414 95000
rect 244794 92000 245414 95000
rect 253794 92000 254414 95000
rect 262794 92000 263414 95000
rect 271794 92000 272414 95000
rect 280794 92000 281414 95000
rect 289794 92000 290414 95000
rect 298794 92000 299414 95000
rect 307794 92000 308414 95000
rect 316794 92000 317414 95000
rect 325794 92000 326414 95000
rect 334794 92000 335414 95000
rect 73794 -1894 74414 68000
rect 82794 -1894 83414 68000
rect 91794 -1894 92414 68000
rect 100794 -1894 101414 68000
rect 109794 -1894 110414 68000
rect 118794 -1894 119414 68000
rect 127794 -1894 128414 68000
rect 136794 -1894 137414 68000
rect 145794 -1894 146414 68000
rect 154794 -1894 155414 68000
rect 163794 -1894 164414 68000
rect 172794 -1894 173414 68000
rect 181794 -1894 182414 68000
rect 190794 -1894 191414 68000
rect 199794 -1894 200414 68000
rect 208794 -1894 209414 68000
rect 217794 -1894 218414 68000
rect 226794 -1894 227414 68000
rect 235794 -1894 236414 68000
rect 244794 -1894 245414 68000
rect 253794 -1894 254414 68000
rect 262794 -1894 263414 68000
rect 271794 -1894 272414 68000
rect 280794 -1894 281414 68000
rect 289794 -1894 290414 68000
rect 298794 -1894 299414 68000
rect 307794 -1894 308414 68000
rect 316794 -1894 317414 68000
rect 325794 -1894 326414 68000
rect 334794 -1894 335414 68000
rect 343794 -1894 344414 705830
rect 352794 -1894 353414 705830
rect 361794 -1894 362414 705830
rect 370794 -1894 371414 705830
rect 379794 -1894 380414 705830
rect 388794 -1894 389414 705830
rect 397794 -1894 398414 705830
rect 406794 -1894 407414 705830
rect 415794 -1894 416414 705830
rect 424794 -1894 425414 705830
rect 433794 -1894 434414 705830
rect 442794 -1894 443414 705830
rect 451794 -1894 452414 705830
rect 460794 -1894 461414 705830
rect 469794 -1894 470414 705830
rect 478794 -1894 479414 705830
rect 487794 -1894 488414 705830
rect 496794 -1894 497414 705830
rect 505794 -1894 506414 705830
rect 514794 -1894 515414 705830
rect 523794 -1894 524414 705830
rect 532794 -1894 533414 705830
rect 541794 -1894 542414 705830
rect 550794 -1894 551414 705830
rect 559794 -1894 560414 705830
rect 568794 -1894 569414 705830
rect 577794 -1894 578414 705830
rect 585310 -934 585930 704870
rect 586270 -1894 586890 705830
<< obsm4 >>
rect 73910 311080 329091 330456
rect 74494 307920 82714 311080
rect 83494 307920 91714 311080
rect 92494 307920 100714 311080
rect 101494 307920 109714 311080
rect 110494 307920 118714 311080
rect 119494 307920 127714 311080
rect 128494 307920 136714 311080
rect 137494 307920 145714 311080
rect 146494 307920 154714 311080
rect 155494 307920 163714 311080
rect 164494 307920 172714 311080
rect 173494 307920 181714 311080
rect 182494 307920 190714 311080
rect 191494 307920 199714 311080
rect 200494 307920 208714 311080
rect 209494 307920 217714 311080
rect 218494 307920 226714 311080
rect 227494 307920 235714 311080
rect 236494 307920 244714 311080
rect 245494 307920 253714 311080
rect 254494 307920 262714 311080
rect 263494 307920 271714 311080
rect 272494 307920 280714 311080
rect 281494 307920 289714 311080
rect 290494 307920 298714 311080
rect 299494 307920 307714 311080
rect 308494 307920 316714 311080
rect 317494 307920 325714 311080
rect 326494 307920 329091 311080
rect 73910 284080 329091 307920
rect 74494 280920 82714 284080
rect 83494 280920 91714 284080
rect 92494 280920 100714 284080
rect 101494 280920 109714 284080
rect 110494 280920 118714 284080
rect 119494 280920 127714 284080
rect 128494 280920 136714 284080
rect 137494 280920 145714 284080
rect 146494 280920 154714 284080
rect 155494 280920 163714 284080
rect 164494 280920 172714 284080
rect 173494 280920 181714 284080
rect 182494 280920 190714 284080
rect 191494 280920 199714 284080
rect 200494 280920 208714 284080
rect 209494 280920 217714 284080
rect 218494 280920 226714 284080
rect 227494 280920 235714 284080
rect 236494 280920 244714 284080
rect 245494 280920 253714 284080
rect 254494 280920 262714 284080
rect 263494 280920 271714 284080
rect 272494 280920 280714 284080
rect 281494 280920 289714 284080
rect 290494 280920 298714 284080
rect 299494 280920 307714 284080
rect 308494 280920 316714 284080
rect 317494 280920 325714 284080
rect 326494 280920 329091 284080
rect 73910 257080 329091 280920
rect 74494 253920 82714 257080
rect 83494 253920 91714 257080
rect 92494 253920 100714 257080
rect 101494 253920 109714 257080
rect 110494 253920 118714 257080
rect 119494 253920 127714 257080
rect 128494 253920 136714 257080
rect 137494 253920 145714 257080
rect 146494 253920 154714 257080
rect 155494 253920 163714 257080
rect 164494 253920 172714 257080
rect 173494 253920 181714 257080
rect 182494 253920 190714 257080
rect 191494 253920 199714 257080
rect 200494 253920 208714 257080
rect 209494 253920 217714 257080
rect 218494 253920 226714 257080
rect 227494 253920 235714 257080
rect 236494 253920 244714 257080
rect 245494 253920 253714 257080
rect 254494 253920 262714 257080
rect 263494 253920 271714 257080
rect 272494 253920 280714 257080
rect 281494 253920 289714 257080
rect 290494 253920 298714 257080
rect 299494 253920 307714 257080
rect 308494 253920 316714 257080
rect 317494 253920 325714 257080
rect 326494 253920 329091 257080
rect 73910 230080 329091 253920
rect 74494 226920 82714 230080
rect 83494 226920 91714 230080
rect 92494 226920 100714 230080
rect 101494 226920 109714 230080
rect 110494 226920 118714 230080
rect 119494 226920 127714 230080
rect 128494 226920 136714 230080
rect 137494 226920 145714 230080
rect 146494 226920 154714 230080
rect 155494 226920 163714 230080
rect 164494 226920 172714 230080
rect 173494 226920 181714 230080
rect 182494 226920 190714 230080
rect 191494 226920 199714 230080
rect 200494 226920 208714 230080
rect 209494 226920 217714 230080
rect 218494 226920 226714 230080
rect 227494 226920 235714 230080
rect 236494 226920 244714 230080
rect 245494 226920 253714 230080
rect 254494 226920 262714 230080
rect 263494 226920 271714 230080
rect 272494 226920 280714 230080
rect 281494 226920 289714 230080
rect 290494 226920 298714 230080
rect 299494 226920 307714 230080
rect 308494 226920 316714 230080
rect 317494 226920 325714 230080
rect 326494 226920 329091 230080
rect 73910 203080 329091 226920
rect 74494 199920 82714 203080
rect 83494 199920 91714 203080
rect 92494 199920 100714 203080
rect 101494 199920 109714 203080
rect 110494 199920 118714 203080
rect 119494 199920 127714 203080
rect 128494 199920 136714 203080
rect 137494 199920 145714 203080
rect 146494 199920 154714 203080
rect 155494 199920 163714 203080
rect 164494 199920 172714 203080
rect 173494 199920 181714 203080
rect 182494 199920 190714 203080
rect 191494 199920 199714 203080
rect 200494 199920 208714 203080
rect 209494 199920 217714 203080
rect 218494 199920 226714 203080
rect 227494 199920 235714 203080
rect 236494 199920 244714 203080
rect 245494 199920 253714 203080
rect 254494 199920 262714 203080
rect 263494 199920 271714 203080
rect 272494 199920 280714 203080
rect 281494 199920 289714 203080
rect 290494 199920 298714 203080
rect 299494 199920 307714 203080
rect 308494 199920 316714 203080
rect 317494 199920 325714 203080
rect 326494 199920 329091 203080
rect 73910 176080 329091 199920
rect 74494 172920 82714 176080
rect 83494 172920 91714 176080
rect 92494 172920 100714 176080
rect 101494 172920 109714 176080
rect 110494 172920 118714 176080
rect 119494 172920 127714 176080
rect 128494 172920 136714 176080
rect 137494 172920 145714 176080
rect 146494 172920 154714 176080
rect 155494 172920 163714 176080
rect 164494 172920 172714 176080
rect 173494 172920 181714 176080
rect 182494 172920 190714 176080
rect 191494 172920 199714 176080
rect 200494 172920 208714 176080
rect 209494 172920 217714 176080
rect 218494 172920 226714 176080
rect 227494 172920 235714 176080
rect 236494 172920 244714 176080
rect 245494 172920 253714 176080
rect 254494 172920 262714 176080
rect 263494 172920 271714 176080
rect 272494 172920 280714 176080
rect 281494 172920 289714 176080
rect 290494 172920 298714 176080
rect 299494 172920 307714 176080
rect 308494 172920 316714 176080
rect 317494 172920 325714 176080
rect 326494 172920 329091 176080
rect 73910 149080 329091 172920
rect 74494 145920 82714 149080
rect 83494 145920 91714 149080
rect 92494 145920 100714 149080
rect 101494 145920 109714 149080
rect 110494 145920 118714 149080
rect 119494 145920 127714 149080
rect 128494 145920 136714 149080
rect 137494 145920 145714 149080
rect 146494 145920 154714 149080
rect 155494 145920 163714 149080
rect 164494 145920 172714 149080
rect 173494 145920 181714 149080
rect 182494 145920 190714 149080
rect 191494 145920 199714 149080
rect 200494 145920 208714 149080
rect 209494 145920 217714 149080
rect 218494 145920 226714 149080
rect 227494 145920 235714 149080
rect 236494 145920 244714 149080
rect 245494 145920 253714 149080
rect 254494 145920 262714 149080
rect 263494 145920 271714 149080
rect 272494 145920 280714 149080
rect 281494 145920 289714 149080
rect 290494 145920 298714 149080
rect 299494 145920 307714 149080
rect 308494 145920 316714 149080
rect 317494 145920 325714 149080
rect 326494 145920 329091 149080
rect 73910 122080 329091 145920
rect 74494 118920 82714 122080
rect 83494 118920 91714 122080
rect 92494 118920 100714 122080
rect 101494 118920 109714 122080
rect 110494 118920 118714 122080
rect 119494 118920 127714 122080
rect 128494 118920 136714 122080
rect 137494 118920 145714 122080
rect 146494 118920 154714 122080
rect 155494 118920 163714 122080
rect 164494 118920 172714 122080
rect 173494 118920 181714 122080
rect 182494 118920 190714 122080
rect 191494 118920 199714 122080
rect 200494 118920 208714 122080
rect 209494 118920 217714 122080
rect 218494 118920 226714 122080
rect 227494 118920 235714 122080
rect 236494 118920 244714 122080
rect 245494 118920 253714 122080
rect 254494 118920 262714 122080
rect 263494 118920 271714 122080
rect 272494 118920 280714 122080
rect 281494 118920 289714 122080
rect 290494 118920 298714 122080
rect 299494 118920 307714 122080
rect 308494 118920 316714 122080
rect 317494 118920 325714 122080
rect 326494 118920 329091 122080
rect 73910 95080 329091 118920
rect 74494 91920 82714 95080
rect 83494 91920 91714 95080
rect 92494 91920 100714 95080
rect 101494 91920 109714 95080
rect 110494 91920 118714 95080
rect 119494 91920 127714 95080
rect 128494 91920 136714 95080
rect 137494 91920 145714 95080
rect 146494 91920 154714 95080
rect 155494 91920 163714 95080
rect 164494 91920 172714 95080
rect 173494 91920 181714 95080
rect 182494 91920 190714 95080
rect 191494 91920 199714 95080
rect 200494 91920 208714 95080
rect 209494 91920 217714 95080
rect 218494 91920 226714 95080
rect 227494 91920 235714 95080
rect 236494 91920 244714 95080
rect 245494 91920 253714 95080
rect 254494 91920 262714 95080
rect 263494 91920 271714 95080
rect 272494 91920 280714 95080
rect 281494 91920 289714 95080
rect 290494 91920 298714 95080
rect 299494 91920 307714 95080
rect 308494 91920 316714 95080
rect 317494 91920 325714 95080
rect 326494 91920 329091 95080
rect 73910 72128 329091 91920
<< metal5 >>
rect -2966 705210 586890 705830
rect -2006 704250 585930 704870
rect -2966 695866 586890 696486
rect -2966 686866 586890 687486
rect -2966 677866 586890 678486
rect -2966 668866 586890 669486
rect -2966 659866 586890 660486
rect -2966 650866 586890 651486
rect -2966 641866 586890 642486
rect -2966 632866 586890 633486
rect -2966 623866 586890 624486
rect -2966 614866 586890 615486
rect -2966 605866 586890 606486
rect -2966 596866 586890 597486
rect -2966 587866 586890 588486
rect -2966 578866 586890 579486
rect -2966 569866 586890 570486
rect -2966 560866 586890 561486
rect -2966 551866 586890 552486
rect -2966 542866 586890 543486
rect -2966 533866 586890 534486
rect -2966 524866 586890 525486
rect -2966 515866 586890 516486
rect -2966 506866 586890 507486
rect -2966 497866 586890 498486
rect -2966 488866 586890 489486
rect -2966 479866 586890 480486
rect -2966 470866 586890 471486
rect -2966 461866 586890 462486
rect -2966 452866 586890 453486
rect -2966 443866 586890 444486
rect -2966 434866 586890 435486
rect -2966 425866 586890 426486
rect -2966 416866 586890 417486
rect -2966 407866 586890 408486
rect -2966 398866 586890 399486
rect -2966 389866 586890 390486
rect -2966 380866 586890 381486
rect -2966 371866 586890 372486
rect -2966 362866 586890 363486
rect -2966 353866 586890 354486
rect -2966 344866 586890 345486
rect -2966 335866 586890 336486
rect -2966 326866 586890 327486
rect -2966 317866 586890 318486
rect 82794 309806 335414 310426
rect -2966 308866 586890 309486
rect -2966 299866 586890 300486
rect -2966 290866 586890 291486
rect 73794 282806 326414 283426
rect -2966 281866 586890 282486
rect -2966 272866 586890 273486
rect -2966 263866 586890 264486
rect 82794 255806 335414 256426
rect -2966 254866 586890 255486
rect -2966 245866 586890 246486
rect -2966 236866 586890 237486
rect 73794 228806 326414 229426
rect -2966 227866 586890 228486
rect -2966 218866 586890 219486
rect -2966 209866 586890 210486
rect 82794 201806 335414 202426
rect -2966 200866 586890 201486
rect -2966 191866 586890 192486
rect -2966 182866 586890 183486
rect 73794 174806 326414 175426
rect -2966 173866 586890 174486
rect -2966 164866 586890 165486
rect -2966 155866 586890 156486
rect 82794 147806 335414 148426
rect -2966 146866 586890 147486
rect -2966 137866 586890 138486
rect -2966 128866 586890 129486
rect 73794 120806 326414 121426
rect -2966 119866 586890 120486
rect -2966 110866 586890 111486
rect -2966 101866 586890 102486
rect 82794 93806 335414 94426
rect -2966 92866 586890 93486
rect -2966 83866 586890 84486
rect -2966 74866 586890 75486
rect -2966 65866 586890 66486
rect -2966 56866 586890 57486
rect -2966 47866 586890 48486
rect -2966 38866 586890 39486
rect -2966 29866 586890 30486
rect -2966 20866 586890 21486
rect -2966 11866 586890 12486
rect -2966 2866 586890 3486
rect -2006 -934 585930 -314
rect -2966 -1894 586890 -1274
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 46 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 47 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 48 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 49 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 50 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 51 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 53 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 54 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 55 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 56 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 57 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 58 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 59 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 60 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 122 nsew signal output
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 123 nsew signal output
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 124 nsew signal output
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 125 nsew signal output
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 126 nsew signal output
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 127 nsew signal output
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 129 nsew signal output
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 130 nsew signal output
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 131 nsew signal output
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 132 nsew signal output
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 133 nsew signal output
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 134 nsew signal output
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 135 nsew signal output
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 136 nsew signal output
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 528 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 531 nsew signal output
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 532 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 20866 586890 21486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 56866 586890 57486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 92866 586890 93486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 532 nsew power input
rlabel metal5 s 73794 120806 326414 121426 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 128866 586890 129486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 164866 586890 165486 6 vccd1
port 532 nsew power input
rlabel metal5 s 73794 174806 326414 175426 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 200866 586890 201486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 532 nsew power input
rlabel metal5 s 73794 228806 326414 229426 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 236866 586890 237486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 272866 586890 273486 6 vccd1
port 532 nsew power input
rlabel metal5 s 73794 282806 326414 283426 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 308866 586890 309486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 344866 586890 345486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 380866 586890 381486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 416866 586890 417486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 452866 586890 453486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 488866 586890 489486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 524866 586890 525486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 560866 586890 561486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 596866 586890 597486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 632866 586890 633486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 668866 586890 669486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 -1894 74414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 -1894 92414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 -1894 110414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 -1894 128414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 -1894 146414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 -1894 164414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 -1894 182414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 -1894 200414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 -1894 218414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 -1894 236414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 -1894 254414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 -1894 272414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 -1894 290414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 -1894 308414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 -1894 326414 68000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 92000 74414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 92000 92414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 92000 110414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 92000 128414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 92000 146414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 92000 164414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 92000 182414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 92000 200414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 92000 218414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 92000 236414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 92000 254414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 92000 272414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 92000 290414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 92000 308414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 92000 326414 95000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 119000 74414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 119000 92414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 119000 110414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 119000 128414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 119000 146414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 119000 164414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 119000 182414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 119000 200414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 119000 218414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 119000 236414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 119000 254414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 119000 272414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 119000 290414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 119000 308414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 119000 326414 122000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 146000 74414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 146000 92414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 146000 110414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 146000 128414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 146000 146414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 146000 164414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 146000 182414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 146000 200414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 146000 218414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 146000 236414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 146000 254414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 146000 272414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 146000 290414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 146000 308414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 146000 326414 149000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 173000 74414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 173000 92414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 173000 110414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 173000 128414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 173000 146414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 173000 164414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 173000 182414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 173000 200414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 173000 218414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 173000 236414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 173000 254414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 173000 272414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 173000 290414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 173000 308414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 173000 326414 176000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 200000 74414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 200000 92414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 200000 110414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 200000 128414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 200000 146414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 200000 164414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 200000 182414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 200000 200414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 200000 218414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 200000 236414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 200000 254414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 200000 272414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 200000 290414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 200000 308414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 200000 326414 203000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 227000 74414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 227000 92414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 227000 110414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 227000 128414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 227000 146414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 227000 164414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 227000 182414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 227000 200414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 227000 218414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 227000 236414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 227000 254414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 227000 272414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 227000 290414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 227000 308414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 227000 326414 230000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 254000 74414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 254000 92414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 254000 110414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 254000 128414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 254000 146414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 254000 164414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 254000 182414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 254000 200414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 254000 218414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 254000 236414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 254000 254414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 254000 272414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 254000 290414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 254000 308414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 254000 326414 257000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 281000 74414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 281000 92414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 281000 110414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 281000 128414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 281000 146414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 281000 164414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 281000 182414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 281000 200414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 281000 218414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 281000 236414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 281000 254414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 281000 272414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 281000 290414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 281000 308414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 281000 326414 284000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 308000 74414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 308000 92414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 308000 110414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 308000 128414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 308000 146414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 308000 164414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 308000 182414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 308000 200414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 308000 218414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 308000 236414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 308000 254414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 308000 272414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 308000 290414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 308000 308414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 308000 326414 311000 6 vccd1
port 532 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 532 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 532 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 19794 -1894 20414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 55794 -1894 56414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 335000 74414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 91794 335000 92414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 335000 110414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 127794 335000 128414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 335000 146414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 163794 335000 164414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 335000 182414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 199794 335000 200414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 335000 218414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 235794 335000 236414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 335000 254414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 271794 335000 272414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 335000 290414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 307794 335000 308414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 335000 326414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 343794 -1894 344414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 379794 -1894 380414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 415794 -1894 416414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 451794 -1894 452414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 487794 -1894 488414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 523794 -1894 524414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 559794 -1894 560414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 11866 586890 12486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 29866 586890 30486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 47866 586890 48486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 65866 586890 66486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 83866 586890 84486 6 vssd1
port 533 nsew ground input
rlabel metal5 s 82794 93806 335414 94426 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 101866 586890 102486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 119866 586890 120486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 137866 586890 138486 6 vssd1
port 533 nsew ground input
rlabel metal5 s 82794 147806 335414 148426 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 155866 586890 156486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 173866 586890 174486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 191866 586890 192486 6 vssd1
port 533 nsew ground input
rlabel metal5 s 82794 201806 335414 202426 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 209866 586890 210486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 227866 586890 228486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 245866 586890 246486 6 vssd1
port 533 nsew ground input
rlabel metal5 s 82794 255806 335414 256426 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 263866 586890 264486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 281866 586890 282486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 299866 586890 300486 6 vssd1
port 533 nsew ground input
rlabel metal5 s 82794 309806 335414 310426 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 317866 586890 318486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 335866 586890 336486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 353866 586890 354486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 371866 586890 372486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 389866 586890 390486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 407866 586890 408486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 425866 586890 426486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 443866 586890 444486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 461866 586890 462486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 479866 586890 480486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 497866 586890 498486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 515866 586890 516486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 533866 586890 534486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 551866 586890 552486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 569866 586890 570486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 587866 586890 588486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 605866 586890 606486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 623866 586890 624486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 641866 586890 642486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 659866 586890 660486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 677866 586890 678486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 695866 586890 696486 6 vssd1
port 533 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 -1894 83414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 -1894 101414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 -1894 119414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 -1894 137414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 -1894 155414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 -1894 173414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 -1894 191414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 -1894 209414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 -1894 227414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 -1894 245414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 -1894 263414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 -1894 281414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 -1894 299414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 -1894 317414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 -1894 335414 68000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 92000 83414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 92000 101414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 92000 119414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 92000 137414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 92000 155414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 92000 173414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 92000 191414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 92000 209414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 92000 227414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 92000 245414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 92000 263414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 92000 281414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 92000 299414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 92000 317414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 92000 335414 95000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 119000 83414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 119000 101414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 119000 119414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 119000 137414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 119000 155414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 119000 173414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 119000 191414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 119000 209414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 119000 227414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 119000 245414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 119000 263414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 119000 281414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 119000 299414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 119000 317414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 119000 335414 122000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 146000 83414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 146000 101414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 146000 119414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 146000 137414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 146000 155414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 146000 173414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 146000 191414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 146000 209414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 146000 227414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 146000 245414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 146000 263414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 146000 281414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 146000 299414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 146000 317414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 146000 335414 149000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 173000 83414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 173000 101414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 173000 119414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 173000 137414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 173000 155414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 173000 173414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 173000 191414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 173000 209414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 173000 227414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 173000 245414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 173000 263414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 173000 281414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 173000 299414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 173000 317414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 173000 335414 176000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 200000 83414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 200000 101414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 200000 119414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 200000 137414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 200000 155414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 200000 173414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 200000 191414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 200000 209414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 200000 227414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 200000 245414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 200000 263414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 200000 281414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 200000 299414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 200000 317414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 200000 335414 203000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 227000 83414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 227000 101414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 227000 119414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 227000 137414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 227000 155414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 227000 173414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 227000 191414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 227000 209414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 227000 227414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 227000 245414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 227000 263414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 227000 281414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 227000 299414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 227000 317414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 227000 335414 230000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 254000 83414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 254000 101414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 254000 119414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 254000 137414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 254000 155414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 254000 173414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 254000 191414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 254000 209414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 254000 227414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 254000 245414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 254000 263414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 254000 281414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 254000 299414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 254000 317414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 254000 335414 257000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 281000 83414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 281000 101414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 281000 119414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 281000 137414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 281000 155414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 281000 173414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 281000 191414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 281000 209414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 281000 227414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 281000 245414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 281000 263414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 281000 281414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 281000 299414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 281000 317414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 281000 335414 284000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 308000 83414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 308000 101414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 308000 119414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 308000 137414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 308000 155414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 308000 173414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 308000 191414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 308000 209414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 308000 227414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 308000 245414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 308000 263414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 308000 281414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 308000 299414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 308000 317414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 308000 335414 311000 6 vssd1
port 533 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 533 nsew ground input
rlabel metal4 s 10794 -1894 11414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 28794 -1894 29414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 46794 -1894 47414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 64794 -1894 65414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 82794 335000 83414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 100794 335000 101414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 118794 335000 119414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 136794 335000 137414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 154794 335000 155414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 172794 335000 173414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 190794 335000 191414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 208794 335000 209414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 226794 335000 227414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 244794 335000 245414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 262794 335000 263414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 280794 335000 281414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 298794 335000 299414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 316794 335000 317414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 334794 335000 335414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 352794 -1894 353414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 370794 -1894 371414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 388794 -1894 389414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 406794 -1894 407414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 424794 -1894 425414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 442794 -1894 443414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 460794 -1894 461414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 478794 -1894 479414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 496794 -1894 497414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 514794 -1894 515414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 532794 -1894 533414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 550794 -1894 551414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 568794 -1894 569414 705830 6 vssd1
port 533 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 533 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 534 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 535 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 536 nsew signal output
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 537 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 538 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 539 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 540 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 541 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 542 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 543 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 544 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 545 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 546 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 547 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 548 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 549 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 550 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 551 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 552 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 553 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 554 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 555 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 556 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 557 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 558 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 559 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 560 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 561 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 562 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 563 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 564 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 565 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 566 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 567 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 568 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 569 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 570 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 571 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 572 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 573 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 574 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 575 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 576 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 577 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 578 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 579 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 580 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 581 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 582 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 583 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 584 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 585 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 586 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 587 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 588 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 589 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 590 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 591 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 592 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 593 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 594 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 595 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 596 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 597 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 598 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 599 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 600 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 601 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 602 nsew signal output
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 603 nsew signal output
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 604 nsew signal output
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 605 nsew signal output
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 606 nsew signal output
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 607 nsew signal output
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 608 nsew signal output
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 609 nsew signal output
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 610 nsew signal output
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 611 nsew signal output
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 612 nsew signal output
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 613 nsew signal output
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 614 nsew signal output
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 615 nsew signal output
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 616 nsew signal output
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 617 nsew signal output
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 618 nsew signal output
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 619 nsew signal output
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 620 nsew signal output
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 621 nsew signal output
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 622 nsew signal output
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 623 nsew signal output
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 624 nsew signal output
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 625 nsew signal output
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 626 nsew signal output
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 627 nsew signal output
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 628 nsew signal output
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 629 nsew signal output
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 630 nsew signal output
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 631 nsew signal output
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 632 nsew signal output
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 633 nsew signal output
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 634 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 635 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 636 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 637 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 638 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 639 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1785376
string GDS_FILE /home/matt/work/asic-workshop/shuttle6/tapeout_100/openlane/user_project_wrapper/runs/user_project_wrapper/results/finishing/user_project_wrapper.magic.gds
string GDS_START 321136
<< end >>

