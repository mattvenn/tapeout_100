magic
tech sky130A
magscale 1 2
timestamp 1656501897
<< metal1 >>
rect 25958 686128 25964 686180
rect 26016 686168 26022 686180
rect 149698 686168 149704 686180
rect 26016 686140 149704 686168
rect 26016 686128 26022 686140
rect 149698 686128 149704 686140
rect 149756 686128 149762 686180
rect 36630 686060 36636 686112
rect 36688 686100 36694 686112
rect 52454 686100 52460 686112
rect 36688 686072 52460 686100
rect 36688 686060 36694 686072
rect 52454 686060 52460 686072
rect 52512 686060 52518 686112
rect 232314 686060 232320 686112
rect 232372 686100 232378 686112
rect 251818 686100 251824 686112
rect 232372 686072 251824 686100
rect 232372 686060 232378 686072
rect 251818 686060 251824 686072
rect 251876 686060 251882 686112
rect 62482 685992 62488 686044
rect 62540 686032 62546 686044
rect 79318 686032 79324 686044
rect 62540 686004 79324 686032
rect 62540 685992 62546 686004
rect 79318 685992 79324 686004
rect 79376 685992 79382 686044
rect 90358 685992 90364 686044
rect 90416 686032 90422 686044
rect 106366 686032 106372 686044
rect 90416 686004 106372 686032
rect 90416 685992 90422 686004
rect 106366 685992 106372 686004
rect 106424 685992 106430 686044
rect 116486 685992 116492 686044
rect 116544 686032 116550 686044
rect 133414 686032 133420 686044
rect 116544 686004 133420 686032
rect 116544 685992 116550 686004
rect 133414 685992 133420 686004
rect 133472 685992 133478 686044
rect 144270 685992 144276 686044
rect 144328 686032 144334 686044
rect 160278 686032 160284 686044
rect 144328 686004 160284 686032
rect 144328 685992 144334 686004
rect 160278 685992 160284 686004
rect 160336 685992 160342 686044
rect 170490 685992 170496 686044
rect 170548 686032 170554 686044
rect 187786 686032 187792 686044
rect 170548 686004 187792 686032
rect 170548 685992 170554 686004
rect 187786 685992 187792 686004
rect 187844 685992 187850 686044
rect 197538 685992 197544 686044
rect 197596 686032 197602 686044
rect 214374 686032 214380 686044
rect 197596 686004 214380 686032
rect 197596 685992 197602 686004
rect 214374 685992 214380 686004
rect 214432 685992 214438 686044
rect 224494 685992 224500 686044
rect 224552 686032 224558 686044
rect 241514 686032 241520 686044
rect 224552 686004 241520 686032
rect 224552 685992 224558 686004
rect 241514 685992 241520 686004
rect 241572 685992 241578 686044
rect 413462 685992 413468 686044
rect 413520 686032 413526 686044
rect 430574 686032 430580 686044
rect 413520 686004 430580 686032
rect 413520 685992 413526 686004
rect 430574 685992 430580 686004
rect 430632 685992 430638 686044
rect 440510 685992 440516 686044
rect 440568 686032 440574 686044
rect 457254 686032 457260 686044
rect 440568 686004 457260 686032
rect 440568 685992 440574 686004
rect 457254 685992 457260 686004
rect 457312 685992 457318 686044
rect 468570 685992 468576 686044
rect 468628 686032 468634 686044
rect 484394 686032 484400 686044
rect 468628 686004 484400 686032
rect 468628 685992 468634 686004
rect 484394 685992 484400 686004
rect 484452 685992 484458 686044
rect 494514 685992 494520 686044
rect 494572 686032 494578 686044
rect 511350 686032 511356 686044
rect 494572 686004 511356 686032
rect 494572 685992 494578 686004
rect 511350 685992 511356 686004
rect 511408 685992 511414 686044
rect 36722 685924 36728 685976
rect 36780 685964 36786 685976
rect 62114 685964 62120 685976
rect 36780 685936 62120 685964
rect 36780 685924 36786 685936
rect 62114 685924 62120 685936
rect 62172 685924 62178 685976
rect 64138 685924 64144 685976
rect 64196 685964 64202 685976
rect 89070 685964 89076 685976
rect 64196 685936 89076 685964
rect 64196 685924 64202 685936
rect 89070 685924 89076 685936
rect 89128 685924 89134 685976
rect 90450 685924 90456 685976
rect 90508 685964 90514 685976
rect 115934 685964 115940 685976
rect 90508 685936 115940 685964
rect 90508 685924 90514 685936
rect 115934 685924 115940 685936
rect 115992 685924 115998 685976
rect 116578 685924 116584 685976
rect 116636 685964 116642 685976
rect 142982 685964 142988 685976
rect 116636 685936 142988 685964
rect 116636 685924 116642 685936
rect 142982 685924 142988 685936
rect 143040 685924 143046 685976
rect 144178 685924 144184 685976
rect 144236 685964 144242 685976
rect 170030 685964 170036 685976
rect 144236 685936 170036 685964
rect 144236 685924 144242 685936
rect 170030 685924 170036 685936
rect 170088 685924 170094 685976
rect 178402 685924 178408 685976
rect 178460 685964 178466 685976
rect 200758 685964 200764 685976
rect 178460 685936 200764 685964
rect 178460 685924 178466 685936
rect 200758 685924 200764 685936
rect 200816 685924 200822 685976
rect 251450 685924 251456 685976
rect 251508 685964 251514 685976
rect 268286 685964 268292 685976
rect 251508 685936 268292 685964
rect 251508 685924 251514 685936
rect 268286 685924 268292 685936
rect 268344 685924 268350 685976
rect 279418 685924 279424 685976
rect 279476 685964 279482 685976
rect 295794 685964 295800 685976
rect 279476 685936 295800 685964
rect 279476 685924 279482 685936
rect 295794 685924 295800 685936
rect 295852 685924 295858 685976
rect 305546 685924 305552 685976
rect 305604 685964 305610 685976
rect 322382 685964 322388 685976
rect 305604 685936 322388 685964
rect 305604 685924 305610 685936
rect 322382 685924 322388 685936
rect 322440 685924 322446 685976
rect 334618 685924 334624 685976
rect 334676 685964 334682 685976
rect 349798 685964 349804 685976
rect 334676 685936 349804 685964
rect 334676 685924 334682 685936
rect 349798 685924 349804 685936
rect 349856 685924 349862 685976
rect 359642 685924 359648 685976
rect 359700 685964 359706 685976
rect 376294 685964 376300 685976
rect 359700 685936 376300 685964
rect 359700 685924 359706 685936
rect 376294 685924 376300 685936
rect 376352 685924 376358 685976
rect 386506 685924 386512 685976
rect 386564 685964 386570 685976
rect 403342 685964 403348 685976
rect 386564 685936 403348 685964
rect 386564 685924 386570 685936
rect 403342 685924 403348 685936
rect 403400 685924 403406 685976
rect 421282 685924 421288 685976
rect 421340 685964 421346 685976
rect 443638 685964 443644 685976
rect 421340 685936 443644 685964
rect 421340 685924 421346 685936
rect 443638 685924 443644 685936
rect 443696 685924 443702 685976
rect 475378 685924 475384 685976
rect 475436 685964 475442 685976
rect 494698 685964 494704 685976
rect 475436 685936 494704 685964
rect 475436 685924 475442 685936
rect 494698 685924 494704 685936
rect 494756 685924 494762 685976
rect 522390 685924 522396 685976
rect 522448 685964 522454 685976
rect 538398 685964 538404 685976
rect 522448 685936 538404 685964
rect 522448 685924 522454 685936
rect 538398 685924 538404 685936
rect 538456 685924 538462 685976
rect 43346 685856 43352 685908
rect 43404 685896 43410 685908
rect 62758 685896 62764 685908
rect 43404 685868 62764 685896
rect 43404 685856 43410 685868
rect 62758 685856 62764 685868
rect 62816 685856 62822 685908
rect 171778 685856 171784 685908
rect 171836 685896 171842 685908
rect 197446 685896 197452 685908
rect 171836 685868 197452 685896
rect 171836 685856 171842 685868
rect 197446 685856 197452 685868
rect 197504 685856 197510 685908
rect 199378 685856 199384 685908
rect 199436 685896 199442 685908
rect 223942 685896 223948 685908
rect 199436 685868 223948 685896
rect 199436 685856 199442 685868
rect 223942 685856 223948 685868
rect 224000 685856 224006 685908
rect 225598 685856 225604 685908
rect 225656 685896 225662 685908
rect 251174 685896 251180 685908
rect 225656 685868 251180 685896
rect 225656 685856 225662 685868
rect 251174 685856 251180 685868
rect 251232 685856 251238 685908
rect 253198 685856 253204 685908
rect 253256 685896 253262 685908
rect 278038 685896 278044 685908
rect 253256 685868 278044 685896
rect 253256 685856 253262 685868
rect 278038 685856 278044 685868
rect 278096 685856 278102 685908
rect 279510 685856 279516 685908
rect 279568 685896 279574 685908
rect 305454 685896 305460 685908
rect 279568 685868 305460 685896
rect 279568 685856 279574 685868
rect 305454 685856 305460 685868
rect 305512 685856 305518 685908
rect 307018 685856 307024 685908
rect 307076 685896 307082 685908
rect 331950 685896 331956 685908
rect 307076 685868 331956 685896
rect 307076 685856 307082 685868
rect 331950 685856 331956 685868
rect 332008 685856 332014 685908
rect 333238 685856 333244 685908
rect 333296 685896 333302 685908
rect 359458 685896 359464 685908
rect 333296 685868 359464 685896
rect 333296 685856 333302 685868
rect 359458 685856 359464 685868
rect 359516 685856 359522 685908
rect 359734 685856 359740 685908
rect 359792 685896 359798 685908
rect 386046 685896 386052 685908
rect 359792 685868 386052 685896
rect 359792 685856 359798 685868
rect 386046 685856 386052 685868
rect 386104 685856 386110 685908
rect 387058 685856 387064 685908
rect 387116 685896 387122 685908
rect 412910 685896 412916 685908
rect 387116 685868 412916 685896
rect 387116 685856 387122 685868
rect 412910 685856 412916 685868
rect 412968 685856 412974 685908
rect 414658 685856 414664 685908
rect 414716 685896 414722 685908
rect 440234 685896 440240 685908
rect 414716 685868 440240 685896
rect 414716 685856 414722 685868
rect 440234 685856 440240 685868
rect 440292 685856 440298 685908
rect 442258 685856 442264 685908
rect 442316 685896 442322 685908
rect 467006 685896 467012 685908
rect 442316 685868 467012 685896
rect 442316 685856 442322 685868
rect 467006 685856 467012 685868
rect 467064 685856 467070 685908
rect 468478 685856 468484 685908
rect 468536 685896 468542 685908
rect 494054 685896 494060 685908
rect 468536 685868 494060 685896
rect 468536 685856 468542 685868
rect 494054 685856 494060 685868
rect 494112 685856 494118 685908
rect 496078 685856 496084 685908
rect 496136 685896 496142 685908
rect 520918 685896 520924 685908
rect 496136 685868 520924 685896
rect 496136 685856 496142 685868
rect 520918 685856 520924 685868
rect 520976 685856 520982 685908
rect 522298 685856 522304 685908
rect 522356 685896 522362 685908
rect 548058 685896 548064 685908
rect 522356 685868 548064 685896
rect 522356 685856 522362 685868
rect 548058 685856 548064 685868
rect 548116 685856 548122 685908
rect 285766 683272 285772 683324
rect 285824 683312 285830 683324
rect 286134 683312 286140 683324
rect 285824 683284 286140 683312
rect 285824 683272 285830 683284
rect 286134 683272 286140 683284
rect 286192 683272 286198 683324
rect 339586 683272 339592 683324
rect 339644 683312 339650 683324
rect 340138 683312 340144 683324
rect 339644 683284 340144 683312
rect 339644 683272 339650 683284
rect 340138 683272 340144 683284
rect 340196 683272 340202 683324
rect 68922 683204 68928 683256
rect 68980 683244 68986 683256
rect 118694 683244 118700 683256
rect 68980 683216 118700 683244
rect 68980 683204 68986 683216
rect 118694 683204 118700 683216
rect 118752 683204 118758 683256
rect 122742 683204 122748 683256
rect 122800 683244 122806 683256
rect 172514 683244 172520 683256
rect 122800 683216 172520 683244
rect 122800 683204 122806 683216
rect 172514 683204 172520 683216
rect 172572 683204 172578 683256
rect 230382 683204 230388 683256
rect 230440 683244 230446 683256
rect 280154 683244 280160 683256
rect 230440 683216 280160 683244
rect 230440 683204 230446 683216
rect 280154 683204 280160 683216
rect 280212 683204 280218 683256
rect 311802 683204 311808 683256
rect 311860 683244 311866 683256
rect 361574 683244 361580 683256
rect 311860 683216 361580 683244
rect 311860 683204 311866 683216
rect 361574 683204 361580 683216
rect 361632 683204 361638 683256
rect 500862 683204 500868 683256
rect 500920 683244 500926 683256
rect 550634 683244 550640 683256
rect 500920 683216 550640 683244
rect 500920 683204 500926 683216
rect 550634 683204 550640 683216
rect 550692 683204 550698 683256
rect 41322 683136 41328 683188
rect 41380 683176 41386 683188
rect 91094 683176 91100 683188
rect 41380 683148 91100 683176
rect 41380 683136 41386 683148
rect 91094 683136 91100 683148
rect 91152 683136 91158 683188
rect 148962 683136 148968 683188
rect 149020 683176 149026 683188
rect 200114 683176 200120 683188
rect 149020 683148 200120 683176
rect 149020 683136 149026 683148
rect 200114 683136 200120 683148
rect 200172 683136 200178 683188
rect 202782 683136 202788 683188
rect 202840 683176 202846 683188
rect 253934 683176 253940 683188
rect 202840 683148 253940 683176
rect 202840 683136 202846 683148
rect 253934 683136 253940 683148
rect 253992 683136 253998 683188
rect 284202 683136 284208 683188
rect 284260 683176 284266 683188
rect 335354 683176 335360 683188
rect 284260 683148 335360 683176
rect 284260 683136 284266 683148
rect 335354 683136 335360 683148
rect 335412 683136 335418 683188
rect 365622 683136 365628 683188
rect 365680 683176 365686 683188
rect 415394 683176 415400 683188
rect 365680 683148 415400 683176
rect 365680 683136 365686 683148
rect 415394 683136 415400 683148
rect 415452 683136 415458 683188
rect 419442 683136 419448 683188
rect 419500 683176 419506 683188
rect 469214 683176 469220 683188
rect 419500 683148 469220 683176
rect 419500 683136 419506 683148
rect 469214 683136 469220 683148
rect 469272 683136 469278 683188
rect 473262 683136 473268 683188
rect 473320 683176 473326 683188
rect 523034 683176 523040 683188
rect 473320 683148 523040 683176
rect 473320 683136 473326 683148
rect 523034 683136 523040 683148
rect 523092 683136 523098 683188
rect 143626 666136 143632 666188
rect 143684 666176 143690 666188
rect 144270 666176 144276 666188
rect 143684 666148 144276 666176
rect 143684 666136 143690 666148
rect 144270 666136 144276 666148
rect 144328 666136 144334 666188
rect 13722 665116 13728 665168
rect 13780 665156 13786 665168
rect 64874 665156 64880 665168
rect 13780 665128 64880 665156
rect 13780 665116 13786 665128
rect 64874 665116 64880 665128
rect 64932 665116 64938 665168
rect 95142 665116 95148 665168
rect 95200 665156 95206 665168
rect 146294 665156 146300 665168
rect 95200 665128 146300 665156
rect 95200 665116 95206 665128
rect 146294 665116 146300 665128
rect 146352 665116 146358 665168
rect 176562 665116 176568 665168
rect 176620 665156 176626 665168
rect 226334 665156 226340 665168
rect 176620 665128 226340 665156
rect 176620 665116 176626 665128
rect 226334 665116 226340 665128
rect 226392 665116 226398 665168
rect 256602 665116 256608 665168
rect 256660 665156 256666 665168
rect 307754 665156 307760 665168
rect 256660 665128 307760 665156
rect 256660 665116 256666 665128
rect 307754 665116 307760 665128
rect 307812 665116 307818 665168
rect 332502 665116 332508 665168
rect 332560 665156 332566 665168
rect 334618 665156 334624 665168
rect 332560 665128 334624 665156
rect 332560 665116 332566 665128
rect 334618 665116 334624 665128
rect 334676 665116 334682 665168
rect 338022 665116 338028 665168
rect 338080 665156 338086 665168
rect 389174 665156 389180 665168
rect 338080 665128 389180 665156
rect 338080 665116 338086 665128
rect 389174 665116 389180 665128
rect 389232 665116 389238 665168
rect 391842 665116 391848 665168
rect 391900 665156 391906 665168
rect 442994 665156 443000 665168
rect 391900 665128 443000 665156
rect 391900 665116 391906 665128
rect 442994 665116 443000 665128
rect 443052 665116 443058 665168
rect 445662 665116 445668 665168
rect 445720 665156 445726 665168
rect 496814 665156 496820 665168
rect 445720 665128 496820 665156
rect 445720 665116 445726 665128
rect 496814 665116 496820 665128
rect 496872 665116 496878 665168
rect 35618 665048 35624 665100
rect 35676 665088 35682 665100
rect 36630 665088 36636 665100
rect 35676 665060 36636 665088
rect 35676 665048 35682 665060
rect 36630 665048 36636 665060
rect 36688 665048 36694 665100
rect 467650 665048 467656 665100
rect 467708 665088 467714 665100
rect 468570 665088 468576 665100
rect 467708 665060 468576 665088
rect 467708 665048 467714 665060
rect 468570 665048 468576 665060
rect 468628 665048 468634 665100
rect 521378 663688 521384 663740
rect 521436 663728 521442 663740
rect 522390 663728 522396 663740
rect 521436 663700 522396 663728
rect 521436 663688 521442 663700
rect 522390 663688 522396 663700
rect 522448 663688 522454 663740
rect 62758 662328 62764 662380
rect 62816 662368 62822 662380
rect 70026 662368 70032 662380
rect 62816 662340 70032 662368
rect 62816 662328 62822 662340
rect 70026 662328 70032 662340
rect 70084 662328 70090 662380
rect 96706 662328 96712 662380
rect 96764 662368 96770 662380
rect 124030 662368 124036 662380
rect 96764 662340 124036 662368
rect 96764 662328 96770 662340
rect 124030 662328 124036 662340
rect 124088 662328 124094 662380
rect 150526 662328 150532 662380
rect 150584 662368 150590 662380
rect 178034 662368 178040 662380
rect 150584 662340 178040 662368
rect 150584 662328 150590 662340
rect 178034 662328 178040 662340
rect 178092 662328 178098 662380
rect 187694 662328 187700 662380
rect 187752 662368 187758 662380
rect 199378 662368 199384 662380
rect 187752 662340 199384 662368
rect 187752 662328 187758 662340
rect 199378 662328 199384 662340
rect 199436 662328 199442 662380
rect 200758 662328 200764 662380
rect 200816 662368 200822 662380
rect 204990 662368 204996 662380
rect 200816 662340 204996 662368
rect 200816 662328 200822 662340
rect 204990 662328 204996 662340
rect 205048 662328 205054 662380
rect 232038 662368 232044 662380
rect 209746 662340 232044 662368
rect 25682 662260 25688 662312
rect 25740 662300 25746 662312
rect 36722 662300 36728 662312
rect 25740 662272 36728 662300
rect 25740 662260 25746 662272
rect 36722 662260 36728 662272
rect 36780 662260 36786 662312
rect 53098 662260 53104 662312
rect 53156 662300 53162 662312
rect 64138 662300 64144 662312
rect 53156 662272 64144 662300
rect 53156 662260 53162 662272
rect 64138 662260 64144 662272
rect 64196 662260 64202 662312
rect 79686 662260 79692 662312
rect 79744 662300 79750 662312
rect 90450 662300 90456 662312
rect 79744 662272 90456 662300
rect 79744 662260 79750 662272
rect 90450 662260 90456 662272
rect 90508 662260 90514 662312
rect 106642 662260 106648 662312
rect 106700 662300 106706 662312
rect 116578 662300 116584 662312
rect 106700 662272 116584 662300
rect 106700 662260 106706 662272
rect 116578 662260 116584 662272
rect 116636 662260 116642 662312
rect 133690 662260 133696 662312
rect 133748 662300 133754 662312
rect 144178 662300 144184 662312
rect 133748 662272 144184 662300
rect 133748 662260 133754 662272
rect 144178 662260 144184 662272
rect 144236 662260 144242 662312
rect 160646 662260 160652 662312
rect 160704 662300 160710 662312
rect 171778 662300 171784 662312
rect 160704 662272 171784 662300
rect 160704 662260 160710 662272
rect 171778 662260 171784 662272
rect 171836 662260 171842 662312
rect 204346 662260 204352 662312
rect 204404 662300 204410 662312
rect 209746 662300 209774 662340
rect 232038 662328 232044 662340
rect 232096 662328 232102 662380
rect 251818 662328 251824 662380
rect 251876 662368 251882 662380
rect 258994 662368 259000 662380
rect 251876 662340 259000 662368
rect 251876 662328 251882 662340
rect 258994 662328 259000 662340
rect 259052 662328 259058 662380
rect 285766 662328 285772 662380
rect 285824 662368 285830 662380
rect 312998 662368 313004 662380
rect 285824 662340 313004 662368
rect 285824 662328 285830 662340
rect 312998 662328 313004 662340
rect 313056 662328 313062 662380
rect 339586 662328 339592 662380
rect 339644 662368 339650 662380
rect 366726 662368 366732 662380
rect 339644 662340 366732 662368
rect 339644 662328 339650 662340
rect 366726 662328 366732 662340
rect 366784 662328 366790 662380
rect 393590 662368 393596 662380
rect 373966 662340 393596 662368
rect 204404 662272 209774 662300
rect 204404 662260 204410 662272
rect 214650 662260 214656 662312
rect 214708 662300 214714 662312
rect 225598 662300 225604 662312
rect 214708 662272 225604 662300
rect 214708 662260 214714 662272
rect 225598 662260 225604 662272
rect 225656 662260 225662 662312
rect 241698 662260 241704 662312
rect 241756 662300 241762 662312
rect 253198 662300 253204 662312
rect 241756 662272 253204 662300
rect 241756 662260 241762 662272
rect 253198 662260 253204 662272
rect 253256 662260 253262 662312
rect 268654 662260 268660 662312
rect 268712 662300 268718 662312
rect 279510 662300 279516 662312
rect 268712 662272 279516 662300
rect 268712 662260 268718 662272
rect 279510 662260 279516 662272
rect 279568 662260 279574 662312
rect 295702 662260 295708 662312
rect 295760 662300 295766 662312
rect 307018 662300 307024 662312
rect 295760 662272 307024 662300
rect 295760 662260 295766 662272
rect 307018 662260 307024 662272
rect 307076 662260 307082 662312
rect 322658 662260 322664 662312
rect 322716 662300 322722 662312
rect 333238 662300 333244 662312
rect 322716 662272 333244 662300
rect 322716 662260 322722 662272
rect 333238 662260 333244 662272
rect 333296 662260 333302 662312
rect 349706 662260 349712 662312
rect 349764 662300 349770 662312
rect 359550 662300 359556 662312
rect 349764 662272 359556 662300
rect 349764 662260 349770 662272
rect 359550 662260 359556 662272
rect 359608 662260 359614 662312
rect 365806 662260 365812 662312
rect 365864 662300 365870 662312
rect 373966 662300 373994 662340
rect 393590 662328 393596 662340
rect 393648 662328 393654 662380
rect 421006 662368 421012 662380
rect 402946 662340 421012 662368
rect 365864 662272 373994 662300
rect 365864 662260 365870 662272
rect 376662 662260 376668 662312
rect 376720 662300 376726 662312
rect 387058 662300 387064 662312
rect 376720 662272 387064 662300
rect 376720 662260 376726 662272
rect 387058 662260 387064 662272
rect 387116 662260 387122 662312
rect 393406 662260 393412 662312
rect 393464 662300 393470 662312
rect 402946 662300 402974 662340
rect 421006 662328 421012 662340
rect 421064 662328 421070 662380
rect 430666 662328 430672 662380
rect 430724 662368 430730 662380
rect 442258 662368 442264 662380
rect 430724 662340 442264 662368
rect 430724 662328 430730 662340
rect 442258 662328 442264 662340
rect 442316 662328 442322 662380
rect 443638 662328 443644 662380
rect 443696 662368 443702 662380
rect 447686 662368 447692 662380
rect 443696 662340 447692 662368
rect 443696 662328 443702 662340
rect 447686 662328 447692 662340
rect 447744 662328 447750 662380
rect 494698 662328 494704 662380
rect 494756 662368 494762 662380
rect 501966 662368 501972 662380
rect 494756 662340 501972 662368
rect 494756 662328 494762 662340
rect 501966 662328 501972 662340
rect 502024 662328 502030 662380
rect 393464 662272 402974 662300
rect 393464 662260 393470 662272
rect 403710 662260 403716 662312
rect 403768 662300 403774 662312
rect 414658 662300 414664 662312
rect 403768 662272 414664 662300
rect 403768 662260 403774 662272
rect 414658 662260 414664 662272
rect 414716 662260 414722 662312
rect 457714 662260 457720 662312
rect 457772 662300 457778 662312
rect 468478 662300 468484 662312
rect 457772 662272 468484 662300
rect 457772 662260 457778 662272
rect 468478 662260 468484 662272
rect 468536 662260 468542 662312
rect 484670 662260 484676 662312
rect 484728 662300 484734 662312
rect 496078 662300 496084 662312
rect 484728 662272 496084 662300
rect 484728 662260 484734 662272
rect 496078 662260 496084 662272
rect 496136 662260 496142 662312
rect 511718 662260 511724 662312
rect 511776 662300 511782 662312
rect 522298 662300 522304 662312
rect 511776 662272 522304 662300
rect 511776 662260 511782 662272
rect 522298 662260 522304 662272
rect 522356 662260 522362 662312
rect 15194 662192 15200 662244
rect 15252 662232 15258 662244
rect 42978 662232 42984 662244
rect 15252 662204 42984 662232
rect 15252 662192 15258 662204
rect 42978 662192 42984 662204
rect 43036 662192 43042 662244
rect 69106 662192 69112 662244
rect 69164 662232 69170 662244
rect 96982 662232 96988 662244
rect 69164 662204 96988 662232
rect 69164 662192 69170 662204
rect 96982 662192 96988 662204
rect 97040 662192 97046 662244
rect 122926 662192 122932 662244
rect 122984 662232 122990 662244
rect 150986 662232 150992 662244
rect 122984 662204 150992 662232
rect 122984 662192 122990 662204
rect 150986 662192 150992 662204
rect 151044 662192 151050 662244
rect 258166 662192 258172 662244
rect 258224 662232 258230 662244
rect 286042 662232 286048 662244
rect 258224 662204 286048 662232
rect 258224 662192 258230 662204
rect 286042 662192 286048 662204
rect 286100 662192 286106 662244
rect 311986 662192 311992 662244
rect 312044 662232 312050 662244
rect 340046 662232 340052 662244
rect 312044 662204 340052 662232
rect 312044 662192 312050 662204
rect 340046 662192 340052 662204
rect 340104 662192 340110 662244
rect 447226 662192 447232 662244
rect 447284 662232 447290 662244
rect 475010 662232 475016 662244
rect 447284 662204 475016 662232
rect 447284 662192 447290 662204
rect 475010 662192 475016 662204
rect 475068 662192 475074 662244
rect 501046 662192 501052 662244
rect 501104 662232 501110 662244
rect 529014 662232 529020 662244
rect 501104 662204 529020 662232
rect 501104 662192 501110 662204
rect 529014 662192 529020 662204
rect 529072 662192 529078 662244
rect 16022 658928 16028 658980
rect 16080 658968 16086 658980
rect 529014 658968 529020 658980
rect 16080 658940 529020 658968
rect 16080 658928 16086 658940
rect 529014 658928 529020 658940
rect 529072 658928 529078 658980
rect 25682 658520 25688 658572
rect 25740 658560 25746 658572
rect 146938 658560 146944 658572
rect 25740 658532 146944 658560
rect 25740 658520 25746 658532
rect 146938 658520 146944 658532
rect 146996 658520 147002 658572
rect 36722 658452 36728 658504
rect 36780 658492 36786 658504
rect 52638 658492 52644 658504
rect 36780 658464 52644 658492
rect 36780 658452 36786 658464
rect 52638 658452 52644 658464
rect 52696 658452 52702 658504
rect 232038 658452 232044 658504
rect 232096 658492 232102 658504
rect 251818 658492 251824 658504
rect 232096 658464 251824 658492
rect 232096 658452 232102 658464
rect 251818 658452 251824 658464
rect 251876 658452 251882 658504
rect 475010 658452 475016 658504
rect 475068 658492 475074 658504
rect 494698 658492 494704 658504
rect 475068 658464 494704 658492
rect 475068 658452 475074 658464
rect 494698 658452 494704 658464
rect 494756 658452 494762 658504
rect 62482 658384 62488 658436
rect 62540 658424 62546 658436
rect 79686 658424 79692 658436
rect 62540 658396 79692 658424
rect 62540 658384 62546 658396
rect 79686 658384 79692 658396
rect 79744 658384 79750 658436
rect 90450 658384 90456 658436
rect 90508 658424 90514 658436
rect 106642 658424 106648 658436
rect 90508 658396 106648 658424
rect 90508 658384 90514 658396
rect 106642 658384 106648 658396
rect 106700 658384 106706 658436
rect 116486 658384 116492 658436
rect 116544 658424 116550 658436
rect 133690 658424 133696 658436
rect 116544 658396 133696 658424
rect 116544 658384 116550 658396
rect 133690 658384 133696 658396
rect 133748 658384 133754 658436
rect 170490 658384 170496 658436
rect 170548 658424 170554 658436
rect 187694 658424 187700 658436
rect 170548 658396 187700 658424
rect 170548 658384 170554 658396
rect 187694 658384 187700 658396
rect 187752 658384 187758 658436
rect 197446 658384 197452 658436
rect 197504 658424 197510 658436
rect 214650 658424 214656 658436
rect 197504 658396 214656 658424
rect 197504 658384 197510 658396
rect 214650 658384 214656 658396
rect 214708 658384 214714 658436
rect 224494 658384 224500 658436
rect 224552 658424 224558 658436
rect 241698 658424 241704 658436
rect 224552 658396 241704 658424
rect 224552 658384 224558 658396
rect 241698 658384 241704 658396
rect 241756 658384 241762 658436
rect 413462 658384 413468 658436
rect 413520 658424 413526 658436
rect 430666 658424 430672 658436
rect 413520 658396 430672 658424
rect 413520 658384 413526 658396
rect 430666 658384 430672 658396
rect 430724 658384 430730 658436
rect 440510 658384 440516 658436
rect 440568 658424 440574 658436
rect 457622 658424 457628 658436
rect 440568 658396 457628 658424
rect 440568 658384 440574 658396
rect 457622 658384 457628 658396
rect 457680 658384 457686 658436
rect 468478 658384 468484 658436
rect 468536 658424 468542 658436
rect 484670 658424 484676 658436
rect 468536 658396 484676 658424
rect 468536 658384 468542 658396
rect 484670 658384 484676 658396
rect 484728 658384 484734 658436
rect 36814 658316 36820 658368
rect 36872 658356 36878 658368
rect 62298 658356 62304 658368
rect 36872 658328 62304 658356
rect 36872 658316 36878 658328
rect 62298 658316 62304 658328
rect 62356 658316 62362 658368
rect 64138 658316 64144 658368
rect 64196 658356 64202 658368
rect 89346 658356 89352 658368
rect 64196 658328 89352 658356
rect 64196 658316 64202 658328
rect 89346 658316 89352 658328
rect 89404 658316 89410 658368
rect 90358 658316 90364 658368
rect 90416 658356 90422 658368
rect 116302 658356 116308 658368
rect 90416 658328 116308 658356
rect 90416 658316 90422 658328
rect 116302 658316 116308 658328
rect 116360 658316 116366 658368
rect 116578 658316 116584 658368
rect 116636 658356 116642 658368
rect 143350 658356 143356 658368
rect 116636 658328 143356 658356
rect 116636 658316 116642 658328
rect 143350 658316 143356 658328
rect 143408 658316 143414 658368
rect 144270 658316 144276 658368
rect 144328 658356 144334 658368
rect 170306 658356 170312 658368
rect 144328 658328 170312 658356
rect 144328 658316 144334 658328
rect 170306 658316 170312 658328
rect 170364 658316 170370 658368
rect 178034 658316 178040 658368
rect 178092 658356 178098 658368
rect 200758 658356 200764 658368
rect 178092 658328 200764 658356
rect 178092 658316 178098 658328
rect 200758 658316 200764 658328
rect 200816 658316 200822 658368
rect 251450 658316 251456 658368
rect 251508 658356 251514 658368
rect 268654 658356 268660 658368
rect 251508 658328 268660 658356
rect 251508 658316 251514 658328
rect 268654 658316 268660 658328
rect 268712 658316 268718 658368
rect 279418 658316 279424 658368
rect 279476 658356 279482 658368
rect 295702 658356 295708 658368
rect 279476 658328 295708 658356
rect 279476 658316 279482 658328
rect 295702 658316 295708 658328
rect 295760 658316 295766 658368
rect 305454 658316 305460 658368
rect 305512 658356 305518 658368
rect 322658 658356 322664 658368
rect 305512 658328 322664 658356
rect 305512 658316 305518 658328
rect 322658 658316 322664 658328
rect 322716 658316 322722 658368
rect 335998 658316 336004 658368
rect 336056 658356 336062 658368
rect 349706 658356 349712 658368
rect 336056 658328 349712 658356
rect 336056 658316 336062 658328
rect 349706 658316 349712 658328
rect 349764 658316 349770 658368
rect 359458 658316 359464 658368
rect 359516 658356 359522 658368
rect 376662 658356 376668 658368
rect 359516 658328 376668 658356
rect 359516 658316 359522 658328
rect 376662 658316 376668 658328
rect 376720 658316 376726 658368
rect 386506 658316 386512 658368
rect 386564 658356 386570 658368
rect 403618 658356 403624 658368
rect 386564 658328 403624 658356
rect 386564 658316 386570 658328
rect 403618 658316 403624 658328
rect 403676 658316 403682 658368
rect 421006 658316 421012 658368
rect 421064 658356 421070 658368
rect 446398 658356 446404 658368
rect 421064 658328 446404 658356
rect 421064 658316 421070 658328
rect 446398 658316 446404 658328
rect 446456 658316 446462 658368
rect 494514 658316 494520 658368
rect 494572 658356 494578 658368
rect 511626 658356 511632 658368
rect 494572 658328 511632 658356
rect 494572 658316 494578 658328
rect 511626 658316 511632 658328
rect 511684 658316 511690 658368
rect 522298 658316 522304 658368
rect 522356 658356 522362 658368
rect 538674 658356 538680 658368
rect 522356 658328 538680 658356
rect 522356 658316 522362 658328
rect 538674 658316 538680 658328
rect 538732 658316 538738 658368
rect 43070 658248 43076 658300
rect 43128 658288 43134 658300
rect 62758 658288 62764 658300
rect 43128 658260 62764 658288
rect 43128 658248 43134 658260
rect 62758 658248 62764 658260
rect 62816 658248 62822 658300
rect 144178 658248 144184 658300
rect 144236 658288 144242 658300
rect 160646 658288 160652 658300
rect 144236 658260 160652 658288
rect 144236 658248 144242 658260
rect 160646 658248 160652 658260
rect 160704 658248 160710 658300
rect 171778 658248 171784 658300
rect 171836 658288 171842 658300
rect 197354 658288 197360 658300
rect 171836 658260 197360 658288
rect 171836 658248 171842 658260
rect 197354 658248 197360 658260
rect 197412 658248 197418 658300
rect 199378 658248 199384 658300
rect 199436 658288 199442 658300
rect 224310 658288 224316 658300
rect 199436 658260 224316 658288
rect 199436 658248 199442 658260
rect 224310 658248 224316 658260
rect 224368 658248 224374 658300
rect 225598 658248 225604 658300
rect 225656 658288 225662 658300
rect 251358 658288 251364 658300
rect 225656 658260 251364 658288
rect 225656 658248 225662 658260
rect 251358 658248 251364 658260
rect 251416 658248 251422 658300
rect 253198 658248 253204 658300
rect 253256 658288 253262 658300
rect 278314 658288 278320 658300
rect 253256 658260 278320 658288
rect 253256 658248 253262 658260
rect 278314 658248 278320 658260
rect 278372 658248 278378 658300
rect 279510 658248 279516 658300
rect 279568 658288 279574 658300
rect 305362 658288 305368 658300
rect 279568 658260 305368 658288
rect 279568 658248 279574 658260
rect 305362 658248 305368 658260
rect 305420 658248 305426 658300
rect 307018 658248 307024 658300
rect 307076 658288 307082 658300
rect 332318 658288 332324 658300
rect 307076 658260 332324 658288
rect 307076 658248 307082 658260
rect 332318 658248 332324 658260
rect 332376 658248 332382 658300
rect 333238 658248 333244 658300
rect 333296 658288 333302 658300
rect 359366 658288 359372 658300
rect 333296 658260 359372 658288
rect 333296 658248 333302 658260
rect 359366 658248 359372 658260
rect 359424 658248 359430 658300
rect 359550 658248 359556 658300
rect 359608 658288 359614 658300
rect 386322 658288 386328 658300
rect 359608 658260 386328 658288
rect 359608 658248 359614 658260
rect 386322 658248 386328 658260
rect 386380 658248 386386 658300
rect 387058 658248 387064 658300
rect 387116 658288 387122 658300
rect 413278 658288 413284 658300
rect 387116 658260 413284 658288
rect 387116 658248 387122 658260
rect 413278 658248 413284 658260
rect 413336 658248 413342 658300
rect 414658 658248 414664 658300
rect 414716 658288 414722 658300
rect 440326 658288 440332 658300
rect 414716 658260 440332 658288
rect 414716 658248 414722 658260
rect 440326 658248 440332 658260
rect 440384 658248 440390 658300
rect 442258 658248 442264 658300
rect 442316 658288 442322 658300
rect 467282 658288 467288 658300
rect 442316 658260 467288 658288
rect 442316 658248 442322 658260
rect 467282 658248 467288 658260
rect 467340 658248 467346 658300
rect 468570 658248 468576 658300
rect 468628 658288 468634 658300
rect 494330 658288 494336 658300
rect 468628 658260 494336 658288
rect 468628 658248 468634 658260
rect 494330 658248 494336 658260
rect 494388 658248 494394 658300
rect 496078 658248 496084 658300
rect 496136 658288 496142 658300
rect 521286 658288 521292 658300
rect 496136 658260 521292 658288
rect 496136 658248 496142 658260
rect 521286 658248 521292 658260
rect 521344 658248 521350 658300
rect 522390 658248 522396 658300
rect 522448 658288 522454 658300
rect 548334 658288 548340 658300
rect 522448 658260 548340 658288
rect 522448 658248 522454 658260
rect 548334 658248 548340 658260
rect 548392 658248 548398 658300
rect 37918 657500 37924 657552
rect 37976 657540 37982 657552
rect 526438 657540 526444 657552
rect 37976 657512 526444 657540
rect 37976 657500 37982 657512
rect 526438 657500 526444 657512
rect 526496 657500 526502 657552
rect 35618 656888 35624 656940
rect 35676 656928 35682 656940
rect 36630 656928 36636 656940
rect 35676 656900 36636 656928
rect 35676 656888 35682 656900
rect 36630 656888 36636 656900
rect 36688 656888 36694 656940
rect 68922 655664 68928 655716
rect 68980 655704 68986 655716
rect 118694 655704 118700 655716
rect 68980 655676 118700 655704
rect 68980 655664 68986 655676
rect 118694 655664 118700 655676
rect 118752 655664 118758 655716
rect 311802 655664 311808 655716
rect 311860 655704 311866 655716
rect 361574 655704 361580 655716
rect 311860 655676 361580 655704
rect 311860 655664 311866 655676
rect 361574 655664 361580 655676
rect 361632 655664 361638 655716
rect 41322 655596 41328 655648
rect 41380 655636 41386 655648
rect 91094 655636 91100 655648
rect 41380 655608 91100 655636
rect 41380 655596 41386 655608
rect 91094 655596 91100 655608
rect 91152 655596 91158 655648
rect 122742 655596 122748 655648
rect 122800 655636 122806 655648
rect 172514 655636 172520 655648
rect 122800 655608 172520 655636
rect 122800 655596 122806 655608
rect 172514 655596 172520 655608
rect 172572 655596 172578 655648
rect 176562 655596 176568 655648
rect 176620 655636 176626 655648
rect 226334 655636 226340 655648
rect 176620 655608 226340 655636
rect 176620 655596 176626 655608
rect 226334 655596 226340 655608
rect 226392 655596 226398 655648
rect 230382 655596 230388 655648
rect 230440 655636 230446 655648
rect 280154 655636 280160 655648
rect 230440 655608 280160 655636
rect 230440 655596 230446 655608
rect 280154 655596 280160 655608
rect 280212 655596 280218 655648
rect 284202 655596 284208 655648
rect 284260 655636 284266 655648
rect 335354 655636 335360 655648
rect 284260 655608 335360 655636
rect 284260 655596 284266 655608
rect 335354 655596 335360 655608
rect 335412 655596 335418 655648
rect 365622 655596 365628 655648
rect 365680 655636 365686 655648
rect 415394 655636 415400 655648
rect 365680 655608 415400 655636
rect 365680 655596 365686 655608
rect 415394 655596 415400 655608
rect 415452 655596 415458 655648
rect 419442 655596 419448 655648
rect 419500 655636 419506 655648
rect 469214 655636 469220 655648
rect 419500 655608 469220 655636
rect 419500 655596 419506 655608
rect 469214 655596 469220 655608
rect 469272 655596 469278 655648
rect 473262 655596 473268 655648
rect 473320 655636 473326 655648
rect 523034 655636 523040 655648
rect 473320 655608 523040 655636
rect 473320 655596 473326 655608
rect 523034 655596 523040 655608
rect 523092 655596 523098 655648
rect 13722 655528 13728 655580
rect 13780 655568 13786 655580
rect 64874 655568 64880 655580
rect 13780 655540 64880 655568
rect 13780 655528 13786 655540
rect 64874 655528 64880 655540
rect 64932 655528 64938 655580
rect 96614 655528 96620 655580
rect 96672 655568 96678 655580
rect 146294 655568 146300 655580
rect 96672 655540 146300 655568
rect 96672 655528 96678 655540
rect 146294 655528 146300 655540
rect 146352 655528 146358 655580
rect 148962 655528 148968 655580
rect 149020 655568 149026 655580
rect 200114 655568 200120 655580
rect 149020 655540 200120 655568
rect 149020 655528 149026 655540
rect 200114 655528 200120 655540
rect 200172 655528 200178 655580
rect 202782 655528 202788 655580
rect 202840 655568 202846 655580
rect 253934 655568 253940 655580
rect 202840 655540 253940 655568
rect 202840 655528 202846 655540
rect 253934 655528 253940 655540
rect 253992 655528 253998 655580
rect 256602 655528 256608 655580
rect 256660 655568 256666 655580
rect 307754 655568 307760 655580
rect 256660 655540 307760 655568
rect 256660 655528 256666 655540
rect 307754 655528 307760 655540
rect 307812 655528 307818 655580
rect 338022 655528 338028 655580
rect 338080 655568 338086 655580
rect 389174 655568 389180 655580
rect 338080 655540 389180 655568
rect 338080 655528 338086 655540
rect 389174 655528 389180 655540
rect 389232 655528 389238 655580
rect 391842 655528 391848 655580
rect 391900 655568 391906 655580
rect 442994 655568 443000 655580
rect 391900 655540 443000 655568
rect 391900 655528 391906 655540
rect 442994 655528 443000 655540
rect 443052 655528 443058 655580
rect 445662 655528 445668 655580
rect 445720 655568 445726 655580
rect 496814 655568 496820 655580
rect 445720 655540 496820 655568
rect 445720 655528 445726 655540
rect 496814 655528 496820 655540
rect 496872 655528 496878 655580
rect 500862 655528 500868 655580
rect 500920 655568 500926 655580
rect 550634 655568 550640 655580
rect 500920 655540 550640 655568
rect 500920 655528 500926 655540
rect 550634 655528 550640 655540
rect 550692 655528 550698 655580
rect 95142 654032 95148 654084
rect 95200 654072 95206 654084
rect 96614 654072 96620 654084
rect 95200 654044 96620 654072
rect 95200 654032 95206 654044
rect 96614 654032 96620 654044
rect 96672 654032 96678 654084
rect 35618 637508 35624 637560
rect 35676 637548 35682 637560
rect 36722 637548 36728 637560
rect 35676 637520 36728 637548
rect 35676 637508 35682 637520
rect 36722 637508 36728 637520
rect 36780 637508 36786 637560
rect 89714 637508 89720 637560
rect 89772 637548 89778 637560
rect 90450 637548 90456 637560
rect 89772 637520 90456 637548
rect 89772 637508 89778 637520
rect 90450 637508 90456 637520
rect 90508 637508 90514 637560
rect 332594 637508 332600 637560
rect 332652 637548 332658 637560
rect 335998 637548 336004 637560
rect 332652 637520 336004 637548
rect 332652 637508 332658 637520
rect 335998 637508 336004 637520
rect 336056 637508 336062 637560
rect 446398 637508 446404 637560
rect 446456 637548 446462 637560
rect 447686 637548 447692 637560
rect 446456 637520 447692 637548
rect 446456 637508 446462 637520
rect 447686 637508 447692 637520
rect 447744 637508 447750 637560
rect 62758 634720 62764 634772
rect 62816 634760 62822 634772
rect 69750 634760 69756 634772
rect 62816 634732 69756 634760
rect 62816 634720 62822 634732
rect 69750 634720 69756 634732
rect 69808 634720 69814 634772
rect 96706 634720 96712 634772
rect 96764 634760 96770 634772
rect 96764 634732 103514 634760
rect 96764 634720 96770 634732
rect 15194 634652 15200 634704
rect 15252 634692 15258 634704
rect 42794 634692 42800 634704
rect 15252 634664 42800 634692
rect 15252 634652 15258 634664
rect 42794 634652 42800 634664
rect 42852 634652 42858 634704
rect 53098 634652 53104 634704
rect 53156 634692 53162 634704
rect 64138 634692 64144 634704
rect 53156 634664 64144 634692
rect 53156 634652 53162 634664
rect 64138 634652 64144 634664
rect 64196 634652 64202 634704
rect 69106 634652 69112 634704
rect 69164 634692 69170 634704
rect 96798 634692 96804 634704
rect 69164 634664 96804 634692
rect 69164 634652 69170 634664
rect 96798 634652 96804 634664
rect 96856 634652 96862 634704
rect 103486 634692 103514 634732
rect 200758 634720 200764 634772
rect 200816 634760 200822 634772
rect 204622 634760 204628 634772
rect 200816 634732 204628 634760
rect 200816 634720 200822 634732
rect 204622 634720 204628 634732
rect 204680 634720 204686 634772
rect 251818 634720 251824 634772
rect 251876 634760 251882 634772
rect 258718 634760 258724 634772
rect 251876 634732 258724 634760
rect 251876 634720 251882 634732
rect 258718 634720 258724 634732
rect 258776 634720 258782 634772
rect 494698 634720 494704 634772
rect 494756 634760 494762 634772
rect 501598 634760 501604 634772
rect 494756 634732 501604 634760
rect 494756 634720 494762 634732
rect 501598 634720 501604 634732
rect 501656 634720 501662 634772
rect 521470 634720 521476 634772
rect 521528 634760 521534 634772
rect 522298 634760 522304 634772
rect 521528 634732 522304 634760
rect 521528 634720 521534 634732
rect 522298 634720 522304 634732
rect 522356 634720 522362 634772
rect 123662 634692 123668 634704
rect 103486 634664 123668 634692
rect 123662 634652 123668 634664
rect 123720 634652 123726 634704
rect 149698 634652 149704 634704
rect 149756 634692 149762 634704
rect 547966 634692 547972 634704
rect 149756 634664 547972 634692
rect 149756 634652 149762 634664
rect 547966 634652 547972 634664
rect 548024 634652 548030 634704
rect 26050 634584 26056 634636
rect 26108 634624 26114 634636
rect 36814 634624 36820 634636
rect 26108 634596 36820 634624
rect 26108 634584 26114 634596
rect 36814 634584 36820 634596
rect 36872 634584 36878 634636
rect 79962 634584 79968 634636
rect 80020 634624 80026 634636
rect 90358 634624 90364 634636
rect 80020 634596 90364 634624
rect 80020 634584 80026 634596
rect 90358 634584 90364 634596
rect 90416 634584 90422 634636
rect 106550 634584 106556 634636
rect 106608 634624 106614 634636
rect 116578 634624 116584 634636
rect 106608 634596 116584 634624
rect 106608 634584 106614 634596
rect 116578 634584 116584 634596
rect 116636 634584 116642 634636
rect 133782 634584 133788 634636
rect 133840 634624 133846 634636
rect 144270 634624 144276 634636
rect 133840 634596 144276 634624
rect 133840 634584 133846 634596
rect 144270 634584 144276 634596
rect 144328 634584 144334 634636
rect 150526 634584 150532 634636
rect 150584 634624 150590 634636
rect 178126 634624 178132 634636
rect 150584 634596 178132 634624
rect 150584 634584 150590 634596
rect 178126 634584 178132 634596
rect 178184 634584 178190 634636
rect 187970 634584 187976 634636
rect 188028 634624 188034 634636
rect 199378 634624 199384 634636
rect 188028 634596 199384 634624
rect 188028 634584 188034 634596
rect 199378 634584 199384 634596
rect 199436 634584 199442 634636
rect 204346 634584 204352 634636
rect 204404 634624 204410 634636
rect 231946 634624 231952 634636
rect 204404 634596 231952 634624
rect 204404 634584 204410 634596
rect 231946 634584 231952 634596
rect 232004 634584 232010 634636
rect 242066 634584 242072 634636
rect 242124 634624 242130 634636
rect 253198 634624 253204 634636
rect 242124 634596 253204 634624
rect 242124 634584 242130 634596
rect 253198 634584 253204 634596
rect 253256 634584 253262 634636
rect 258166 634584 258172 634636
rect 258224 634624 258230 634636
rect 258224 634596 281764 634624
rect 258224 634584 258230 634596
rect 122926 634516 122932 634568
rect 122984 634556 122990 634568
rect 150710 634556 150716 634568
rect 122984 634528 150716 634556
rect 122984 634516 122990 634528
rect 150710 634516 150716 634528
rect 150768 634516 150774 634568
rect 160554 634516 160560 634568
rect 160612 634556 160618 634568
rect 171778 634556 171784 634568
rect 160612 634528 171784 634556
rect 160612 634516 160618 634528
rect 171778 634516 171784 634528
rect 171836 634516 171842 634568
rect 215018 634516 215024 634568
rect 215076 634556 215082 634568
rect 225598 634556 225604 634568
rect 215076 634528 225604 634556
rect 215076 634516 215082 634528
rect 225598 634516 225604 634528
rect 225656 634516 225662 634568
rect 268930 634516 268936 634568
rect 268988 634556 268994 634568
rect 279510 634556 279516 634568
rect 268988 634528 279516 634556
rect 268988 634516 268994 634528
rect 279510 634516 279516 634528
rect 279568 634516 279574 634568
rect 281736 634556 281764 634596
rect 285766 634584 285772 634636
rect 285824 634624 285830 634636
rect 312630 634624 312636 634636
rect 285824 634596 312636 634624
rect 285824 634584 285830 634596
rect 312630 634584 312636 634596
rect 312688 634584 312694 634636
rect 340138 634624 340144 634636
rect 316006 634596 340144 634624
rect 286134 634556 286140 634568
rect 281736 634528 286140 634556
rect 286134 634516 286140 634528
rect 286192 634516 286198 634568
rect 295978 634516 295984 634568
rect 296036 634556 296042 634568
rect 307018 634556 307024 634568
rect 296036 634528 307024 634556
rect 296036 634516 296042 634528
rect 307018 634516 307024 634528
rect 307076 634516 307082 634568
rect 311986 634516 311992 634568
rect 312044 634556 312050 634568
rect 316006 634556 316034 634596
rect 340138 634584 340144 634596
rect 340196 634584 340202 634636
rect 366726 634624 366732 634636
rect 344986 634596 366732 634624
rect 312044 634528 316034 634556
rect 312044 634516 312050 634528
rect 322842 634516 322848 634568
rect 322900 634556 322906 634568
rect 333238 634556 333244 634568
rect 322900 634528 333244 634556
rect 322900 634516 322906 634528
rect 333238 634516 333244 634528
rect 333296 634516 333302 634568
rect 339586 634516 339592 634568
rect 339644 634556 339650 634568
rect 344986 634556 345014 634596
rect 366726 634584 366732 634596
rect 366784 634584 366790 634636
rect 393590 634624 393596 634636
rect 373966 634596 393596 634624
rect 339644 634528 345014 634556
rect 339644 634516 339650 634528
rect 350074 634516 350080 634568
rect 350132 634556 350138 634568
rect 359550 634556 359556 634568
rect 350132 634528 359556 634556
rect 350132 634516 350138 634528
rect 359550 634516 359556 634528
rect 359608 634516 359614 634568
rect 365806 634516 365812 634568
rect 365864 634556 365870 634568
rect 373966 634556 373994 634596
rect 393590 634584 393596 634596
rect 393648 634584 393654 634636
rect 420914 634624 420920 634636
rect 402946 634596 420920 634624
rect 365864 634528 373994 634556
rect 365864 634516 365870 634528
rect 376570 634516 376576 634568
rect 376628 634556 376634 634568
rect 387058 634556 387064 634568
rect 376628 634528 387064 634556
rect 376628 634516 376634 634528
rect 387058 634516 387064 634528
rect 387116 634516 387122 634568
rect 393406 634516 393412 634568
rect 393464 634556 393470 634568
rect 402946 634556 402974 634596
rect 420914 634584 420920 634596
rect 420972 634584 420978 634636
rect 431034 634584 431040 634636
rect 431092 634624 431098 634636
rect 442258 634624 442264 634636
rect 431092 634596 442264 634624
rect 431092 634584 431098 634596
rect 442258 634584 442264 634596
rect 442316 634584 442322 634636
rect 447226 634584 447232 634636
rect 447284 634624 447290 634636
rect 474734 634624 474740 634636
rect 447284 634596 474740 634624
rect 447284 634584 447290 634596
rect 474734 634584 474740 634596
rect 474792 634584 474798 634636
rect 484946 634584 484952 634636
rect 485004 634624 485010 634636
rect 496078 634624 496084 634636
rect 485004 634596 496084 634624
rect 485004 634584 485010 634596
rect 496078 634584 496084 634596
rect 496136 634584 496142 634636
rect 501046 634584 501052 634636
rect 501104 634624 501110 634636
rect 528646 634624 528652 634636
rect 501104 634596 528652 634624
rect 501104 634584 501110 634596
rect 528646 634584 528652 634596
rect 528704 634584 528710 634636
rect 393464 634528 402974 634556
rect 393464 634516 393470 634528
rect 403986 634516 403992 634568
rect 404044 634556 404050 634568
rect 414658 634556 414664 634568
rect 404044 634528 414664 634556
rect 404044 634516 404050 634528
rect 414658 634516 414664 634528
rect 414716 634516 414722 634568
rect 458082 634516 458088 634568
rect 458140 634556 458146 634568
rect 468570 634556 468576 634568
rect 458140 634528 468576 634556
rect 458140 634516 458146 634528
rect 468570 634516 468576 634528
rect 468628 634516 468634 634568
rect 511810 634516 511816 634568
rect 511868 634556 511874 634568
rect 522390 634556 522396 634568
rect 511868 634528 522396 634556
rect 511868 634516 511874 634528
rect 522390 634516 522396 634528
rect 522448 634516 522454 634568
rect 36538 634448 36544 634500
rect 36596 634488 36602 634500
rect 538398 634488 538404 634500
rect 36596 634460 538404 634488
rect 36596 634448 36602 634460
rect 538398 634448 538404 634460
rect 538456 634448 538462 634500
rect 16298 632680 16304 632732
rect 16356 632720 16362 632732
rect 528738 632720 528744 632732
rect 16356 632692 528744 632720
rect 16356 632680 16362 632692
rect 528738 632680 528744 632692
rect 528796 632680 528802 632732
rect 25958 632340 25964 632392
rect 26016 632380 26022 632392
rect 148318 632380 148324 632392
rect 26016 632352 148324 632380
rect 26016 632340 26022 632352
rect 148318 632340 148324 632352
rect 148376 632340 148382 632392
rect 36722 632272 36728 632324
rect 36780 632312 36786 632324
rect 52454 632312 52460 632324
rect 36780 632284 52460 632312
rect 36780 632272 36786 632284
rect 52454 632272 52460 632284
rect 52512 632272 52518 632324
rect 232314 632272 232320 632324
rect 232372 632312 232378 632324
rect 251818 632312 251824 632324
rect 232372 632284 251824 632312
rect 232372 632272 232378 632284
rect 251818 632272 251824 632284
rect 251876 632272 251882 632324
rect 475378 632272 475384 632324
rect 475436 632312 475442 632324
rect 494698 632312 494704 632324
rect 475436 632284 494704 632312
rect 475436 632272 475442 632284
rect 494698 632272 494704 632284
rect 494756 632272 494762 632324
rect 62482 632204 62488 632256
rect 62540 632244 62546 632256
rect 79318 632244 79324 632256
rect 62540 632216 79324 632244
rect 62540 632204 62546 632216
rect 79318 632204 79324 632216
rect 79376 632204 79382 632256
rect 90358 632204 90364 632256
rect 90416 632244 90422 632256
rect 106366 632244 106372 632256
rect 90416 632216 106372 632244
rect 90416 632204 90422 632216
rect 106366 632204 106372 632216
rect 106424 632204 106430 632256
rect 116486 632204 116492 632256
rect 116544 632244 116550 632256
rect 133414 632244 133420 632256
rect 116544 632216 133420 632244
rect 116544 632204 116550 632216
rect 133414 632204 133420 632216
rect 133472 632204 133478 632256
rect 170490 632204 170496 632256
rect 170548 632244 170554 632256
rect 187786 632244 187792 632256
rect 170548 632216 187792 632244
rect 170548 632204 170554 632216
rect 187786 632204 187792 632216
rect 187844 632204 187850 632256
rect 197538 632204 197544 632256
rect 197596 632244 197602 632256
rect 214374 632244 214380 632256
rect 197596 632216 214380 632244
rect 197596 632204 197602 632216
rect 214374 632204 214380 632216
rect 214432 632204 214438 632256
rect 224494 632204 224500 632256
rect 224552 632244 224558 632256
rect 241514 632244 241520 632256
rect 224552 632216 241520 632244
rect 224552 632204 224558 632216
rect 241514 632204 241520 632216
rect 241572 632204 241578 632256
rect 413462 632204 413468 632256
rect 413520 632244 413526 632256
rect 430574 632244 430580 632256
rect 413520 632216 430580 632244
rect 413520 632204 413526 632216
rect 430574 632204 430580 632216
rect 430632 632204 430638 632256
rect 440510 632204 440516 632256
rect 440568 632244 440574 632256
rect 457254 632244 457260 632256
rect 440568 632216 457260 632244
rect 440568 632204 440574 632216
rect 457254 632204 457260 632216
rect 457312 632204 457318 632256
rect 468570 632204 468576 632256
rect 468628 632244 468634 632256
rect 484394 632244 484400 632256
rect 468628 632216 484400 632244
rect 468628 632204 468634 632216
rect 484394 632204 484400 632216
rect 484452 632204 484458 632256
rect 36814 632136 36820 632188
rect 36872 632176 36878 632188
rect 62114 632176 62120 632188
rect 36872 632148 62120 632176
rect 36872 632136 36878 632148
rect 62114 632136 62120 632148
rect 62172 632136 62178 632188
rect 64138 632136 64144 632188
rect 64196 632176 64202 632188
rect 89070 632176 89076 632188
rect 64196 632148 89076 632176
rect 64196 632136 64202 632148
rect 89070 632136 89076 632148
rect 89128 632136 89134 632188
rect 90450 632136 90456 632188
rect 90508 632176 90514 632188
rect 115934 632176 115940 632188
rect 90508 632148 115940 632176
rect 90508 632136 90514 632148
rect 115934 632136 115940 632148
rect 115992 632136 115998 632188
rect 116578 632136 116584 632188
rect 116636 632176 116642 632188
rect 142982 632176 142988 632188
rect 116636 632148 142988 632176
rect 116636 632136 116642 632148
rect 142982 632136 142988 632148
rect 143040 632136 143046 632188
rect 144270 632136 144276 632188
rect 144328 632176 144334 632188
rect 170030 632176 170036 632188
rect 144328 632148 170036 632176
rect 144328 632136 144334 632148
rect 170030 632136 170036 632148
rect 170088 632136 170094 632188
rect 178402 632136 178408 632188
rect 178460 632176 178466 632188
rect 200758 632176 200764 632188
rect 178460 632148 200764 632176
rect 178460 632136 178466 632148
rect 200758 632136 200764 632148
rect 200816 632136 200822 632188
rect 251450 632136 251456 632188
rect 251508 632176 251514 632188
rect 268286 632176 268292 632188
rect 251508 632148 268292 632176
rect 251508 632136 251514 632148
rect 268286 632136 268292 632148
rect 268344 632136 268350 632188
rect 279418 632136 279424 632188
rect 279476 632176 279482 632188
rect 295794 632176 295800 632188
rect 279476 632148 295800 632176
rect 279476 632136 279482 632148
rect 295794 632136 295800 632148
rect 295852 632136 295858 632188
rect 305638 632136 305644 632188
rect 305696 632176 305702 632188
rect 322382 632176 322388 632188
rect 305696 632148 322388 632176
rect 305696 632136 305702 632148
rect 322382 632136 322388 632148
rect 322440 632136 322446 632188
rect 335998 632136 336004 632188
rect 336056 632176 336062 632188
rect 349798 632176 349804 632188
rect 336056 632148 349804 632176
rect 336056 632136 336062 632148
rect 349798 632136 349804 632148
rect 349856 632136 349862 632188
rect 359550 632136 359556 632188
rect 359608 632176 359614 632188
rect 376294 632176 376300 632188
rect 359608 632148 376300 632176
rect 359608 632136 359614 632148
rect 376294 632136 376300 632148
rect 376352 632136 376358 632188
rect 386506 632136 386512 632188
rect 386564 632176 386570 632188
rect 403342 632176 403348 632188
rect 386564 632148 403348 632176
rect 386564 632136 386570 632148
rect 403342 632136 403348 632148
rect 403400 632136 403406 632188
rect 421282 632136 421288 632188
rect 421340 632176 421346 632188
rect 445018 632176 445024 632188
rect 421340 632148 445024 632176
rect 421340 632136 421346 632148
rect 445018 632136 445024 632148
rect 445076 632136 445082 632188
rect 494514 632136 494520 632188
rect 494572 632176 494578 632188
rect 511350 632176 511356 632188
rect 494572 632148 511356 632176
rect 494572 632136 494578 632148
rect 511350 632136 511356 632148
rect 511408 632136 511414 632188
rect 522298 632136 522304 632188
rect 522356 632176 522362 632188
rect 538398 632176 538404 632188
rect 522356 632148 538404 632176
rect 522356 632136 522362 632148
rect 538398 632136 538404 632148
rect 538456 632136 538462 632188
rect 43346 632068 43352 632120
rect 43404 632108 43410 632120
rect 62758 632108 62764 632120
rect 43404 632080 62764 632108
rect 43404 632068 43410 632080
rect 62758 632068 62764 632080
rect 62816 632068 62822 632120
rect 144178 632068 144184 632120
rect 144236 632108 144242 632120
rect 160278 632108 160284 632120
rect 144236 632080 160284 632108
rect 144236 632068 144242 632080
rect 160278 632068 160284 632080
rect 160336 632068 160342 632120
rect 171778 632068 171784 632120
rect 171836 632108 171842 632120
rect 197446 632108 197452 632120
rect 171836 632080 197452 632108
rect 171836 632068 171842 632080
rect 197446 632068 197452 632080
rect 197504 632068 197510 632120
rect 199378 632068 199384 632120
rect 199436 632108 199442 632120
rect 223942 632108 223948 632120
rect 199436 632080 223948 632108
rect 199436 632068 199442 632080
rect 223942 632068 223948 632080
rect 224000 632068 224006 632120
rect 225598 632068 225604 632120
rect 225656 632108 225662 632120
rect 251174 632108 251180 632120
rect 225656 632080 251180 632108
rect 225656 632068 225662 632080
rect 251174 632068 251180 632080
rect 251232 632068 251238 632120
rect 253198 632068 253204 632120
rect 253256 632108 253262 632120
rect 278038 632108 278044 632120
rect 253256 632080 278044 632108
rect 253256 632068 253262 632080
rect 278038 632068 278044 632080
rect 278096 632068 278102 632120
rect 279510 632068 279516 632120
rect 279568 632108 279574 632120
rect 305546 632108 305552 632120
rect 279568 632080 305552 632108
rect 279568 632068 279574 632080
rect 305546 632068 305552 632080
rect 305604 632068 305610 632120
rect 307018 632068 307024 632120
rect 307076 632108 307082 632120
rect 331950 632108 331956 632120
rect 307076 632080 331956 632108
rect 307076 632068 307082 632080
rect 331950 632068 331956 632080
rect 332008 632068 332014 632120
rect 333238 632068 333244 632120
rect 333296 632108 333302 632120
rect 359458 632108 359464 632120
rect 333296 632080 359464 632108
rect 333296 632068 333302 632080
rect 359458 632068 359464 632080
rect 359516 632068 359522 632120
rect 359734 632068 359740 632120
rect 359792 632108 359798 632120
rect 386046 632108 386052 632120
rect 359792 632080 386052 632108
rect 359792 632068 359798 632080
rect 386046 632068 386052 632080
rect 386104 632068 386110 632120
rect 387058 632068 387064 632120
rect 387116 632108 387122 632120
rect 413002 632108 413008 632120
rect 387116 632080 413008 632108
rect 387116 632068 387122 632080
rect 413002 632068 413008 632080
rect 413060 632068 413066 632120
rect 414658 632068 414664 632120
rect 414716 632108 414722 632120
rect 440234 632108 440240 632120
rect 414716 632080 440240 632108
rect 414716 632068 414722 632080
rect 440234 632068 440240 632080
rect 440292 632068 440298 632120
rect 442258 632068 442264 632120
rect 442316 632108 442322 632120
rect 467006 632108 467012 632120
rect 442316 632080 467012 632108
rect 442316 632068 442322 632080
rect 467006 632068 467012 632080
rect 467064 632068 467070 632120
rect 468478 632068 468484 632120
rect 468536 632108 468542 632120
rect 494054 632108 494060 632120
rect 468536 632080 494060 632108
rect 468536 632068 468542 632080
rect 494054 632068 494060 632080
rect 494112 632068 494118 632120
rect 496078 632068 496084 632120
rect 496136 632108 496142 632120
rect 520918 632108 520924 632120
rect 496136 632080 520924 632108
rect 496136 632068 496142 632080
rect 520918 632068 520924 632080
rect 520976 632068 520982 632120
rect 522390 632068 522396 632120
rect 522448 632108 522454 632120
rect 548058 632108 548064 632120
rect 522448 632080 548064 632108
rect 522448 632068 522454 632080
rect 548058 632068 548064 632080
rect 548116 632068 548122 632120
rect 37918 629892 37924 629944
rect 37976 629932 37982 629944
rect 526438 629932 526444 629944
rect 37976 629904 526444 629932
rect 37976 629892 37982 629904
rect 526438 629892 526444 629904
rect 526496 629892 526502 629944
rect 285766 629280 285772 629332
rect 285824 629320 285830 629332
rect 286134 629320 286140 629332
rect 285824 629292 286140 629320
rect 285824 629280 285830 629292
rect 286134 629280 286140 629292
rect 286192 629280 286198 629332
rect 339586 629280 339592 629332
rect 339644 629320 339650 629332
rect 340138 629320 340144 629332
rect 339644 629292 340144 629320
rect 339644 629280 339650 629292
rect 340138 629280 340144 629292
rect 340196 629280 340202 629332
rect 13722 611260 13728 611312
rect 13780 611300 13786 611312
rect 64874 611300 64880 611312
rect 13780 611272 64880 611300
rect 13780 611260 13786 611272
rect 64874 611260 64880 611272
rect 64932 611260 64938 611312
rect 95142 611260 95148 611312
rect 95200 611300 95206 611312
rect 146294 611300 146300 611312
rect 95200 611272 146300 611300
rect 95200 611260 95206 611272
rect 146294 611260 146300 611272
rect 146352 611260 146358 611312
rect 148962 611260 148968 611312
rect 149020 611300 149026 611312
rect 200114 611300 200120 611312
rect 149020 611272 200120 611300
rect 149020 611260 149026 611272
rect 200114 611260 200120 611272
rect 200172 611260 200178 611312
rect 202782 611260 202788 611312
rect 202840 611300 202846 611312
rect 253934 611300 253940 611312
rect 202840 611272 253940 611300
rect 202840 611260 202846 611272
rect 253934 611260 253940 611272
rect 253992 611260 253998 611312
rect 256602 611260 256608 611312
rect 256660 611300 256666 611312
rect 307754 611300 307760 611312
rect 256660 611272 307760 611300
rect 256660 611260 256666 611272
rect 307754 611260 307760 611272
rect 307812 611260 307818 611312
rect 338022 611260 338028 611312
rect 338080 611300 338086 611312
rect 389174 611300 389180 611312
rect 338080 611272 389180 611300
rect 338080 611260 338086 611272
rect 389174 611260 389180 611272
rect 389232 611260 389238 611312
rect 391842 611260 391848 611312
rect 391900 611300 391906 611312
rect 442994 611300 443000 611312
rect 391900 611272 443000 611300
rect 391900 611260 391906 611272
rect 442994 611260 443000 611272
rect 443052 611260 443058 611312
rect 445662 611260 445668 611312
rect 445720 611300 445726 611312
rect 496814 611300 496820 611312
rect 445720 611272 496820 611300
rect 445720 611260 445726 611272
rect 496814 611260 496820 611272
rect 496872 611260 496878 611312
rect 500862 611260 500868 611312
rect 500920 611300 500926 611312
rect 550634 611300 550640 611312
rect 500920 611272 550640 611300
rect 500920 611260 500926 611272
rect 550634 611260 550640 611272
rect 550692 611260 550698 611312
rect 35618 611192 35624 611244
rect 35676 611232 35682 611244
rect 36722 611232 36728 611244
rect 35676 611204 36728 611232
rect 35676 611192 35682 611204
rect 36722 611192 36728 611204
rect 36780 611192 36786 611244
rect 41322 611192 41328 611244
rect 41380 611232 41386 611244
rect 91094 611232 91100 611244
rect 41380 611204 91100 611232
rect 41380 611192 41386 611204
rect 91094 611192 91100 611204
rect 91152 611192 91158 611244
rect 122742 611192 122748 611244
rect 122800 611232 122806 611244
rect 172514 611232 172520 611244
rect 122800 611204 172520 611232
rect 122800 611192 122806 611204
rect 172514 611192 172520 611204
rect 172572 611192 172578 611244
rect 176562 611192 176568 611244
rect 176620 611232 176626 611244
rect 226334 611232 226340 611244
rect 176620 611204 226340 611232
rect 176620 611192 176626 611204
rect 226334 611192 226340 611204
rect 226392 611192 226398 611244
rect 230382 611192 230388 611244
rect 230440 611232 230446 611244
rect 280154 611232 280160 611244
rect 230440 611204 280160 611232
rect 230440 611192 230446 611204
rect 280154 611192 280160 611204
rect 280212 611192 280218 611244
rect 284202 611192 284208 611244
rect 284260 611232 284266 611244
rect 335354 611232 335360 611244
rect 284260 611204 335360 611232
rect 284260 611192 284266 611204
rect 335354 611192 335360 611204
rect 335412 611192 335418 611244
rect 365622 611192 365628 611244
rect 365680 611232 365686 611244
rect 415394 611232 415400 611244
rect 365680 611204 415400 611232
rect 365680 611192 365686 611204
rect 415394 611192 415400 611204
rect 415452 611192 415458 611244
rect 419442 611192 419448 611244
rect 419500 611232 419506 611244
rect 469214 611232 469220 611244
rect 419500 611204 469220 611232
rect 419500 611192 419506 611204
rect 469214 611192 469220 611204
rect 469272 611192 469278 611244
rect 473262 611192 473268 611244
rect 473320 611232 473326 611244
rect 523034 611232 523040 611244
rect 473320 611204 523040 611232
rect 473320 611192 473326 611204
rect 523034 611192 523040 611204
rect 523092 611192 523098 611244
rect 68922 611124 68928 611176
rect 68980 611164 68986 611176
rect 118694 611164 118700 611176
rect 68980 611136 118700 611164
rect 68980 611124 68986 611136
rect 118694 611124 118700 611136
rect 118752 611124 118758 611176
rect 311802 611124 311808 611176
rect 311860 611164 311866 611176
rect 361574 611164 361580 611176
rect 311860 611136 361580 611164
rect 311860 611124 311866 611136
rect 361574 611124 361580 611136
rect 361632 611124 361638 611176
rect 445018 611124 445024 611176
rect 445076 611164 445082 611176
rect 447686 611164 447692 611176
rect 445076 611136 447692 611164
rect 445076 611124 445082 611136
rect 447686 611124 447692 611136
rect 447744 611124 447750 611176
rect 467650 611124 467656 611176
rect 467708 611164 467714 611176
rect 468570 611164 468576 611176
rect 467708 611136 468576 611164
rect 467708 611124 467714 611136
rect 468570 611124 468576 611136
rect 468628 611124 468634 611176
rect 332594 610648 332600 610700
rect 332652 610688 332658 610700
rect 335998 610688 336004 610700
rect 332652 610660 336004 610688
rect 332652 610648 332658 610660
rect 335998 610648 336004 610660
rect 336056 610648 336062 610700
rect 52730 608540 52736 608592
rect 52788 608580 52794 608592
rect 64138 608580 64144 608592
rect 52788 608552 64144 608580
rect 52788 608540 52794 608552
rect 64138 608540 64144 608552
rect 64196 608540 64202 608592
rect 69106 608540 69112 608592
rect 69164 608580 69170 608592
rect 69164 608552 74534 608580
rect 69164 608540 69170 608552
rect 15194 608472 15200 608524
rect 15252 608512 15258 608524
rect 42978 608512 42984 608524
rect 15252 608484 42984 608512
rect 15252 608472 15258 608484
rect 42978 608472 42984 608484
rect 43036 608472 43042 608524
rect 62758 608472 62764 608524
rect 62816 608512 62822 608524
rect 70026 608512 70032 608524
rect 62816 608484 70032 608512
rect 62816 608472 62822 608484
rect 70026 608472 70032 608484
rect 70084 608472 70090 608524
rect 74506 608512 74534 608552
rect 96706 608540 96712 608592
rect 96764 608580 96770 608592
rect 96764 608552 103514 608580
rect 96764 608540 96770 608552
rect 96982 608512 96988 608524
rect 74506 608484 96988 608512
rect 96982 608472 96988 608484
rect 97040 608472 97046 608524
rect 103486 608512 103514 608552
rect 146938 608540 146944 608592
rect 146996 608580 147002 608592
rect 146996 608552 151814 608580
rect 146996 608540 147002 608552
rect 124030 608512 124036 608524
rect 103486 608484 124036 608512
rect 124030 608472 124036 608484
rect 124088 608472 124094 608524
rect 133690 608472 133696 608524
rect 133748 608512 133754 608524
rect 144270 608512 144276 608524
rect 133748 608484 144276 608512
rect 133748 608472 133754 608484
rect 144270 608472 144276 608484
rect 144328 608472 144334 608524
rect 150526 608472 150532 608524
rect 150584 608512 150590 608524
rect 151786 608512 151814 608552
rect 200758 608540 200764 608592
rect 200816 608580 200822 608592
rect 204990 608580 204996 608592
rect 200816 608552 204996 608580
rect 200816 608540 200822 608552
rect 204990 608540 204996 608552
rect 205048 608540 205054 608592
rect 251818 608540 251824 608592
rect 251876 608580 251882 608592
rect 258994 608580 259000 608592
rect 251876 608552 259000 608580
rect 251876 608540 251882 608552
rect 258994 608540 259000 608552
rect 259052 608540 259058 608592
rect 494698 608540 494704 608592
rect 494756 608580 494762 608592
rect 501966 608580 501972 608592
rect 494756 608552 501972 608580
rect 494756 608540 494762 608552
rect 501966 608540 501972 608552
rect 502024 608540 502030 608592
rect 548334 608512 548340 608524
rect 150584 608484 151124 608512
rect 151786 608484 548340 608512
rect 150584 608472 150590 608484
rect 25682 608404 25688 608456
rect 25740 608444 25746 608456
rect 36814 608444 36820 608456
rect 25740 608416 36820 608444
rect 25740 608404 25746 608416
rect 36814 608404 36820 608416
rect 36872 608404 36878 608456
rect 79686 608404 79692 608456
rect 79744 608444 79750 608456
rect 90450 608444 90456 608456
rect 79744 608416 90456 608444
rect 79744 608404 79750 608416
rect 90450 608404 90456 608416
rect 90508 608404 90514 608456
rect 106642 608404 106648 608456
rect 106700 608444 106706 608456
rect 116578 608444 116584 608456
rect 106700 608416 116584 608444
rect 106700 608404 106706 608416
rect 116578 608404 116584 608416
rect 116636 608404 116642 608456
rect 122926 608404 122932 608456
rect 122984 608444 122990 608456
rect 150986 608444 150992 608456
rect 122984 608416 150992 608444
rect 122984 608404 122990 608416
rect 150986 608404 150992 608416
rect 151044 608404 151050 608456
rect 151096 608444 151124 608484
rect 548334 608472 548340 608484
rect 548392 608472 548398 608524
rect 178034 608444 178040 608456
rect 151096 608416 178040 608444
rect 178034 608404 178040 608416
rect 178092 608404 178098 608456
rect 187694 608404 187700 608456
rect 187752 608444 187758 608456
rect 199378 608444 199384 608456
rect 187752 608416 199384 608444
rect 187752 608404 187758 608416
rect 199378 608404 199384 608416
rect 199436 608404 199442 608456
rect 204346 608404 204352 608456
rect 204404 608444 204410 608456
rect 232038 608444 232044 608456
rect 204404 608416 232044 608444
rect 204404 608404 204410 608416
rect 232038 608404 232044 608416
rect 232096 608404 232102 608456
rect 241698 608404 241704 608456
rect 241756 608444 241762 608456
rect 253198 608444 253204 608456
rect 241756 608416 253204 608444
rect 241756 608404 241762 608416
rect 253198 608404 253204 608416
rect 253256 608404 253262 608456
rect 258166 608404 258172 608456
rect 258224 608444 258230 608456
rect 286042 608444 286048 608456
rect 258224 608416 286048 608444
rect 258224 608404 258230 608416
rect 286042 608404 286048 608416
rect 286100 608404 286106 608456
rect 312998 608444 313004 608456
rect 287026 608416 313004 608444
rect 160646 608336 160652 608388
rect 160704 608376 160710 608388
rect 171778 608376 171784 608388
rect 160704 608348 171784 608376
rect 160704 608336 160710 608348
rect 171778 608336 171784 608348
rect 171836 608336 171842 608388
rect 214650 608336 214656 608388
rect 214708 608376 214714 608388
rect 225598 608376 225604 608388
rect 214708 608348 225604 608376
rect 214708 608336 214714 608348
rect 225598 608336 225604 608348
rect 225656 608336 225662 608388
rect 268654 608336 268660 608388
rect 268712 608376 268718 608388
rect 279510 608376 279516 608388
rect 268712 608348 279516 608376
rect 268712 608336 268718 608348
rect 279510 608336 279516 608348
rect 279568 608336 279574 608388
rect 285766 608336 285772 608388
rect 285824 608376 285830 608388
rect 287026 608376 287054 608416
rect 312998 608404 313004 608416
rect 313056 608404 313062 608456
rect 340046 608444 340052 608456
rect 316006 608416 340052 608444
rect 285824 608348 287054 608376
rect 285824 608336 285830 608348
rect 295702 608336 295708 608388
rect 295760 608376 295766 608388
rect 307018 608376 307024 608388
rect 295760 608348 307024 608376
rect 295760 608336 295766 608348
rect 307018 608336 307024 608348
rect 307076 608336 307082 608388
rect 311986 608336 311992 608388
rect 312044 608376 312050 608388
rect 316006 608376 316034 608416
rect 340046 608404 340052 608416
rect 340104 608404 340110 608456
rect 367002 608444 367008 608456
rect 344986 608416 367008 608444
rect 312044 608348 316034 608376
rect 312044 608336 312050 608348
rect 322658 608336 322664 608388
rect 322716 608376 322722 608388
rect 333238 608376 333244 608388
rect 322716 608348 333244 608376
rect 322716 608336 322722 608348
rect 333238 608336 333244 608348
rect 333296 608336 333302 608388
rect 339586 608336 339592 608388
rect 339644 608376 339650 608388
rect 344986 608376 345014 608416
rect 367002 608404 367008 608416
rect 367060 608404 367066 608456
rect 393958 608444 393964 608456
rect 373966 608416 393964 608444
rect 339644 608348 345014 608376
rect 339644 608336 339650 608348
rect 349706 608336 349712 608388
rect 349764 608376 349770 608388
rect 359550 608376 359556 608388
rect 349764 608348 359556 608376
rect 349764 608336 349770 608348
rect 359550 608336 359556 608348
rect 359608 608336 359614 608388
rect 365806 608336 365812 608388
rect 365864 608376 365870 608388
rect 373966 608376 373994 608416
rect 393958 608404 393964 608416
rect 394016 608404 394022 608456
rect 421006 608444 421012 608456
rect 402946 608416 421012 608444
rect 365864 608348 373994 608376
rect 365864 608336 365870 608348
rect 376662 608336 376668 608388
rect 376720 608376 376726 608388
rect 387058 608376 387064 608388
rect 376720 608348 387064 608376
rect 376720 608336 376726 608348
rect 387058 608336 387064 608348
rect 387116 608336 387122 608388
rect 393406 608336 393412 608388
rect 393464 608376 393470 608388
rect 402946 608376 402974 608416
rect 421006 608404 421012 608416
rect 421064 608404 421070 608456
rect 430666 608404 430672 608456
rect 430724 608444 430730 608456
rect 442258 608444 442264 608456
rect 430724 608416 442264 608444
rect 430724 608404 430730 608416
rect 442258 608404 442264 608416
rect 442316 608404 442322 608456
rect 447226 608404 447232 608456
rect 447284 608444 447290 608456
rect 475010 608444 475016 608456
rect 447284 608416 475016 608444
rect 447284 608404 447290 608416
rect 475010 608404 475016 608416
rect 475068 608404 475074 608456
rect 484670 608404 484676 608456
rect 484728 608444 484734 608456
rect 496078 608444 496084 608456
rect 484728 608416 496084 608444
rect 484728 608404 484734 608416
rect 496078 608404 496084 608416
rect 496136 608404 496142 608456
rect 501046 608404 501052 608456
rect 501104 608444 501110 608456
rect 529014 608444 529020 608456
rect 501104 608416 529020 608444
rect 501104 608404 501110 608416
rect 529014 608404 529020 608416
rect 529072 608404 529078 608456
rect 393464 608348 402974 608376
rect 393464 608336 393470 608348
rect 403710 608336 403716 608388
rect 403768 608376 403774 608388
rect 414658 608376 414664 608388
rect 403768 608348 414664 608376
rect 403768 608336 403774 608348
rect 414658 608336 414664 608348
rect 414716 608336 414722 608388
rect 457714 608336 457720 608388
rect 457772 608376 457778 608388
rect 468478 608376 468484 608388
rect 457772 608348 468484 608376
rect 457772 608336 457778 608348
rect 468478 608336 468484 608348
rect 468536 608336 468542 608388
rect 511718 608336 511724 608388
rect 511776 608376 511782 608388
rect 522390 608376 522396 608388
rect 511776 608348 522396 608376
rect 511776 608336 511782 608348
rect 522390 608336 522396 608348
rect 522448 608336 522454 608388
rect 36630 608268 36636 608320
rect 36688 608308 36694 608320
rect 538674 608308 538680 608320
rect 36688 608280 538680 608308
rect 36688 608268 36694 608280
rect 538674 608268 538680 608280
rect 538732 608268 538738 608320
rect 15286 605072 15292 605124
rect 15344 605112 15350 605124
rect 529014 605112 529020 605124
rect 15344 605084 529020 605112
rect 15344 605072 15350 605084
rect 529014 605072 529020 605084
rect 529072 605072 529078 605124
rect 25682 604732 25688 604784
rect 25740 604772 25746 604784
rect 146938 604772 146944 604784
rect 25740 604744 146944 604772
rect 25740 604732 25746 604744
rect 146938 604732 146944 604744
rect 146996 604732 147002 604784
rect 36722 604664 36728 604716
rect 36780 604704 36786 604716
rect 52638 604704 52644 604716
rect 36780 604676 52644 604704
rect 36780 604664 36786 604676
rect 52638 604664 52644 604676
rect 52696 604664 52702 604716
rect 232038 604664 232044 604716
rect 232096 604704 232102 604716
rect 251818 604704 251824 604716
rect 232096 604676 251824 604704
rect 232096 604664 232102 604676
rect 251818 604664 251824 604676
rect 251876 604664 251882 604716
rect 475010 604664 475016 604716
rect 475068 604704 475074 604716
rect 494698 604704 494704 604716
rect 475068 604676 494704 604704
rect 475068 604664 475074 604676
rect 494698 604664 494704 604676
rect 494756 604664 494762 604716
rect 62482 604596 62488 604648
rect 62540 604636 62546 604648
rect 79686 604636 79692 604648
rect 62540 604608 79692 604636
rect 62540 604596 62546 604608
rect 79686 604596 79692 604608
rect 79744 604596 79750 604648
rect 90450 604596 90456 604648
rect 90508 604636 90514 604648
rect 106642 604636 106648 604648
rect 90508 604608 106648 604636
rect 90508 604596 90514 604608
rect 106642 604596 106648 604608
rect 106700 604596 106706 604648
rect 116486 604596 116492 604648
rect 116544 604636 116550 604648
rect 133690 604636 133696 604648
rect 116544 604608 133696 604636
rect 116544 604596 116550 604608
rect 133690 604596 133696 604608
rect 133748 604596 133754 604648
rect 170490 604596 170496 604648
rect 170548 604636 170554 604648
rect 187694 604636 187700 604648
rect 170548 604608 187700 604636
rect 170548 604596 170554 604608
rect 187694 604596 187700 604608
rect 187752 604596 187758 604648
rect 197446 604596 197452 604648
rect 197504 604636 197510 604648
rect 214650 604636 214656 604648
rect 197504 604608 214656 604636
rect 197504 604596 197510 604608
rect 214650 604596 214656 604608
rect 214708 604596 214714 604648
rect 224494 604596 224500 604648
rect 224552 604636 224558 604648
rect 241698 604636 241704 604648
rect 224552 604608 241704 604636
rect 224552 604596 224558 604608
rect 241698 604596 241704 604608
rect 241756 604596 241762 604648
rect 413462 604596 413468 604648
rect 413520 604636 413526 604648
rect 430666 604636 430672 604648
rect 413520 604608 430672 604636
rect 413520 604596 413526 604608
rect 430666 604596 430672 604608
rect 430724 604596 430730 604648
rect 440510 604596 440516 604648
rect 440568 604636 440574 604648
rect 457622 604636 457628 604648
rect 440568 604608 457628 604636
rect 440568 604596 440574 604608
rect 457622 604596 457628 604608
rect 457680 604596 457686 604648
rect 468570 604596 468576 604648
rect 468628 604636 468634 604648
rect 484670 604636 484676 604648
rect 468628 604608 484676 604636
rect 468628 604596 468634 604608
rect 484670 604596 484676 604608
rect 484728 604596 484734 604648
rect 36814 604528 36820 604580
rect 36872 604568 36878 604580
rect 62298 604568 62304 604580
rect 36872 604540 62304 604568
rect 36872 604528 36878 604540
rect 62298 604528 62304 604540
rect 62356 604528 62362 604580
rect 64138 604528 64144 604580
rect 64196 604568 64202 604580
rect 89346 604568 89352 604580
rect 64196 604540 89352 604568
rect 64196 604528 64202 604540
rect 89346 604528 89352 604540
rect 89404 604528 89410 604580
rect 90358 604528 90364 604580
rect 90416 604568 90422 604580
rect 116302 604568 116308 604580
rect 90416 604540 116308 604568
rect 90416 604528 90422 604540
rect 116302 604528 116308 604540
rect 116360 604528 116366 604580
rect 116578 604528 116584 604580
rect 116636 604568 116642 604580
rect 143350 604568 143356 604580
rect 116636 604540 143356 604568
rect 116636 604528 116642 604540
rect 143350 604528 143356 604540
rect 143408 604528 143414 604580
rect 144270 604528 144276 604580
rect 144328 604568 144334 604580
rect 170306 604568 170312 604580
rect 144328 604540 170312 604568
rect 144328 604528 144334 604540
rect 170306 604528 170312 604540
rect 170364 604528 170370 604580
rect 178034 604528 178040 604580
rect 178092 604568 178098 604580
rect 200758 604568 200764 604580
rect 178092 604540 200764 604568
rect 178092 604528 178098 604540
rect 200758 604528 200764 604540
rect 200816 604528 200822 604580
rect 251450 604528 251456 604580
rect 251508 604568 251514 604580
rect 268654 604568 268660 604580
rect 251508 604540 268660 604568
rect 251508 604528 251514 604540
rect 268654 604528 268660 604540
rect 268712 604528 268718 604580
rect 279510 604528 279516 604580
rect 279568 604568 279574 604580
rect 295702 604568 295708 604580
rect 279568 604540 295708 604568
rect 279568 604528 279574 604540
rect 295702 604528 295708 604540
rect 295760 604528 295766 604580
rect 305454 604528 305460 604580
rect 305512 604568 305518 604580
rect 322658 604568 322664 604580
rect 305512 604540 322664 604568
rect 305512 604528 305518 604540
rect 322658 604528 322664 604540
rect 322716 604528 322722 604580
rect 335998 604528 336004 604580
rect 336056 604568 336062 604580
rect 349706 604568 349712 604580
rect 336056 604540 349712 604568
rect 336056 604528 336062 604540
rect 349706 604528 349712 604540
rect 349764 604528 349770 604580
rect 359458 604528 359464 604580
rect 359516 604568 359522 604580
rect 376662 604568 376668 604580
rect 359516 604540 376668 604568
rect 359516 604528 359522 604540
rect 376662 604528 376668 604540
rect 376720 604528 376726 604580
rect 386506 604528 386512 604580
rect 386564 604568 386570 604580
rect 403618 604568 403624 604580
rect 386564 604540 403624 604568
rect 386564 604528 386570 604540
rect 403618 604528 403624 604540
rect 403676 604528 403682 604580
rect 421006 604528 421012 604580
rect 421064 604568 421070 604580
rect 445018 604568 445024 604580
rect 421064 604540 445024 604568
rect 421064 604528 421070 604540
rect 445018 604528 445024 604540
rect 445076 604528 445082 604580
rect 494514 604528 494520 604580
rect 494572 604568 494578 604580
rect 511626 604568 511632 604580
rect 494572 604540 511632 604568
rect 494572 604528 494578 604540
rect 511626 604528 511632 604540
rect 511684 604528 511690 604580
rect 522298 604528 522304 604580
rect 522356 604568 522362 604580
rect 538674 604568 538680 604580
rect 522356 604540 538680 604568
rect 522356 604528 522362 604540
rect 538674 604528 538680 604540
rect 538732 604528 538738 604580
rect 43070 604460 43076 604512
rect 43128 604500 43134 604512
rect 62758 604500 62764 604512
rect 43128 604472 62764 604500
rect 43128 604460 43134 604472
rect 62758 604460 62764 604472
rect 62816 604460 62822 604512
rect 144178 604460 144184 604512
rect 144236 604500 144242 604512
rect 160646 604500 160652 604512
rect 144236 604472 160652 604500
rect 144236 604460 144242 604472
rect 160646 604460 160652 604472
rect 160704 604460 160710 604512
rect 171778 604460 171784 604512
rect 171836 604500 171842 604512
rect 197354 604500 197360 604512
rect 171836 604472 197360 604500
rect 171836 604460 171842 604472
rect 197354 604460 197360 604472
rect 197412 604460 197418 604512
rect 199378 604460 199384 604512
rect 199436 604500 199442 604512
rect 224310 604500 224316 604512
rect 199436 604472 224316 604500
rect 199436 604460 199442 604472
rect 224310 604460 224316 604472
rect 224368 604460 224374 604512
rect 225598 604460 225604 604512
rect 225656 604500 225662 604512
rect 251358 604500 251364 604512
rect 225656 604472 251364 604500
rect 225656 604460 225662 604472
rect 251358 604460 251364 604472
rect 251416 604460 251422 604512
rect 253198 604460 253204 604512
rect 253256 604500 253262 604512
rect 278314 604500 278320 604512
rect 253256 604472 278320 604500
rect 253256 604460 253262 604472
rect 278314 604460 278320 604472
rect 278372 604460 278378 604512
rect 279418 604460 279424 604512
rect 279476 604500 279482 604512
rect 305362 604500 305368 604512
rect 279476 604472 305368 604500
rect 279476 604460 279482 604472
rect 305362 604460 305368 604472
rect 305420 604460 305426 604512
rect 307018 604460 307024 604512
rect 307076 604500 307082 604512
rect 332318 604500 332324 604512
rect 307076 604472 332324 604500
rect 307076 604460 307082 604472
rect 332318 604460 332324 604472
rect 332376 604460 332382 604512
rect 333238 604460 333244 604512
rect 333296 604500 333302 604512
rect 359366 604500 359372 604512
rect 333296 604472 359372 604500
rect 333296 604460 333302 604472
rect 359366 604460 359372 604472
rect 359424 604460 359430 604512
rect 359550 604460 359556 604512
rect 359608 604500 359614 604512
rect 386322 604500 386328 604512
rect 359608 604472 386328 604500
rect 359608 604460 359614 604472
rect 386322 604460 386328 604472
rect 386380 604460 386386 604512
rect 387058 604460 387064 604512
rect 387116 604500 387122 604512
rect 413278 604500 413284 604512
rect 387116 604472 413284 604500
rect 387116 604460 387122 604472
rect 413278 604460 413284 604472
rect 413336 604460 413342 604512
rect 414658 604460 414664 604512
rect 414716 604500 414722 604512
rect 440326 604500 440332 604512
rect 414716 604472 440332 604500
rect 414716 604460 414722 604472
rect 440326 604460 440332 604472
rect 440384 604460 440390 604512
rect 442258 604460 442264 604512
rect 442316 604500 442322 604512
rect 467282 604500 467288 604512
rect 442316 604472 467288 604500
rect 442316 604460 442322 604472
rect 467282 604460 467288 604472
rect 467340 604460 467346 604512
rect 468478 604460 468484 604512
rect 468536 604500 468542 604512
rect 494330 604500 494336 604512
rect 468536 604472 494336 604500
rect 468536 604460 468542 604472
rect 494330 604460 494336 604472
rect 494388 604460 494394 604512
rect 496078 604460 496084 604512
rect 496136 604500 496142 604512
rect 521286 604500 521292 604512
rect 496136 604472 521292 604500
rect 496136 604460 496142 604472
rect 521286 604460 521292 604472
rect 521344 604460 521350 604512
rect 522390 604460 522396 604512
rect 522448 604500 522454 604512
rect 548334 604500 548340 604512
rect 522448 604472 548340 604500
rect 522448 604460 522454 604472
rect 548334 604460 548340 604472
rect 548392 604460 548398 604512
rect 37918 602352 37924 602404
rect 37976 602392 37982 602404
rect 526438 602392 526444 602404
rect 37976 602364 526444 602392
rect 37976 602352 37982 602364
rect 526438 602352 526444 602364
rect 526496 602352 526502 602404
rect 35618 601672 35624 601724
rect 35676 601712 35682 601724
rect 36630 601712 36636 601724
rect 35676 601684 36636 601712
rect 35676 601672 35682 601684
rect 36630 601672 36636 601684
rect 36688 601672 36694 601724
rect 278774 584740 278780 584792
rect 278832 584780 278838 584792
rect 279510 584780 279516 584792
rect 278832 584752 279516 584780
rect 278832 584740 278838 584752
rect 279510 584740 279516 584752
rect 279568 584740 279574 584792
rect 445018 583720 445024 583772
rect 445076 583760 445082 583772
rect 447686 583760 447692 583772
rect 445076 583732 447692 583760
rect 445076 583720 445082 583732
rect 447686 583720 447692 583732
rect 447744 583720 447750 583772
rect 13722 583652 13728 583704
rect 13780 583692 13786 583704
rect 64874 583692 64880 583704
rect 13780 583664 64880 583692
rect 13780 583652 13786 583664
rect 64874 583652 64880 583664
rect 64932 583652 64938 583704
rect 89714 583652 89720 583704
rect 89772 583692 89778 583704
rect 90450 583692 90456 583704
rect 89772 583664 90456 583692
rect 89772 583652 89778 583664
rect 90450 583652 90456 583664
rect 90508 583652 90514 583704
rect 95142 583652 95148 583704
rect 95200 583692 95206 583704
rect 146294 583692 146300 583704
rect 95200 583664 146300 583692
rect 95200 583652 95206 583664
rect 146294 583652 146300 583664
rect 146352 583652 146358 583704
rect 148962 583652 148968 583704
rect 149020 583692 149026 583704
rect 200114 583692 200120 583704
rect 149020 583664 200120 583692
rect 149020 583652 149026 583664
rect 200114 583652 200120 583664
rect 200172 583652 200178 583704
rect 202782 583652 202788 583704
rect 202840 583692 202846 583704
rect 253934 583692 253940 583704
rect 202840 583664 253940 583692
rect 202840 583652 202846 583664
rect 253934 583652 253940 583664
rect 253992 583652 253998 583704
rect 256602 583652 256608 583704
rect 256660 583692 256666 583704
rect 307754 583692 307760 583704
rect 256660 583664 307760 583692
rect 256660 583652 256666 583664
rect 307754 583652 307760 583664
rect 307812 583652 307818 583704
rect 332594 583652 332600 583704
rect 332652 583692 332658 583704
rect 335998 583692 336004 583704
rect 332652 583664 336004 583692
rect 332652 583652 332658 583664
rect 335998 583652 336004 583664
rect 336056 583652 336062 583704
rect 338022 583652 338028 583704
rect 338080 583692 338086 583704
rect 389174 583692 389180 583704
rect 338080 583664 389180 583692
rect 338080 583652 338086 583664
rect 389174 583652 389180 583664
rect 389232 583652 389238 583704
rect 391842 583652 391848 583704
rect 391900 583692 391906 583704
rect 442994 583692 443000 583704
rect 391900 583664 443000 583692
rect 391900 583652 391906 583664
rect 442994 583652 443000 583664
rect 443052 583652 443058 583704
rect 445662 583652 445668 583704
rect 445720 583692 445726 583704
rect 496814 583692 496820 583704
rect 445720 583664 496820 583692
rect 445720 583652 445726 583664
rect 496814 583652 496820 583664
rect 496872 583652 496878 583704
rect 500862 583652 500868 583704
rect 500920 583692 500926 583704
rect 550634 583692 550640 583704
rect 500920 583664 550640 583692
rect 500920 583652 500926 583664
rect 550634 583652 550640 583664
rect 550692 583652 550698 583704
rect 35618 583584 35624 583636
rect 35676 583624 35682 583636
rect 36722 583624 36728 583636
rect 35676 583596 36728 583624
rect 35676 583584 35682 583596
rect 36722 583584 36728 583596
rect 36780 583584 36786 583636
rect 41322 583584 41328 583636
rect 41380 583624 41386 583636
rect 91094 583624 91100 583636
rect 41380 583596 91100 583624
rect 41380 583584 41386 583596
rect 91094 583584 91100 583596
rect 91152 583584 91158 583636
rect 116210 583584 116216 583636
rect 116268 583624 116274 583636
rect 116486 583624 116492 583636
rect 116268 583596 116492 583624
rect 116268 583584 116274 583596
rect 116486 583584 116492 583596
rect 116544 583584 116550 583636
rect 122742 583584 122748 583636
rect 122800 583624 122806 583636
rect 172514 583624 172520 583636
rect 122800 583596 172520 583624
rect 122800 583584 122806 583596
rect 172514 583584 172520 583596
rect 172572 583584 172578 583636
rect 176562 583584 176568 583636
rect 176620 583624 176626 583636
rect 226334 583624 226340 583636
rect 176620 583596 226340 583624
rect 176620 583584 176626 583596
rect 226334 583584 226340 583596
rect 226392 583584 226398 583636
rect 230382 583584 230388 583636
rect 230440 583624 230446 583636
rect 280154 583624 280160 583636
rect 230440 583596 280160 583624
rect 230440 583584 230446 583596
rect 280154 583584 280160 583596
rect 280212 583584 280218 583636
rect 284202 583584 284208 583636
rect 284260 583624 284266 583636
rect 335354 583624 335360 583636
rect 284260 583596 335360 583624
rect 284260 583584 284266 583596
rect 335354 583584 335360 583596
rect 335412 583584 335418 583636
rect 365622 583584 365628 583636
rect 365680 583624 365686 583636
rect 415394 583624 415400 583636
rect 365680 583596 415400 583624
rect 365680 583584 365686 583596
rect 415394 583584 415400 583596
rect 415452 583584 415458 583636
rect 419442 583584 419448 583636
rect 419500 583624 419506 583636
rect 469214 583624 469220 583636
rect 419500 583596 469220 583624
rect 419500 583584 419506 583596
rect 469214 583584 469220 583596
rect 469272 583584 469278 583636
rect 473262 583584 473268 583636
rect 473320 583624 473326 583636
rect 523034 583624 523040 583636
rect 473320 583596 523040 583624
rect 473320 583584 473326 583596
rect 523034 583584 523040 583596
rect 523092 583584 523098 583636
rect 68922 583516 68928 583568
rect 68980 583556 68986 583568
rect 118694 583556 118700 583568
rect 68980 583528 118700 583556
rect 68980 583516 68986 583528
rect 118694 583516 118700 583528
rect 118752 583516 118758 583568
rect 170214 583516 170220 583568
rect 170272 583556 170278 583568
rect 170490 583556 170496 583568
rect 170272 583528 170496 583556
rect 170272 583516 170278 583528
rect 170490 583516 170496 583528
rect 170548 583516 170554 583568
rect 200758 583516 200764 583568
rect 200816 583556 200822 583568
rect 204622 583556 204628 583568
rect 200816 583528 204628 583556
rect 200816 583516 200822 583528
rect 204622 583516 204628 583528
rect 204680 583516 204686 583568
rect 311802 583516 311808 583568
rect 311860 583556 311866 583568
rect 361574 583556 361580 583568
rect 311860 583528 361580 583556
rect 311860 583516 311866 583528
rect 361574 583516 361580 583528
rect 361632 583516 361638 583568
rect 467650 583516 467656 583568
rect 467708 583556 467714 583568
rect 468570 583556 468576 583568
rect 467708 583528 468576 583556
rect 467708 583516 467714 583528
rect 468570 583516 468576 583528
rect 468628 583516 468634 583568
rect 62758 580932 62764 580984
rect 62816 580972 62822 580984
rect 69750 580972 69756 580984
rect 62816 580944 69756 580972
rect 62816 580932 62822 580944
rect 69750 580932 69756 580944
rect 69808 580932 69814 580984
rect 96706 580932 96712 580984
rect 96764 580972 96770 580984
rect 96764 580944 103514 580972
rect 96764 580932 96770 580944
rect 15194 580864 15200 580916
rect 15252 580904 15258 580916
rect 42794 580904 42800 580916
rect 15252 580876 42800 580904
rect 15252 580864 15258 580876
rect 42794 580864 42800 580876
rect 42852 580864 42858 580916
rect 53098 580864 53104 580916
rect 53156 580904 53162 580916
rect 64138 580904 64144 580916
rect 53156 580876 64144 580904
rect 53156 580864 53162 580876
rect 64138 580864 64144 580876
rect 64196 580864 64202 580916
rect 69106 580864 69112 580916
rect 69164 580904 69170 580916
rect 96798 580904 96804 580916
rect 69164 580876 96804 580904
rect 69164 580864 69170 580876
rect 96798 580864 96804 580876
rect 96856 580864 96862 580916
rect 103486 580904 103514 580944
rect 251818 580932 251824 580984
rect 251876 580972 251882 580984
rect 258718 580972 258724 580984
rect 251876 580944 258724 580972
rect 251876 580932 251882 580944
rect 258718 580932 258724 580944
rect 258776 580932 258782 580984
rect 494698 580932 494704 580984
rect 494756 580972 494762 580984
rect 501598 580972 501604 580984
rect 494756 580944 501604 580972
rect 494756 580932 494762 580944
rect 501598 580932 501604 580944
rect 501656 580932 501662 580984
rect 123662 580904 123668 580916
rect 103486 580876 123668 580904
rect 123662 580864 123668 580876
rect 123720 580864 123726 580916
rect 148318 580864 148324 580916
rect 148376 580904 148382 580916
rect 548058 580904 548064 580916
rect 148376 580876 548064 580904
rect 148376 580864 148382 580876
rect 548058 580864 548064 580876
rect 548116 580864 548122 580916
rect 25958 580796 25964 580848
rect 26016 580836 26022 580848
rect 36814 580836 36820 580848
rect 26016 580808 36820 580836
rect 26016 580796 26022 580808
rect 36814 580796 36820 580808
rect 36872 580796 36878 580848
rect 79962 580796 79968 580848
rect 80020 580836 80026 580848
rect 90358 580836 90364 580848
rect 80020 580808 90364 580836
rect 80020 580796 80026 580808
rect 90358 580796 90364 580808
rect 90416 580796 90422 580848
rect 106550 580796 106556 580848
rect 106608 580836 106614 580848
rect 116578 580836 116584 580848
rect 106608 580808 116584 580836
rect 106608 580796 106614 580808
rect 116578 580796 116584 580808
rect 116636 580796 116642 580848
rect 133782 580796 133788 580848
rect 133840 580836 133846 580848
rect 144270 580836 144276 580848
rect 133840 580808 144276 580836
rect 133840 580796 133846 580808
rect 144270 580796 144276 580808
rect 144328 580796 144334 580848
rect 150526 580796 150532 580848
rect 150584 580836 150590 580848
rect 178126 580836 178132 580848
rect 150584 580808 178132 580836
rect 150584 580796 150590 580808
rect 178126 580796 178132 580808
rect 178184 580796 178190 580848
rect 187970 580796 187976 580848
rect 188028 580836 188034 580848
rect 199378 580836 199384 580848
rect 188028 580808 199384 580836
rect 188028 580796 188034 580808
rect 199378 580796 199384 580808
rect 199436 580796 199442 580848
rect 204346 580796 204352 580848
rect 204404 580836 204410 580848
rect 231854 580836 231860 580848
rect 204404 580808 231860 580836
rect 204404 580796 204410 580808
rect 231854 580796 231860 580808
rect 231912 580796 231918 580848
rect 242066 580796 242072 580848
rect 242124 580836 242130 580848
rect 253198 580836 253204 580848
rect 242124 580808 253204 580836
rect 242124 580796 242130 580808
rect 253198 580796 253204 580808
rect 253256 580796 253262 580848
rect 258166 580796 258172 580848
rect 258224 580836 258230 580848
rect 286134 580836 286140 580848
rect 258224 580808 286140 580836
rect 258224 580796 258230 580808
rect 286134 580796 286140 580808
rect 286192 580796 286198 580848
rect 312630 580836 312636 580848
rect 287026 580808 312636 580836
rect 122926 580728 122932 580780
rect 122984 580768 122990 580780
rect 150710 580768 150716 580780
rect 122984 580740 150716 580768
rect 122984 580728 122990 580740
rect 150710 580728 150716 580740
rect 150768 580728 150774 580780
rect 160554 580728 160560 580780
rect 160612 580768 160618 580780
rect 171778 580768 171784 580780
rect 160612 580740 171784 580768
rect 160612 580728 160618 580740
rect 171778 580728 171784 580740
rect 171836 580728 171842 580780
rect 215018 580728 215024 580780
rect 215076 580768 215082 580780
rect 225598 580768 225604 580780
rect 215076 580740 225604 580768
rect 215076 580728 215082 580740
rect 225598 580728 225604 580740
rect 225656 580728 225662 580780
rect 268930 580728 268936 580780
rect 268988 580768 268994 580780
rect 279418 580768 279424 580780
rect 268988 580740 279424 580768
rect 268988 580728 268994 580740
rect 279418 580728 279424 580740
rect 279476 580728 279482 580780
rect 285766 580728 285772 580780
rect 285824 580768 285830 580780
rect 287026 580768 287054 580808
rect 312630 580796 312636 580808
rect 312688 580796 312694 580848
rect 340138 580836 340144 580848
rect 316006 580808 340144 580836
rect 285824 580740 287054 580768
rect 285824 580728 285830 580740
rect 295978 580728 295984 580780
rect 296036 580768 296042 580780
rect 307018 580768 307024 580780
rect 296036 580740 307024 580768
rect 296036 580728 296042 580740
rect 307018 580728 307024 580740
rect 307076 580728 307082 580780
rect 311986 580728 311992 580780
rect 312044 580768 312050 580780
rect 316006 580768 316034 580808
rect 340138 580796 340144 580808
rect 340196 580796 340202 580848
rect 366726 580836 366732 580848
rect 344986 580808 366732 580836
rect 312044 580740 316034 580768
rect 312044 580728 312050 580740
rect 322842 580728 322848 580780
rect 322900 580768 322906 580780
rect 333238 580768 333244 580780
rect 322900 580740 333244 580768
rect 322900 580728 322906 580740
rect 333238 580728 333244 580740
rect 333296 580728 333302 580780
rect 339586 580728 339592 580780
rect 339644 580768 339650 580780
rect 344986 580768 345014 580808
rect 366726 580796 366732 580808
rect 366784 580796 366790 580848
rect 393590 580836 393596 580848
rect 373966 580808 393596 580836
rect 339644 580740 345014 580768
rect 339644 580728 339650 580740
rect 350074 580728 350080 580780
rect 350132 580768 350138 580780
rect 359550 580768 359556 580780
rect 350132 580740 359556 580768
rect 350132 580728 350138 580740
rect 359550 580728 359556 580740
rect 359608 580728 359614 580780
rect 365806 580728 365812 580780
rect 365864 580768 365870 580780
rect 373966 580768 373994 580808
rect 393590 580796 393596 580808
rect 393648 580796 393654 580848
rect 420914 580836 420920 580848
rect 402946 580808 420920 580836
rect 365864 580740 373994 580768
rect 365864 580728 365870 580740
rect 376570 580728 376576 580780
rect 376628 580768 376634 580780
rect 387058 580768 387064 580780
rect 376628 580740 387064 580768
rect 376628 580728 376634 580740
rect 387058 580728 387064 580740
rect 387116 580728 387122 580780
rect 393406 580728 393412 580780
rect 393464 580768 393470 580780
rect 402946 580768 402974 580808
rect 420914 580796 420920 580808
rect 420972 580796 420978 580848
rect 431034 580796 431040 580848
rect 431092 580836 431098 580848
rect 442258 580836 442264 580848
rect 431092 580808 442264 580836
rect 431092 580796 431098 580808
rect 442258 580796 442264 580808
rect 442316 580796 442322 580848
rect 447226 580796 447232 580848
rect 447284 580836 447290 580848
rect 474734 580836 474740 580848
rect 447284 580808 474740 580836
rect 447284 580796 447290 580808
rect 474734 580796 474740 580808
rect 474792 580796 474798 580848
rect 484946 580796 484952 580848
rect 485004 580836 485010 580848
rect 496078 580836 496084 580848
rect 485004 580808 496084 580836
rect 485004 580796 485010 580808
rect 496078 580796 496084 580808
rect 496136 580796 496142 580848
rect 501046 580796 501052 580848
rect 501104 580836 501110 580848
rect 528738 580836 528744 580848
rect 501104 580808 528744 580836
rect 501104 580796 501110 580808
rect 528738 580796 528744 580808
rect 528796 580796 528802 580848
rect 393464 580740 402974 580768
rect 393464 580728 393470 580740
rect 403986 580728 403992 580780
rect 404044 580768 404050 580780
rect 414658 580768 414664 580780
rect 404044 580740 414664 580768
rect 404044 580728 404050 580740
rect 414658 580728 414664 580740
rect 414716 580728 414722 580780
rect 458082 580728 458088 580780
rect 458140 580768 458146 580780
rect 468478 580768 468484 580780
rect 458140 580740 468484 580768
rect 458140 580728 458146 580740
rect 468478 580728 468484 580740
rect 468536 580728 468542 580780
rect 511902 580728 511908 580780
rect 511960 580768 511966 580780
rect 522390 580768 522396 580780
rect 511960 580740 522396 580768
rect 511960 580728 511966 580740
rect 522390 580728 522396 580740
rect 522448 580728 522454 580780
rect 36538 580660 36544 580712
rect 36596 580700 36602 580712
rect 538398 580700 538404 580712
rect 36596 580672 538404 580700
rect 36596 580660 36602 580672
rect 538398 580660 538404 580672
rect 538456 580660 538462 580712
rect 16298 578892 16304 578944
rect 16356 578932 16362 578944
rect 528646 578932 528652 578944
rect 16356 578904 528652 578932
rect 16356 578892 16362 578904
rect 528646 578892 528652 578904
rect 528704 578892 528710 578944
rect 26050 578484 26056 578536
rect 26108 578524 26114 578536
rect 149698 578524 149704 578536
rect 26108 578496 149704 578524
rect 26108 578484 26114 578496
rect 149698 578484 149704 578496
rect 149756 578484 149762 578536
rect 36722 578416 36728 578468
rect 36780 578456 36786 578468
rect 52454 578456 52460 578468
rect 36780 578428 52460 578456
rect 36780 578416 36786 578428
rect 52454 578416 52460 578428
rect 52512 578416 52518 578468
rect 232314 578416 232320 578468
rect 232372 578456 232378 578468
rect 251818 578456 251824 578468
rect 232372 578428 251824 578456
rect 232372 578416 232378 578428
rect 251818 578416 251824 578428
rect 251876 578416 251882 578468
rect 475378 578416 475384 578468
rect 475436 578456 475442 578468
rect 494698 578456 494704 578468
rect 475436 578428 494704 578456
rect 475436 578416 475442 578428
rect 494698 578416 494704 578428
rect 494756 578416 494762 578468
rect 62482 578348 62488 578400
rect 62540 578388 62546 578400
rect 79318 578388 79324 578400
rect 62540 578360 79324 578388
rect 62540 578348 62546 578360
rect 79318 578348 79324 578360
rect 79376 578348 79382 578400
rect 90450 578348 90456 578400
rect 90508 578388 90514 578400
rect 106458 578388 106464 578400
rect 90508 578360 106464 578388
rect 90508 578348 90514 578360
rect 106458 578348 106464 578360
rect 106516 578348 106522 578400
rect 116486 578348 116492 578400
rect 116544 578388 116550 578400
rect 133414 578388 133420 578400
rect 116544 578360 133420 578388
rect 116544 578348 116550 578360
rect 133414 578348 133420 578360
rect 133472 578348 133478 578400
rect 144178 578348 144184 578400
rect 144236 578388 144242 578400
rect 160278 578388 160284 578400
rect 144236 578360 160284 578388
rect 144236 578348 144242 578360
rect 160278 578348 160284 578360
rect 160336 578348 160342 578400
rect 170490 578348 170496 578400
rect 170548 578388 170554 578400
rect 187786 578388 187792 578400
rect 170548 578360 187792 578388
rect 170548 578348 170554 578360
rect 187786 578348 187792 578360
rect 187844 578348 187850 578400
rect 197538 578348 197544 578400
rect 197596 578388 197602 578400
rect 214374 578388 214380 578400
rect 197596 578360 214380 578388
rect 197596 578348 197602 578360
rect 214374 578348 214380 578360
rect 214432 578348 214438 578400
rect 224494 578348 224500 578400
rect 224552 578388 224558 578400
rect 241606 578388 241612 578400
rect 224552 578360 241612 578388
rect 224552 578348 224558 578360
rect 241606 578348 241612 578360
rect 241664 578348 241670 578400
rect 413462 578348 413468 578400
rect 413520 578388 413526 578400
rect 430574 578388 430580 578400
rect 413520 578360 430580 578388
rect 413520 578348 413526 578360
rect 430574 578348 430580 578360
rect 430632 578348 430638 578400
rect 440510 578348 440516 578400
rect 440568 578388 440574 578400
rect 457254 578388 457260 578400
rect 440568 578360 457260 578388
rect 440568 578348 440574 578360
rect 457254 578348 457260 578360
rect 457312 578348 457318 578400
rect 468478 578348 468484 578400
rect 468536 578388 468542 578400
rect 484394 578388 484400 578400
rect 468536 578360 484400 578388
rect 468536 578348 468542 578360
rect 484394 578348 484400 578360
rect 484452 578348 484458 578400
rect 36814 578280 36820 578332
rect 36872 578320 36878 578332
rect 62114 578320 62120 578332
rect 36872 578292 62120 578320
rect 36872 578280 36878 578292
rect 62114 578280 62120 578292
rect 62172 578280 62178 578332
rect 64138 578280 64144 578332
rect 64196 578320 64202 578332
rect 89070 578320 89076 578332
rect 64196 578292 89076 578320
rect 64196 578280 64202 578292
rect 89070 578280 89076 578292
rect 89128 578280 89134 578332
rect 90358 578280 90364 578332
rect 90416 578320 90422 578332
rect 116118 578320 116124 578332
rect 90416 578292 116124 578320
rect 90416 578280 90422 578292
rect 116118 578280 116124 578292
rect 116176 578280 116182 578332
rect 116578 578280 116584 578332
rect 116636 578320 116642 578332
rect 142982 578320 142988 578332
rect 116636 578292 142988 578320
rect 116636 578280 116642 578292
rect 142982 578280 142988 578292
rect 143040 578280 143046 578332
rect 144270 578280 144276 578332
rect 144328 578320 144334 578332
rect 170030 578320 170036 578332
rect 144328 578292 170036 578320
rect 144328 578280 144334 578292
rect 170030 578280 170036 578292
rect 170088 578280 170094 578332
rect 178402 578280 178408 578332
rect 178460 578320 178466 578332
rect 200758 578320 200764 578332
rect 178460 578292 200764 578320
rect 178460 578280 178466 578292
rect 200758 578280 200764 578292
rect 200816 578280 200822 578332
rect 251450 578280 251456 578332
rect 251508 578320 251514 578332
rect 268286 578320 268292 578332
rect 251508 578292 268292 578320
rect 251508 578280 251514 578292
rect 268286 578280 268292 578292
rect 268344 578280 268350 578332
rect 279418 578280 279424 578332
rect 279476 578320 279482 578332
rect 295794 578320 295800 578332
rect 279476 578292 295800 578320
rect 279476 578280 279482 578292
rect 295794 578280 295800 578292
rect 295852 578280 295858 578332
rect 305546 578280 305552 578332
rect 305604 578320 305610 578332
rect 322382 578320 322388 578332
rect 305604 578292 322388 578320
rect 305604 578280 305610 578292
rect 322382 578280 322388 578292
rect 322440 578280 322446 578332
rect 335998 578280 336004 578332
rect 336056 578320 336062 578332
rect 349798 578320 349804 578332
rect 336056 578292 349804 578320
rect 336056 578280 336062 578292
rect 349798 578280 349804 578292
rect 349856 578280 349862 578332
rect 359642 578280 359648 578332
rect 359700 578320 359706 578332
rect 376294 578320 376300 578332
rect 359700 578292 376300 578320
rect 359700 578280 359706 578292
rect 376294 578280 376300 578292
rect 376352 578280 376358 578332
rect 386506 578280 386512 578332
rect 386564 578320 386570 578332
rect 403342 578320 403348 578332
rect 386564 578292 403348 578320
rect 386564 578280 386570 578292
rect 403342 578280 403348 578292
rect 403400 578280 403406 578332
rect 421282 578280 421288 578332
rect 421340 578320 421346 578332
rect 446398 578320 446404 578332
rect 421340 578292 446404 578320
rect 421340 578280 421346 578292
rect 446398 578280 446404 578292
rect 446456 578280 446462 578332
rect 494514 578280 494520 578332
rect 494572 578320 494578 578332
rect 511350 578320 511356 578332
rect 494572 578292 511356 578320
rect 494572 578280 494578 578292
rect 511350 578280 511356 578292
rect 511408 578280 511414 578332
rect 522390 578280 522396 578332
rect 522448 578320 522454 578332
rect 538398 578320 538404 578332
rect 522448 578292 538404 578320
rect 522448 578280 522454 578292
rect 538398 578280 538404 578292
rect 538456 578280 538462 578332
rect 43346 578212 43352 578264
rect 43404 578252 43410 578264
rect 62758 578252 62764 578264
rect 43404 578224 62764 578252
rect 43404 578212 43410 578224
rect 62758 578212 62764 578224
rect 62816 578212 62822 578264
rect 171778 578212 171784 578264
rect 171836 578252 171842 578264
rect 197446 578252 197452 578264
rect 171836 578224 197452 578252
rect 171836 578212 171842 578224
rect 197446 578212 197452 578224
rect 197504 578212 197510 578264
rect 199378 578212 199384 578264
rect 199436 578252 199442 578264
rect 223942 578252 223948 578264
rect 199436 578224 223948 578252
rect 199436 578212 199442 578224
rect 223942 578212 223948 578224
rect 224000 578212 224006 578264
rect 225598 578212 225604 578264
rect 225656 578252 225662 578264
rect 251266 578252 251272 578264
rect 225656 578224 251272 578252
rect 225656 578212 225662 578224
rect 251266 578212 251272 578224
rect 251324 578212 251330 578264
rect 253198 578212 253204 578264
rect 253256 578252 253262 578264
rect 278038 578252 278044 578264
rect 253256 578224 278044 578252
rect 253256 578212 253262 578224
rect 278038 578212 278044 578224
rect 278096 578212 278102 578264
rect 279510 578212 279516 578264
rect 279568 578252 279574 578264
rect 305454 578252 305460 578264
rect 279568 578224 305460 578252
rect 279568 578212 279574 578224
rect 305454 578212 305460 578224
rect 305512 578212 305518 578264
rect 307018 578212 307024 578264
rect 307076 578252 307082 578264
rect 331950 578252 331956 578264
rect 307076 578224 331956 578252
rect 307076 578212 307082 578224
rect 331950 578212 331956 578224
rect 332008 578212 332014 578264
rect 333238 578212 333244 578264
rect 333296 578252 333302 578264
rect 359458 578252 359464 578264
rect 333296 578224 359464 578252
rect 333296 578212 333302 578224
rect 359458 578212 359464 578224
rect 359516 578212 359522 578264
rect 359734 578212 359740 578264
rect 359792 578252 359798 578264
rect 386046 578252 386052 578264
rect 359792 578224 386052 578252
rect 359792 578212 359798 578224
rect 386046 578212 386052 578224
rect 386104 578212 386110 578264
rect 387058 578212 387064 578264
rect 387116 578252 387122 578264
rect 412910 578252 412916 578264
rect 387116 578224 412916 578252
rect 387116 578212 387122 578224
rect 412910 578212 412916 578224
rect 412968 578212 412974 578264
rect 414658 578212 414664 578264
rect 414716 578252 414722 578264
rect 440234 578252 440240 578264
rect 414716 578224 440240 578252
rect 414716 578212 414722 578224
rect 440234 578212 440240 578224
rect 440292 578212 440298 578264
rect 442258 578212 442264 578264
rect 442316 578252 442322 578264
rect 467006 578252 467012 578264
rect 442316 578224 467012 578252
rect 442316 578212 442322 578224
rect 467006 578212 467012 578224
rect 467064 578212 467070 578264
rect 468570 578212 468576 578264
rect 468628 578252 468634 578264
rect 494054 578252 494060 578264
rect 468628 578224 494060 578252
rect 468628 578212 468634 578224
rect 494054 578212 494060 578224
rect 494112 578212 494118 578264
rect 496078 578212 496084 578264
rect 496136 578252 496142 578264
rect 520918 578252 520924 578264
rect 496136 578224 520924 578252
rect 496136 578212 496142 578224
rect 520918 578212 520924 578224
rect 520976 578212 520982 578264
rect 522298 578212 522304 578264
rect 522356 578252 522362 578264
rect 547966 578252 547972 578264
rect 522356 578224 547972 578252
rect 522356 578212 522362 578224
rect 547966 578212 547972 578224
rect 548024 578212 548030 578264
rect 37918 576104 37924 576156
rect 37976 576144 37982 576156
rect 526438 576144 526444 576156
rect 37976 576116 526444 576144
rect 37976 576104 37982 576116
rect 526438 576104 526444 576116
rect 526496 576104 526502 576156
rect 285766 575356 285772 575408
rect 285824 575396 285830 575408
rect 286134 575396 286140 575408
rect 285824 575368 286140 575396
rect 285824 575356 285830 575368
rect 286134 575356 286140 575368
rect 286192 575356 286198 575408
rect 339586 575288 339592 575340
rect 339644 575328 339650 575340
rect 340138 575328 340144 575340
rect 339644 575300 340144 575328
rect 339644 575288 339650 575300
rect 340138 575288 340144 575300
rect 340196 575288 340202 575340
rect 89714 562300 89720 562352
rect 89772 562340 89778 562352
rect 90450 562340 90456 562352
rect 89772 562312 90456 562340
rect 89772 562300 89778 562312
rect 90450 562300 90456 562312
rect 90508 562300 90514 562352
rect 13722 557472 13728 557524
rect 13780 557512 13786 557524
rect 64874 557512 64880 557524
rect 13780 557484 64880 557512
rect 13780 557472 13786 557484
rect 64874 557472 64880 557484
rect 64932 557472 64938 557524
rect 95142 557472 95148 557524
rect 95200 557512 95206 557524
rect 146294 557512 146300 557524
rect 95200 557484 146300 557512
rect 95200 557472 95206 557484
rect 146294 557472 146300 557484
rect 146352 557472 146358 557524
rect 148962 557472 148968 557524
rect 149020 557512 149026 557524
rect 200114 557512 200120 557524
rect 149020 557484 200120 557512
rect 149020 557472 149026 557484
rect 200114 557472 200120 557484
rect 200172 557472 200178 557524
rect 202782 557472 202788 557524
rect 202840 557512 202846 557524
rect 253934 557512 253940 557524
rect 202840 557484 253940 557512
rect 202840 557472 202846 557484
rect 253934 557472 253940 557484
rect 253992 557472 253998 557524
rect 256602 557472 256608 557524
rect 256660 557512 256666 557524
rect 307754 557512 307760 557524
rect 256660 557484 307760 557512
rect 256660 557472 256666 557484
rect 307754 557472 307760 557484
rect 307812 557472 307818 557524
rect 338022 557472 338028 557524
rect 338080 557512 338086 557524
rect 389174 557512 389180 557524
rect 338080 557484 389180 557512
rect 338080 557472 338086 557484
rect 389174 557472 389180 557484
rect 389232 557472 389238 557524
rect 391842 557472 391848 557524
rect 391900 557512 391906 557524
rect 442994 557512 443000 557524
rect 391900 557484 443000 557512
rect 391900 557472 391906 557484
rect 442994 557472 443000 557484
rect 443052 557472 443058 557524
rect 445662 557472 445668 557524
rect 445720 557512 445726 557524
rect 496814 557512 496820 557524
rect 445720 557484 496820 557512
rect 445720 557472 445726 557484
rect 496814 557472 496820 557484
rect 496872 557472 496878 557524
rect 500862 557472 500868 557524
rect 500920 557512 500926 557524
rect 550634 557512 550640 557524
rect 500920 557484 550640 557512
rect 500920 557472 500926 557484
rect 550634 557472 550640 557484
rect 550692 557472 550698 557524
rect 35618 557404 35624 557456
rect 35676 557444 35682 557456
rect 36722 557444 36728 557456
rect 35676 557416 36728 557444
rect 35676 557404 35682 557416
rect 36722 557404 36728 557416
rect 36780 557404 36786 557456
rect 41322 557404 41328 557456
rect 41380 557444 41386 557456
rect 91094 557444 91100 557456
rect 41380 557416 91100 557444
rect 41380 557404 41386 557416
rect 91094 557404 91100 557416
rect 91152 557404 91158 557456
rect 122742 557404 122748 557456
rect 122800 557444 122806 557456
rect 172514 557444 172520 557456
rect 122800 557416 172520 557444
rect 122800 557404 122806 557416
rect 172514 557404 172520 557416
rect 172572 557404 172578 557456
rect 176562 557404 176568 557456
rect 176620 557444 176626 557456
rect 226334 557444 226340 557456
rect 176620 557416 226340 557444
rect 176620 557404 176626 557416
rect 226334 557404 226340 557416
rect 226392 557404 226398 557456
rect 230382 557404 230388 557456
rect 230440 557444 230446 557456
rect 280154 557444 280160 557456
rect 230440 557416 280160 557444
rect 230440 557404 230446 557416
rect 280154 557404 280160 557416
rect 280212 557404 280218 557456
rect 284202 557404 284208 557456
rect 284260 557444 284266 557456
rect 335354 557444 335360 557456
rect 284260 557416 335360 557444
rect 284260 557404 284266 557416
rect 335354 557404 335360 557416
rect 335412 557404 335418 557456
rect 365622 557404 365628 557456
rect 365680 557444 365686 557456
rect 415394 557444 415400 557456
rect 365680 557416 415400 557444
rect 365680 557404 365686 557416
rect 415394 557404 415400 557416
rect 415452 557404 415458 557456
rect 419442 557404 419448 557456
rect 419500 557444 419506 557456
rect 469214 557444 469220 557456
rect 419500 557416 444374 557444
rect 419500 557404 419506 557416
rect 68922 557336 68928 557388
rect 68980 557376 68986 557388
rect 118694 557376 118700 557388
rect 68980 557348 118700 557376
rect 68980 557336 68986 557348
rect 118694 557336 118700 557348
rect 118752 557336 118758 557388
rect 311802 557336 311808 557388
rect 311860 557376 311866 557388
rect 361574 557376 361580 557388
rect 311860 557348 361580 557376
rect 311860 557336 311866 557348
rect 361574 557336 361580 557348
rect 361632 557336 361638 557388
rect 444346 557308 444374 557416
rect 454006 557416 469220 557444
rect 454006 557308 454034 557416
rect 469214 557404 469220 557416
rect 469272 557404 469278 557456
rect 473262 557404 473268 557456
rect 473320 557444 473326 557456
rect 523034 557444 523040 557456
rect 473320 557416 523040 557444
rect 473320 557404 473326 557416
rect 523034 557404 523040 557416
rect 523092 557404 523098 557456
rect 444346 557280 454034 557308
rect 446398 556724 446404 556776
rect 446456 556764 446462 556776
rect 447686 556764 447692 556776
rect 446456 556736 447692 556764
rect 446456 556724 446462 556736
rect 447686 556724 447692 556736
rect 447744 556724 447750 556776
rect 521746 556724 521752 556776
rect 521804 556764 521810 556776
rect 522390 556764 522396 556776
rect 521804 556736 522396 556764
rect 521804 556724 521810 556736
rect 522390 556724 522396 556736
rect 522448 556724 522454 556776
rect 52730 554684 52736 554736
rect 52788 554724 52794 554736
rect 64138 554724 64144 554736
rect 52788 554696 64144 554724
rect 52788 554684 52794 554696
rect 64138 554684 64144 554696
rect 64196 554684 64202 554736
rect 69106 554684 69112 554736
rect 69164 554724 69170 554736
rect 69164 554696 74534 554724
rect 69164 554684 69170 554696
rect 15194 554616 15200 554668
rect 15252 554656 15258 554668
rect 42978 554656 42984 554668
rect 15252 554628 42984 554656
rect 15252 554616 15258 554628
rect 42978 554616 42984 554628
rect 43036 554616 43042 554668
rect 62758 554616 62764 554668
rect 62816 554656 62822 554668
rect 70026 554656 70032 554668
rect 62816 554628 70032 554656
rect 62816 554616 62822 554628
rect 70026 554616 70032 554628
rect 70084 554616 70090 554668
rect 74506 554656 74534 554696
rect 96706 554684 96712 554736
rect 96764 554724 96770 554736
rect 96764 554696 103514 554724
rect 96764 554684 96770 554696
rect 96982 554656 96988 554668
rect 74506 554628 96988 554656
rect 96982 554616 96988 554628
rect 97040 554616 97046 554668
rect 103486 554656 103514 554696
rect 146938 554684 146944 554736
rect 146996 554724 147002 554736
rect 146996 554696 151814 554724
rect 146996 554684 147002 554696
rect 124030 554656 124036 554668
rect 103486 554628 124036 554656
rect 124030 554616 124036 554628
rect 124088 554616 124094 554668
rect 133690 554616 133696 554668
rect 133748 554656 133754 554668
rect 144270 554656 144276 554668
rect 133748 554628 144276 554656
rect 133748 554616 133754 554628
rect 144270 554616 144276 554628
rect 144328 554616 144334 554668
rect 150526 554616 150532 554668
rect 150584 554656 150590 554668
rect 151786 554656 151814 554696
rect 200758 554684 200764 554736
rect 200816 554724 200822 554736
rect 204990 554724 204996 554736
rect 200816 554696 204996 554724
rect 200816 554684 200822 554696
rect 204990 554684 204996 554696
rect 205048 554684 205054 554736
rect 251818 554684 251824 554736
rect 251876 554724 251882 554736
rect 258994 554724 259000 554736
rect 251876 554696 259000 554724
rect 251876 554684 251882 554696
rect 258994 554684 259000 554696
rect 259052 554684 259058 554736
rect 332318 554684 332324 554736
rect 332376 554724 332382 554736
rect 335998 554724 336004 554736
rect 332376 554696 336004 554724
rect 332376 554684 332382 554696
rect 335998 554684 336004 554696
rect 336056 554684 336062 554736
rect 494698 554684 494704 554736
rect 494756 554724 494762 554736
rect 501966 554724 501972 554736
rect 494756 554696 501972 554724
rect 494756 554684 494762 554696
rect 501966 554684 501972 554696
rect 502024 554684 502030 554736
rect 548334 554656 548340 554668
rect 150584 554628 151124 554656
rect 151786 554628 548340 554656
rect 150584 554616 150590 554628
rect 25682 554548 25688 554600
rect 25740 554588 25746 554600
rect 36814 554588 36820 554600
rect 25740 554560 36820 554588
rect 25740 554548 25746 554560
rect 36814 554548 36820 554560
rect 36872 554548 36878 554600
rect 79686 554548 79692 554600
rect 79744 554588 79750 554600
rect 90358 554588 90364 554600
rect 79744 554560 90364 554588
rect 79744 554548 79750 554560
rect 90358 554548 90364 554560
rect 90416 554548 90422 554600
rect 106642 554548 106648 554600
rect 106700 554588 106706 554600
rect 116578 554588 116584 554600
rect 106700 554560 116584 554588
rect 106700 554548 106706 554560
rect 116578 554548 116584 554560
rect 116636 554548 116642 554600
rect 122926 554548 122932 554600
rect 122984 554588 122990 554600
rect 150986 554588 150992 554600
rect 122984 554560 150992 554588
rect 122984 554548 122990 554560
rect 150986 554548 150992 554560
rect 151044 554548 151050 554600
rect 151096 554588 151124 554628
rect 548334 554616 548340 554628
rect 548392 554616 548398 554668
rect 178034 554588 178040 554600
rect 151096 554560 178040 554588
rect 178034 554548 178040 554560
rect 178092 554548 178098 554600
rect 187694 554548 187700 554600
rect 187752 554588 187758 554600
rect 199378 554588 199384 554600
rect 187752 554560 199384 554588
rect 187752 554548 187758 554560
rect 199378 554548 199384 554560
rect 199436 554548 199442 554600
rect 204346 554548 204352 554600
rect 204404 554588 204410 554600
rect 232038 554588 232044 554600
rect 204404 554560 232044 554588
rect 204404 554548 204410 554560
rect 232038 554548 232044 554560
rect 232096 554548 232102 554600
rect 241698 554548 241704 554600
rect 241756 554588 241762 554600
rect 253198 554588 253204 554600
rect 241756 554560 253204 554588
rect 241756 554548 241762 554560
rect 253198 554548 253204 554560
rect 253256 554548 253262 554600
rect 258166 554548 258172 554600
rect 258224 554588 258230 554600
rect 286042 554588 286048 554600
rect 258224 554560 286048 554588
rect 258224 554548 258230 554560
rect 286042 554548 286048 554560
rect 286100 554548 286106 554600
rect 312998 554588 313004 554600
rect 287026 554560 313004 554588
rect 160646 554480 160652 554532
rect 160704 554520 160710 554532
rect 171778 554520 171784 554532
rect 160704 554492 171784 554520
rect 160704 554480 160710 554492
rect 171778 554480 171784 554492
rect 171836 554480 171842 554532
rect 214650 554480 214656 554532
rect 214708 554520 214714 554532
rect 225598 554520 225604 554532
rect 214708 554492 225604 554520
rect 214708 554480 214714 554492
rect 225598 554480 225604 554492
rect 225656 554480 225662 554532
rect 268654 554480 268660 554532
rect 268712 554520 268718 554532
rect 279510 554520 279516 554532
rect 268712 554492 279516 554520
rect 268712 554480 268718 554492
rect 279510 554480 279516 554492
rect 279568 554480 279574 554532
rect 285766 554480 285772 554532
rect 285824 554520 285830 554532
rect 287026 554520 287054 554560
rect 312998 554548 313004 554560
rect 313056 554548 313062 554600
rect 340046 554588 340052 554600
rect 316006 554560 340052 554588
rect 285824 554492 287054 554520
rect 285824 554480 285830 554492
rect 295702 554480 295708 554532
rect 295760 554520 295766 554532
rect 307018 554520 307024 554532
rect 295760 554492 307024 554520
rect 295760 554480 295766 554492
rect 307018 554480 307024 554492
rect 307076 554480 307082 554532
rect 311986 554480 311992 554532
rect 312044 554520 312050 554532
rect 316006 554520 316034 554560
rect 340046 554548 340052 554560
rect 340104 554548 340110 554600
rect 367002 554588 367008 554600
rect 344986 554560 367008 554588
rect 312044 554492 316034 554520
rect 312044 554480 312050 554492
rect 322658 554480 322664 554532
rect 322716 554520 322722 554532
rect 333238 554520 333244 554532
rect 322716 554492 333244 554520
rect 322716 554480 322722 554492
rect 333238 554480 333244 554492
rect 333296 554480 333302 554532
rect 339586 554480 339592 554532
rect 339644 554520 339650 554532
rect 344986 554520 345014 554560
rect 367002 554548 367008 554560
rect 367060 554548 367066 554600
rect 393958 554588 393964 554600
rect 373966 554560 393964 554588
rect 339644 554492 345014 554520
rect 339644 554480 339650 554492
rect 349706 554480 349712 554532
rect 349764 554520 349770 554532
rect 359550 554520 359556 554532
rect 349764 554492 359556 554520
rect 349764 554480 349770 554492
rect 359550 554480 359556 554492
rect 359608 554480 359614 554532
rect 365806 554480 365812 554532
rect 365864 554520 365870 554532
rect 373966 554520 373994 554560
rect 393958 554548 393964 554560
rect 394016 554548 394022 554600
rect 421006 554588 421012 554600
rect 402946 554560 421012 554588
rect 365864 554492 373994 554520
rect 365864 554480 365870 554492
rect 376662 554480 376668 554532
rect 376720 554520 376726 554532
rect 387058 554520 387064 554532
rect 376720 554492 387064 554520
rect 376720 554480 376726 554492
rect 387058 554480 387064 554492
rect 387116 554480 387122 554532
rect 393406 554480 393412 554532
rect 393464 554520 393470 554532
rect 402946 554520 402974 554560
rect 421006 554548 421012 554560
rect 421064 554548 421070 554600
rect 430666 554548 430672 554600
rect 430724 554588 430730 554600
rect 442258 554588 442264 554600
rect 430724 554560 442264 554588
rect 430724 554548 430730 554560
rect 442258 554548 442264 554560
rect 442316 554548 442322 554600
rect 447226 554548 447232 554600
rect 447284 554588 447290 554600
rect 475010 554588 475016 554600
rect 447284 554560 475016 554588
rect 447284 554548 447290 554560
rect 475010 554548 475016 554560
rect 475068 554548 475074 554600
rect 484670 554548 484676 554600
rect 484728 554588 484734 554600
rect 496078 554588 496084 554600
rect 484728 554560 496084 554588
rect 484728 554548 484734 554560
rect 496078 554548 496084 554560
rect 496136 554548 496142 554600
rect 501046 554548 501052 554600
rect 501104 554588 501110 554600
rect 529014 554588 529020 554600
rect 501104 554560 529020 554588
rect 501104 554548 501110 554560
rect 529014 554548 529020 554560
rect 529072 554548 529078 554600
rect 393464 554492 402974 554520
rect 393464 554480 393470 554492
rect 403710 554480 403716 554532
rect 403768 554520 403774 554532
rect 414658 554520 414664 554532
rect 403768 554492 414664 554520
rect 403768 554480 403774 554492
rect 414658 554480 414664 554492
rect 414716 554480 414722 554532
rect 457714 554480 457720 554532
rect 457772 554520 457778 554532
rect 468570 554520 468576 554532
rect 457772 554492 468576 554520
rect 457772 554480 457778 554492
rect 468570 554480 468576 554492
rect 468628 554480 468634 554532
rect 511718 554480 511724 554532
rect 511776 554520 511782 554532
rect 522298 554520 522304 554532
rect 511776 554492 522304 554520
rect 511776 554480 511782 554492
rect 522298 554480 522304 554492
rect 522356 554480 522362 554532
rect 36630 554412 36636 554464
rect 36688 554452 36694 554464
rect 538674 554452 538680 554464
rect 36688 554424 538680 554452
rect 36688 554412 36694 554424
rect 538674 554412 538680 554424
rect 538732 554412 538738 554464
rect 16022 551284 16028 551336
rect 16080 551324 16086 551336
rect 529014 551324 529020 551336
rect 16080 551296 529020 551324
rect 16080 551284 16086 551296
rect 529014 551284 529020 551296
rect 529072 551284 529078 551336
rect 25682 550876 25688 550928
rect 25740 550916 25746 550928
rect 146938 550916 146944 550928
rect 25740 550888 146944 550916
rect 25740 550876 25746 550888
rect 146938 550876 146944 550888
rect 146996 550876 147002 550928
rect 36630 550808 36636 550860
rect 36688 550848 36694 550860
rect 52638 550848 52644 550860
rect 36688 550820 52644 550848
rect 36688 550808 36694 550820
rect 52638 550808 52644 550820
rect 52696 550808 52702 550860
rect 232038 550808 232044 550860
rect 232096 550848 232102 550860
rect 251818 550848 251824 550860
rect 232096 550820 251824 550848
rect 232096 550808 232102 550820
rect 251818 550808 251824 550820
rect 251876 550808 251882 550860
rect 475010 550808 475016 550860
rect 475068 550848 475074 550860
rect 494698 550848 494704 550860
rect 475068 550820 494704 550848
rect 475068 550808 475074 550820
rect 494698 550808 494704 550820
rect 494756 550808 494762 550860
rect 62482 550740 62488 550792
rect 62540 550780 62546 550792
rect 79686 550780 79692 550792
rect 62540 550752 79692 550780
rect 62540 550740 62546 550752
rect 79686 550740 79692 550752
rect 79744 550740 79750 550792
rect 90450 550740 90456 550792
rect 90508 550780 90514 550792
rect 106642 550780 106648 550792
rect 90508 550752 106648 550780
rect 90508 550740 90514 550752
rect 106642 550740 106648 550752
rect 106700 550740 106706 550792
rect 116486 550740 116492 550792
rect 116544 550780 116550 550792
rect 133690 550780 133696 550792
rect 116544 550752 133696 550780
rect 116544 550740 116550 550752
rect 133690 550740 133696 550752
rect 133748 550740 133754 550792
rect 170490 550740 170496 550792
rect 170548 550780 170554 550792
rect 187694 550780 187700 550792
rect 170548 550752 187700 550780
rect 170548 550740 170554 550752
rect 187694 550740 187700 550752
rect 187752 550740 187758 550792
rect 197446 550740 197452 550792
rect 197504 550780 197510 550792
rect 214650 550780 214656 550792
rect 197504 550752 214656 550780
rect 197504 550740 197510 550752
rect 214650 550740 214656 550752
rect 214708 550740 214714 550792
rect 224494 550740 224500 550792
rect 224552 550780 224558 550792
rect 241698 550780 241704 550792
rect 224552 550752 241704 550780
rect 224552 550740 224558 550752
rect 241698 550740 241704 550752
rect 241756 550740 241762 550792
rect 413462 550740 413468 550792
rect 413520 550780 413526 550792
rect 430666 550780 430672 550792
rect 413520 550752 430672 550780
rect 413520 550740 413526 550752
rect 430666 550740 430672 550752
rect 430724 550740 430730 550792
rect 440510 550740 440516 550792
rect 440568 550780 440574 550792
rect 457622 550780 457628 550792
rect 440568 550752 457628 550780
rect 440568 550740 440574 550752
rect 457622 550740 457628 550752
rect 457680 550740 457686 550792
rect 468478 550740 468484 550792
rect 468536 550780 468542 550792
rect 484670 550780 484676 550792
rect 468536 550752 484676 550780
rect 468536 550740 468542 550752
rect 484670 550740 484676 550752
rect 484728 550740 484734 550792
rect 36814 550672 36820 550724
rect 36872 550712 36878 550724
rect 62298 550712 62304 550724
rect 36872 550684 62304 550712
rect 36872 550672 36878 550684
rect 62298 550672 62304 550684
rect 62356 550672 62362 550724
rect 64138 550672 64144 550724
rect 64196 550712 64202 550724
rect 89346 550712 89352 550724
rect 64196 550684 89352 550712
rect 64196 550672 64202 550684
rect 89346 550672 89352 550684
rect 89404 550672 89410 550724
rect 90358 550672 90364 550724
rect 90416 550712 90422 550724
rect 116302 550712 116308 550724
rect 90416 550684 116308 550712
rect 90416 550672 90422 550684
rect 116302 550672 116308 550684
rect 116360 550672 116366 550724
rect 116578 550672 116584 550724
rect 116636 550712 116642 550724
rect 143350 550712 143356 550724
rect 116636 550684 143356 550712
rect 116636 550672 116642 550684
rect 143350 550672 143356 550684
rect 143408 550672 143414 550724
rect 144270 550672 144276 550724
rect 144328 550712 144334 550724
rect 170306 550712 170312 550724
rect 144328 550684 170312 550712
rect 144328 550672 144334 550684
rect 170306 550672 170312 550684
rect 170364 550672 170370 550724
rect 178034 550672 178040 550724
rect 178092 550712 178098 550724
rect 200758 550712 200764 550724
rect 178092 550684 200764 550712
rect 178092 550672 178098 550684
rect 200758 550672 200764 550684
rect 200816 550672 200822 550724
rect 251450 550672 251456 550724
rect 251508 550712 251514 550724
rect 268654 550712 268660 550724
rect 251508 550684 268660 550712
rect 251508 550672 251514 550684
rect 268654 550672 268660 550684
rect 268712 550672 268718 550724
rect 279510 550672 279516 550724
rect 279568 550712 279574 550724
rect 295702 550712 295708 550724
rect 279568 550684 295708 550712
rect 279568 550672 279574 550684
rect 295702 550672 295708 550684
rect 295760 550672 295766 550724
rect 305454 550672 305460 550724
rect 305512 550712 305518 550724
rect 322658 550712 322664 550724
rect 305512 550684 322664 550712
rect 305512 550672 305518 550684
rect 322658 550672 322664 550684
rect 322716 550672 322722 550724
rect 334618 550672 334624 550724
rect 334676 550712 334682 550724
rect 349706 550712 349712 550724
rect 334676 550684 349712 550712
rect 334676 550672 334682 550684
rect 349706 550672 349712 550684
rect 349764 550672 349770 550724
rect 359458 550672 359464 550724
rect 359516 550712 359522 550724
rect 376662 550712 376668 550724
rect 359516 550684 376668 550712
rect 359516 550672 359522 550684
rect 376662 550672 376668 550684
rect 376720 550672 376726 550724
rect 386506 550672 386512 550724
rect 386564 550712 386570 550724
rect 403618 550712 403624 550724
rect 386564 550684 403624 550712
rect 386564 550672 386570 550684
rect 403618 550672 403624 550684
rect 403676 550672 403682 550724
rect 421006 550672 421012 550724
rect 421064 550712 421070 550724
rect 443638 550712 443644 550724
rect 421064 550684 443644 550712
rect 421064 550672 421070 550684
rect 443638 550672 443644 550684
rect 443696 550672 443702 550724
rect 494514 550672 494520 550724
rect 494572 550712 494578 550724
rect 511626 550712 511632 550724
rect 494572 550684 511632 550712
rect 494572 550672 494578 550684
rect 511626 550672 511632 550684
rect 511684 550672 511690 550724
rect 522298 550672 522304 550724
rect 522356 550712 522362 550724
rect 538674 550712 538680 550724
rect 522356 550684 538680 550712
rect 522356 550672 522362 550684
rect 538674 550672 538680 550684
rect 538732 550672 538738 550724
rect 43070 550604 43076 550656
rect 43128 550644 43134 550656
rect 62758 550644 62764 550656
rect 43128 550616 62764 550644
rect 43128 550604 43134 550616
rect 62758 550604 62764 550616
rect 62816 550604 62822 550656
rect 144178 550604 144184 550656
rect 144236 550644 144242 550656
rect 160646 550644 160652 550656
rect 144236 550616 160652 550644
rect 144236 550604 144242 550616
rect 160646 550604 160652 550616
rect 160704 550604 160710 550656
rect 171778 550604 171784 550656
rect 171836 550644 171842 550656
rect 197354 550644 197360 550656
rect 171836 550616 197360 550644
rect 171836 550604 171842 550616
rect 197354 550604 197360 550616
rect 197412 550604 197418 550656
rect 199378 550604 199384 550656
rect 199436 550644 199442 550656
rect 224310 550644 224316 550656
rect 199436 550616 224316 550644
rect 199436 550604 199442 550616
rect 224310 550604 224316 550616
rect 224368 550604 224374 550656
rect 225598 550604 225604 550656
rect 225656 550644 225662 550656
rect 251358 550644 251364 550656
rect 225656 550616 251364 550644
rect 225656 550604 225662 550616
rect 251358 550604 251364 550616
rect 251416 550604 251422 550656
rect 253198 550604 253204 550656
rect 253256 550644 253262 550656
rect 278314 550644 278320 550656
rect 253256 550616 278320 550644
rect 253256 550604 253262 550616
rect 278314 550604 278320 550616
rect 278372 550604 278378 550656
rect 279418 550604 279424 550656
rect 279476 550644 279482 550656
rect 305362 550644 305368 550656
rect 279476 550616 305368 550644
rect 279476 550604 279482 550616
rect 305362 550604 305368 550616
rect 305420 550604 305426 550656
rect 307018 550604 307024 550656
rect 307076 550644 307082 550656
rect 332318 550644 332324 550656
rect 307076 550616 332324 550644
rect 307076 550604 307082 550616
rect 332318 550604 332324 550616
rect 332376 550604 332382 550656
rect 333238 550604 333244 550656
rect 333296 550644 333302 550656
rect 359366 550644 359372 550656
rect 333296 550616 359372 550644
rect 333296 550604 333302 550616
rect 359366 550604 359372 550616
rect 359424 550604 359430 550656
rect 359550 550604 359556 550656
rect 359608 550644 359614 550656
rect 386322 550644 386328 550656
rect 359608 550616 386328 550644
rect 359608 550604 359614 550616
rect 386322 550604 386328 550616
rect 386380 550604 386386 550656
rect 387058 550604 387064 550656
rect 387116 550644 387122 550656
rect 413278 550644 413284 550656
rect 387116 550616 413284 550644
rect 387116 550604 387122 550616
rect 413278 550604 413284 550616
rect 413336 550604 413342 550656
rect 414658 550604 414664 550656
rect 414716 550644 414722 550656
rect 440326 550644 440332 550656
rect 414716 550616 440332 550644
rect 414716 550604 414722 550616
rect 440326 550604 440332 550616
rect 440384 550604 440390 550656
rect 442258 550604 442264 550656
rect 442316 550644 442322 550656
rect 467282 550644 467288 550656
rect 442316 550616 467288 550644
rect 442316 550604 442322 550616
rect 467282 550604 467288 550616
rect 467340 550604 467346 550656
rect 468570 550604 468576 550656
rect 468628 550644 468634 550656
rect 494330 550644 494336 550656
rect 468628 550616 494336 550644
rect 468628 550604 468634 550616
rect 494330 550604 494336 550616
rect 494388 550604 494394 550656
rect 496078 550604 496084 550656
rect 496136 550644 496142 550656
rect 521286 550644 521292 550656
rect 496136 550616 521292 550644
rect 496136 550604 496142 550616
rect 521286 550604 521292 550616
rect 521344 550604 521350 550656
rect 522390 550604 522396 550656
rect 522448 550644 522454 550656
rect 548334 550644 548340 550656
rect 522448 550616 548340 550644
rect 522448 550604 522454 550616
rect 548334 550604 548340 550616
rect 548392 550604 548398 550656
rect 37918 548496 37924 548548
rect 37976 548536 37982 548548
rect 526438 548536 526444 548548
rect 37976 548508 526444 548536
rect 37976 548496 37982 548508
rect 526438 548496 526444 548508
rect 526496 548496 526502 548548
rect 35618 547884 35624 547936
rect 35676 547924 35682 547936
rect 36722 547924 36728 547936
rect 35676 547896 36728 547924
rect 35676 547884 35682 547896
rect 36722 547884 36728 547896
rect 36780 547884 36786 547936
rect 89714 533604 89720 533656
rect 89772 533644 89778 533656
rect 90450 533644 90456 533656
rect 89772 533616 90456 533644
rect 89772 533604 89778 533616
rect 90450 533604 90456 533616
rect 90508 533604 90514 533656
rect 13722 529864 13728 529916
rect 13780 529904 13786 529916
rect 64874 529904 64880 529916
rect 13780 529876 64880 529904
rect 13780 529864 13786 529876
rect 64874 529864 64880 529876
rect 64932 529864 64938 529916
rect 95142 529864 95148 529916
rect 95200 529904 95206 529916
rect 146294 529904 146300 529916
rect 95200 529876 146300 529904
rect 95200 529864 95206 529876
rect 146294 529864 146300 529876
rect 146352 529864 146358 529916
rect 148962 529864 148968 529916
rect 149020 529904 149026 529916
rect 200114 529904 200120 529916
rect 149020 529876 200120 529904
rect 149020 529864 149026 529876
rect 200114 529864 200120 529876
rect 200172 529864 200178 529916
rect 202782 529864 202788 529916
rect 202840 529904 202846 529916
rect 253934 529904 253940 529916
rect 202840 529876 253940 529904
rect 202840 529864 202846 529876
rect 253934 529864 253940 529876
rect 253992 529864 253998 529916
rect 256602 529864 256608 529916
rect 256660 529904 256666 529916
rect 307754 529904 307760 529916
rect 256660 529876 307760 529904
rect 256660 529864 256666 529876
rect 307754 529864 307760 529876
rect 307812 529864 307818 529916
rect 332502 529864 332508 529916
rect 332560 529904 332566 529916
rect 334618 529904 334624 529916
rect 332560 529876 334624 529904
rect 332560 529864 332566 529876
rect 334618 529864 334624 529876
rect 334676 529864 334682 529916
rect 338022 529864 338028 529916
rect 338080 529904 338086 529916
rect 389174 529904 389180 529916
rect 338080 529876 389180 529904
rect 338080 529864 338086 529876
rect 389174 529864 389180 529876
rect 389232 529864 389238 529916
rect 391842 529864 391848 529916
rect 391900 529904 391906 529916
rect 442994 529904 443000 529916
rect 391900 529876 443000 529904
rect 391900 529864 391906 529876
rect 442994 529864 443000 529876
rect 443052 529864 443058 529916
rect 445662 529864 445668 529916
rect 445720 529904 445726 529916
rect 496814 529904 496820 529916
rect 445720 529876 496820 529904
rect 445720 529864 445726 529876
rect 496814 529864 496820 529876
rect 496872 529864 496878 529916
rect 500862 529864 500868 529916
rect 500920 529904 500926 529916
rect 550634 529904 550640 529916
rect 500920 529876 550640 529904
rect 500920 529864 500926 529876
rect 550634 529864 550640 529876
rect 550692 529864 550698 529916
rect 35618 529796 35624 529848
rect 35676 529836 35682 529848
rect 36630 529836 36636 529848
rect 35676 529808 36636 529836
rect 35676 529796 35682 529808
rect 36630 529796 36636 529808
rect 36688 529796 36694 529848
rect 41322 529796 41328 529848
rect 41380 529836 41386 529848
rect 91094 529836 91100 529848
rect 41380 529808 91100 529836
rect 41380 529796 41386 529808
rect 91094 529796 91100 529808
rect 91152 529796 91158 529848
rect 122742 529796 122748 529848
rect 122800 529836 122806 529848
rect 172514 529836 172520 529848
rect 122800 529808 172520 529836
rect 122800 529796 122806 529808
rect 172514 529796 172520 529808
rect 172572 529796 172578 529848
rect 176562 529796 176568 529848
rect 176620 529836 176626 529848
rect 226334 529836 226340 529848
rect 176620 529808 226340 529836
rect 176620 529796 176626 529808
rect 226334 529796 226340 529808
rect 226392 529796 226398 529848
rect 230382 529796 230388 529848
rect 230440 529836 230446 529848
rect 230440 529808 277394 529836
rect 230440 529796 230446 529808
rect 68922 529728 68928 529780
rect 68980 529768 68986 529780
rect 118694 529768 118700 529780
rect 68980 529740 118700 529768
rect 68980 529728 68986 529740
rect 118694 529728 118700 529740
rect 118752 529728 118758 529780
rect 277366 529768 277394 529808
rect 278682 529796 278688 529848
rect 278740 529836 278746 529848
rect 279510 529836 279516 529848
rect 278740 529808 279516 529836
rect 278740 529796 278746 529808
rect 279510 529796 279516 529808
rect 279568 529796 279574 529848
rect 284202 529796 284208 529848
rect 284260 529836 284266 529848
rect 335354 529836 335360 529848
rect 284260 529808 335360 529836
rect 284260 529796 284266 529808
rect 335354 529796 335360 529808
rect 335412 529796 335418 529848
rect 365622 529796 365628 529848
rect 365680 529836 365686 529848
rect 415394 529836 415400 529848
rect 365680 529808 415400 529836
rect 365680 529796 365686 529808
rect 415394 529796 415400 529808
rect 415452 529796 415458 529848
rect 419442 529796 419448 529848
rect 419500 529836 419506 529848
rect 469214 529836 469220 529848
rect 419500 529808 469220 529836
rect 419500 529796 419506 529808
rect 469214 529796 469220 529808
rect 469272 529796 469278 529848
rect 473262 529796 473268 529848
rect 473320 529836 473326 529848
rect 523034 529836 523040 529848
rect 473320 529808 523040 529836
rect 473320 529796 473326 529808
rect 523034 529796 523040 529808
rect 523092 529796 523098 529848
rect 280154 529768 280160 529780
rect 277366 529740 280160 529768
rect 280154 529728 280160 529740
rect 280212 529728 280218 529780
rect 311802 529728 311808 529780
rect 311860 529768 311866 529780
rect 361574 529768 361580 529780
rect 311860 529740 361580 529768
rect 311860 529728 311866 529740
rect 361574 529728 361580 529740
rect 361632 529728 361638 529780
rect 116210 529592 116216 529644
rect 116268 529632 116274 529644
rect 116486 529632 116492 529644
rect 116268 529604 116492 529632
rect 116268 529592 116274 529604
rect 116486 529592 116492 529604
rect 116544 529592 116550 529644
rect 170214 529592 170220 529644
rect 170272 529632 170278 529644
rect 170490 529632 170496 529644
rect 170272 529604 170496 529632
rect 170272 529592 170278 529604
rect 170490 529592 170496 529604
rect 170548 529592 170554 529644
rect 53098 527076 53104 527128
rect 53156 527116 53162 527128
rect 64138 527116 64144 527128
rect 53156 527088 64144 527116
rect 53156 527076 53162 527088
rect 64138 527076 64144 527088
rect 64196 527076 64202 527128
rect 69106 527076 69112 527128
rect 69164 527116 69170 527128
rect 69164 527088 74534 527116
rect 69164 527076 69170 527088
rect 15194 527008 15200 527060
rect 15252 527048 15258 527060
rect 42794 527048 42800 527060
rect 15252 527020 42800 527048
rect 15252 527008 15258 527020
rect 42794 527008 42800 527020
rect 42852 527008 42858 527060
rect 62758 527008 62764 527060
rect 62816 527048 62822 527060
rect 69750 527048 69756 527060
rect 62816 527020 69756 527048
rect 62816 527008 62822 527020
rect 69750 527008 69756 527020
rect 69808 527008 69814 527060
rect 74506 527048 74534 527088
rect 96706 527076 96712 527128
rect 96764 527116 96770 527128
rect 96764 527088 103514 527116
rect 96764 527076 96770 527088
rect 96798 527048 96804 527060
rect 74506 527020 96804 527048
rect 96798 527008 96804 527020
rect 96856 527008 96862 527060
rect 103486 527048 103514 527088
rect 200758 527076 200764 527128
rect 200816 527116 200822 527128
rect 204622 527116 204628 527128
rect 200816 527088 204628 527116
rect 200816 527076 200822 527088
rect 204622 527076 204628 527088
rect 204680 527076 204686 527128
rect 251818 527076 251824 527128
rect 251876 527116 251882 527128
rect 258718 527116 258724 527128
rect 251876 527088 258724 527116
rect 251876 527076 251882 527088
rect 258718 527076 258724 527088
rect 258776 527076 258782 527128
rect 443638 527076 443644 527128
rect 443696 527116 443702 527128
rect 447686 527116 447692 527128
rect 443696 527088 447692 527116
rect 443696 527076 443702 527088
rect 447686 527076 447692 527088
rect 447744 527076 447750 527128
rect 494698 527076 494704 527128
rect 494756 527116 494762 527128
rect 501598 527116 501604 527128
rect 494756 527088 501604 527116
rect 494756 527076 494762 527088
rect 501598 527076 501604 527088
rect 501656 527076 501662 527128
rect 123662 527048 123668 527060
rect 103486 527020 123668 527048
rect 123662 527008 123668 527020
rect 123720 527008 123726 527060
rect 149698 527008 149704 527060
rect 149756 527048 149762 527060
rect 547966 527048 547972 527060
rect 149756 527020 547972 527048
rect 149756 527008 149762 527020
rect 547966 527008 547972 527020
rect 548024 527008 548030 527060
rect 26050 526940 26056 526992
rect 26108 526980 26114 526992
rect 36814 526980 36820 526992
rect 26108 526952 36820 526980
rect 26108 526940 26114 526952
rect 36814 526940 36820 526952
rect 36872 526940 36878 526992
rect 79962 526940 79968 526992
rect 80020 526980 80026 526992
rect 90358 526980 90364 526992
rect 80020 526952 90364 526980
rect 80020 526940 80026 526952
rect 90358 526940 90364 526952
rect 90416 526940 90422 526992
rect 106550 526940 106556 526992
rect 106608 526980 106614 526992
rect 116578 526980 116584 526992
rect 106608 526952 116584 526980
rect 106608 526940 106614 526952
rect 116578 526940 116584 526952
rect 116636 526940 116642 526992
rect 133782 526940 133788 526992
rect 133840 526980 133846 526992
rect 144270 526980 144276 526992
rect 133840 526952 144276 526980
rect 133840 526940 133846 526952
rect 144270 526940 144276 526952
rect 144328 526940 144334 526992
rect 150526 526940 150532 526992
rect 150584 526980 150590 526992
rect 178126 526980 178132 526992
rect 150584 526952 178132 526980
rect 150584 526940 150590 526952
rect 178126 526940 178132 526952
rect 178184 526940 178190 526992
rect 187970 526940 187976 526992
rect 188028 526980 188034 526992
rect 199378 526980 199384 526992
rect 188028 526952 199384 526980
rect 188028 526940 188034 526952
rect 199378 526940 199384 526952
rect 199436 526940 199442 526992
rect 204346 526940 204352 526992
rect 204404 526980 204410 526992
rect 231946 526980 231952 526992
rect 204404 526952 231952 526980
rect 204404 526940 204410 526952
rect 231946 526940 231952 526952
rect 232004 526940 232010 526992
rect 242066 526940 242072 526992
rect 242124 526980 242130 526992
rect 253198 526980 253204 526992
rect 242124 526952 253204 526980
rect 242124 526940 242130 526952
rect 253198 526940 253204 526952
rect 253256 526940 253262 526992
rect 258166 526940 258172 526992
rect 258224 526980 258230 526992
rect 258224 526952 279924 526980
rect 258224 526940 258230 526952
rect 122926 526872 122932 526924
rect 122984 526912 122990 526924
rect 150710 526912 150716 526924
rect 122984 526884 150716 526912
rect 122984 526872 122990 526884
rect 150710 526872 150716 526884
rect 150768 526872 150774 526924
rect 160554 526872 160560 526924
rect 160612 526912 160618 526924
rect 171778 526912 171784 526924
rect 160612 526884 171784 526912
rect 160612 526872 160618 526884
rect 171778 526872 171784 526884
rect 171836 526872 171842 526924
rect 215018 526872 215024 526924
rect 215076 526912 215082 526924
rect 225598 526912 225604 526924
rect 215076 526884 225604 526912
rect 215076 526872 215082 526884
rect 225598 526872 225604 526884
rect 225656 526872 225662 526924
rect 268930 526872 268936 526924
rect 268988 526912 268994 526924
rect 279418 526912 279424 526924
rect 268988 526884 279424 526912
rect 268988 526872 268994 526884
rect 279418 526872 279424 526884
rect 279476 526872 279482 526924
rect 279896 526912 279924 526952
rect 285766 526940 285772 526992
rect 285824 526980 285830 526992
rect 312630 526980 312636 526992
rect 285824 526952 312636 526980
rect 285824 526940 285830 526952
rect 312630 526940 312636 526952
rect 312688 526940 312694 526992
rect 340138 526980 340144 526992
rect 316006 526952 340144 526980
rect 286134 526912 286140 526924
rect 279896 526884 286140 526912
rect 286134 526872 286140 526884
rect 286192 526872 286198 526924
rect 295978 526872 295984 526924
rect 296036 526912 296042 526924
rect 307018 526912 307024 526924
rect 296036 526884 307024 526912
rect 296036 526872 296042 526884
rect 307018 526872 307024 526884
rect 307076 526872 307082 526924
rect 311986 526872 311992 526924
rect 312044 526912 312050 526924
rect 316006 526912 316034 526952
rect 340138 526940 340144 526952
rect 340196 526940 340202 526992
rect 366726 526980 366732 526992
rect 344986 526952 366732 526980
rect 312044 526884 316034 526912
rect 312044 526872 312050 526884
rect 322842 526872 322848 526924
rect 322900 526912 322906 526924
rect 333238 526912 333244 526924
rect 322900 526884 333244 526912
rect 322900 526872 322906 526884
rect 333238 526872 333244 526884
rect 333296 526872 333302 526924
rect 339586 526872 339592 526924
rect 339644 526912 339650 526924
rect 344986 526912 345014 526952
rect 366726 526940 366732 526952
rect 366784 526940 366790 526992
rect 393590 526980 393596 526992
rect 373966 526952 393596 526980
rect 339644 526884 345014 526912
rect 339644 526872 339650 526884
rect 350074 526872 350080 526924
rect 350132 526912 350138 526924
rect 359550 526912 359556 526924
rect 350132 526884 359556 526912
rect 350132 526872 350138 526884
rect 359550 526872 359556 526884
rect 359608 526872 359614 526924
rect 365806 526872 365812 526924
rect 365864 526912 365870 526924
rect 373966 526912 373994 526952
rect 393590 526940 393596 526952
rect 393648 526940 393654 526992
rect 420914 526980 420920 526992
rect 402946 526952 420920 526980
rect 365864 526884 373994 526912
rect 365864 526872 365870 526884
rect 376570 526872 376576 526924
rect 376628 526912 376634 526924
rect 387058 526912 387064 526924
rect 376628 526884 387064 526912
rect 376628 526872 376634 526884
rect 387058 526872 387064 526884
rect 387116 526872 387122 526924
rect 393406 526872 393412 526924
rect 393464 526912 393470 526924
rect 402946 526912 402974 526952
rect 420914 526940 420920 526952
rect 420972 526940 420978 526992
rect 431034 526940 431040 526992
rect 431092 526980 431098 526992
rect 442258 526980 442264 526992
rect 431092 526952 442264 526980
rect 431092 526940 431098 526952
rect 442258 526940 442264 526952
rect 442316 526940 442322 526992
rect 447226 526940 447232 526992
rect 447284 526980 447290 526992
rect 474734 526980 474740 526992
rect 447284 526952 474740 526980
rect 447284 526940 447290 526952
rect 474734 526940 474740 526952
rect 474792 526940 474798 526992
rect 484946 526940 484952 526992
rect 485004 526980 485010 526992
rect 496078 526980 496084 526992
rect 485004 526952 496084 526980
rect 485004 526940 485010 526952
rect 496078 526940 496084 526952
rect 496136 526940 496142 526992
rect 501046 526940 501052 526992
rect 501104 526980 501110 526992
rect 528646 526980 528652 526992
rect 501104 526952 528652 526980
rect 501104 526940 501110 526952
rect 528646 526940 528652 526952
rect 528704 526940 528710 526992
rect 393464 526884 402974 526912
rect 393464 526872 393470 526884
rect 403986 526872 403992 526924
rect 404044 526912 404050 526924
rect 414658 526912 414664 526924
rect 404044 526884 414664 526912
rect 404044 526872 404050 526884
rect 414658 526872 414664 526884
rect 414716 526872 414722 526924
rect 458082 526872 458088 526924
rect 458140 526912 458146 526924
rect 468570 526912 468576 526924
rect 458140 526884 468576 526912
rect 458140 526872 458146 526884
rect 468570 526872 468576 526884
rect 468628 526872 468634 526924
rect 511810 526872 511816 526924
rect 511868 526912 511874 526924
rect 522390 526912 522396 526924
rect 511868 526884 522396 526912
rect 511868 526872 511874 526884
rect 522390 526872 522396 526884
rect 522448 526872 522454 526924
rect 36538 526804 36544 526856
rect 36596 526844 36602 526856
rect 538398 526844 538404 526856
rect 36596 526816 538404 526844
rect 36596 526804 36602 526816
rect 538398 526804 538404 526816
rect 538456 526804 538462 526856
rect 527082 525716 527088 525768
rect 527140 525756 527146 525768
rect 579798 525756 579804 525768
rect 527140 525728 579804 525756
rect 527140 525716 527146 525728
rect 579798 525716 579804 525728
rect 579856 525716 579862 525768
rect 16298 523676 16304 523728
rect 16356 523716 16362 523728
rect 528738 523716 528744 523728
rect 16356 523688 528744 523716
rect 16356 523676 16362 523688
rect 528738 523676 528744 523688
rect 528796 523676 528802 523728
rect 25958 523268 25964 523320
rect 26016 523308 26022 523320
rect 149698 523308 149704 523320
rect 26016 523280 149704 523308
rect 26016 523268 26022 523280
rect 149698 523268 149704 523280
rect 149756 523268 149762 523320
rect 36814 523200 36820 523252
rect 36872 523240 36878 523252
rect 52454 523240 52460 523252
rect 36872 523212 52460 523240
rect 36872 523200 36878 523212
rect 52454 523200 52460 523212
rect 52512 523200 52518 523252
rect 232314 523200 232320 523252
rect 232372 523240 232378 523252
rect 251818 523240 251824 523252
rect 232372 523212 251824 523240
rect 232372 523200 232378 523212
rect 251818 523200 251824 523212
rect 251876 523200 251882 523252
rect 475378 523200 475384 523252
rect 475436 523240 475442 523252
rect 494698 523240 494704 523252
rect 475436 523212 494704 523240
rect 475436 523200 475442 523212
rect 494698 523200 494704 523212
rect 494756 523200 494762 523252
rect 62482 523132 62488 523184
rect 62540 523172 62546 523184
rect 79318 523172 79324 523184
rect 62540 523144 79324 523172
rect 62540 523132 62546 523144
rect 79318 523132 79324 523144
rect 79376 523132 79382 523184
rect 90450 523132 90456 523184
rect 90508 523172 90514 523184
rect 106366 523172 106372 523184
rect 90508 523144 106372 523172
rect 90508 523132 90514 523144
rect 106366 523132 106372 523144
rect 106424 523132 106430 523184
rect 116486 523132 116492 523184
rect 116544 523172 116550 523184
rect 133414 523172 133420 523184
rect 116544 523144 133420 523172
rect 116544 523132 116550 523144
rect 133414 523132 133420 523144
rect 133472 523132 133478 523184
rect 144178 523132 144184 523184
rect 144236 523172 144242 523184
rect 160278 523172 160284 523184
rect 144236 523144 160284 523172
rect 144236 523132 144242 523144
rect 160278 523132 160284 523144
rect 160336 523132 160342 523184
rect 170490 523132 170496 523184
rect 170548 523172 170554 523184
rect 187786 523172 187792 523184
rect 170548 523144 187792 523172
rect 170548 523132 170554 523144
rect 187786 523132 187792 523144
rect 187844 523132 187850 523184
rect 197538 523132 197544 523184
rect 197596 523172 197602 523184
rect 214374 523172 214380 523184
rect 197596 523144 214380 523172
rect 197596 523132 197602 523144
rect 214374 523132 214380 523144
rect 214432 523132 214438 523184
rect 224494 523132 224500 523184
rect 224552 523172 224558 523184
rect 241514 523172 241520 523184
rect 224552 523144 241520 523172
rect 224552 523132 224558 523144
rect 241514 523132 241520 523144
rect 241572 523132 241578 523184
rect 413462 523132 413468 523184
rect 413520 523172 413526 523184
rect 430574 523172 430580 523184
rect 413520 523144 430580 523172
rect 413520 523132 413526 523144
rect 430574 523132 430580 523144
rect 430632 523132 430638 523184
rect 440510 523132 440516 523184
rect 440568 523172 440574 523184
rect 457254 523172 457260 523184
rect 440568 523144 457260 523172
rect 440568 523132 440574 523144
rect 457254 523132 457260 523144
rect 457312 523132 457318 523184
rect 468478 523132 468484 523184
rect 468536 523172 468542 523184
rect 484394 523172 484400 523184
rect 468536 523144 484400 523172
rect 468536 523132 468542 523144
rect 484394 523132 484400 523144
rect 484452 523132 484458 523184
rect 36538 523064 36544 523116
rect 36596 523104 36602 523116
rect 62114 523104 62120 523116
rect 36596 523076 62120 523104
rect 36596 523064 36602 523076
rect 62114 523064 62120 523076
rect 62172 523064 62178 523116
rect 64138 523064 64144 523116
rect 64196 523104 64202 523116
rect 89070 523104 89076 523116
rect 64196 523076 89076 523104
rect 64196 523064 64202 523076
rect 89070 523064 89076 523076
rect 89128 523064 89134 523116
rect 90358 523064 90364 523116
rect 90416 523104 90422 523116
rect 115934 523104 115940 523116
rect 90416 523076 115940 523104
rect 90416 523064 90422 523076
rect 115934 523064 115940 523076
rect 115992 523064 115998 523116
rect 116578 523064 116584 523116
rect 116636 523104 116642 523116
rect 142982 523104 142988 523116
rect 116636 523076 142988 523104
rect 116636 523064 116642 523076
rect 142982 523064 142988 523076
rect 143040 523064 143046 523116
rect 144270 523064 144276 523116
rect 144328 523104 144334 523116
rect 170030 523104 170036 523116
rect 144328 523076 170036 523104
rect 144328 523064 144334 523076
rect 170030 523064 170036 523076
rect 170088 523064 170094 523116
rect 178402 523064 178408 523116
rect 178460 523104 178466 523116
rect 200758 523104 200764 523116
rect 178460 523076 200764 523104
rect 178460 523064 178466 523076
rect 200758 523064 200764 523076
rect 200816 523064 200822 523116
rect 251450 523064 251456 523116
rect 251508 523104 251514 523116
rect 268286 523104 268292 523116
rect 251508 523076 268292 523104
rect 251508 523064 251514 523076
rect 268286 523064 268292 523076
rect 268344 523064 268350 523116
rect 279510 523064 279516 523116
rect 279568 523104 279574 523116
rect 295794 523104 295800 523116
rect 279568 523076 295800 523104
rect 279568 523064 279574 523076
rect 295794 523064 295800 523076
rect 295852 523064 295858 523116
rect 305546 523064 305552 523116
rect 305604 523104 305610 523116
rect 322382 523104 322388 523116
rect 305604 523076 322388 523104
rect 305604 523064 305610 523076
rect 322382 523064 322388 523076
rect 322440 523064 322446 523116
rect 334618 523064 334624 523116
rect 334676 523104 334682 523116
rect 349798 523104 349804 523116
rect 334676 523076 349804 523104
rect 334676 523064 334682 523076
rect 349798 523064 349804 523076
rect 349856 523064 349862 523116
rect 359550 523064 359556 523116
rect 359608 523104 359614 523116
rect 376294 523104 376300 523116
rect 359608 523076 376300 523104
rect 359608 523064 359614 523076
rect 376294 523064 376300 523076
rect 376352 523064 376358 523116
rect 386506 523064 386512 523116
rect 386564 523104 386570 523116
rect 403342 523104 403348 523116
rect 386564 523076 403348 523104
rect 386564 523064 386570 523076
rect 403342 523064 403348 523076
rect 403400 523064 403406 523116
rect 421282 523064 421288 523116
rect 421340 523104 421346 523116
rect 443638 523104 443644 523116
rect 421340 523076 443644 523104
rect 421340 523064 421346 523076
rect 443638 523064 443644 523076
rect 443696 523064 443702 523116
rect 494514 523064 494520 523116
rect 494572 523104 494578 523116
rect 511350 523104 511356 523116
rect 494572 523076 511356 523104
rect 494572 523064 494578 523076
rect 511350 523064 511356 523076
rect 511408 523064 511414 523116
rect 522390 523064 522396 523116
rect 522448 523104 522454 523116
rect 538398 523104 538404 523116
rect 522448 523076 538404 523104
rect 522448 523064 522454 523076
rect 538398 523064 538404 523076
rect 538456 523064 538462 523116
rect 43346 522996 43352 523048
rect 43404 523036 43410 523048
rect 62758 523036 62764 523048
rect 43404 523008 62764 523036
rect 43404 522996 43410 523008
rect 62758 522996 62764 523008
rect 62816 522996 62822 523048
rect 171778 522996 171784 523048
rect 171836 523036 171842 523048
rect 197446 523036 197452 523048
rect 171836 523008 197452 523036
rect 171836 522996 171842 523008
rect 197446 522996 197452 523008
rect 197504 522996 197510 523048
rect 199378 522996 199384 523048
rect 199436 523036 199442 523048
rect 223942 523036 223948 523048
rect 199436 523008 223948 523036
rect 199436 522996 199442 523008
rect 223942 522996 223948 523008
rect 224000 522996 224006 523048
rect 225598 522996 225604 523048
rect 225656 523036 225662 523048
rect 251174 523036 251180 523048
rect 225656 523008 251180 523036
rect 225656 522996 225662 523008
rect 251174 522996 251180 523008
rect 251232 522996 251238 523048
rect 253198 522996 253204 523048
rect 253256 523036 253262 523048
rect 278038 523036 278044 523048
rect 253256 523008 278044 523036
rect 253256 522996 253262 523008
rect 278038 522996 278044 523008
rect 278096 522996 278102 523048
rect 279418 522996 279424 523048
rect 279476 523036 279482 523048
rect 305454 523036 305460 523048
rect 279476 523008 305460 523036
rect 279476 522996 279482 523008
rect 305454 522996 305460 523008
rect 305512 522996 305518 523048
rect 307018 522996 307024 523048
rect 307076 523036 307082 523048
rect 331950 523036 331956 523048
rect 307076 523008 331956 523036
rect 307076 522996 307082 523008
rect 331950 522996 331956 523008
rect 332008 522996 332014 523048
rect 333238 522996 333244 523048
rect 333296 523036 333302 523048
rect 359458 523036 359464 523048
rect 333296 523008 359464 523036
rect 333296 522996 333302 523008
rect 359458 522996 359464 523008
rect 359516 522996 359522 523048
rect 359734 522996 359740 523048
rect 359792 523036 359798 523048
rect 386046 523036 386052 523048
rect 359792 523008 386052 523036
rect 359792 522996 359798 523008
rect 386046 522996 386052 523008
rect 386104 522996 386110 523048
rect 387058 522996 387064 523048
rect 387116 523036 387122 523048
rect 412910 523036 412916 523048
rect 387116 523008 412916 523036
rect 387116 522996 387122 523008
rect 412910 522996 412916 523008
rect 412968 522996 412974 523048
rect 414658 522996 414664 523048
rect 414716 523036 414722 523048
rect 440234 523036 440240 523048
rect 414716 523008 440240 523036
rect 414716 522996 414722 523008
rect 440234 522996 440240 523008
rect 440292 522996 440298 523048
rect 442258 522996 442264 523048
rect 442316 523036 442322 523048
rect 467006 523036 467012 523048
rect 442316 523008 467012 523036
rect 442316 522996 442322 523008
rect 467006 522996 467012 523008
rect 467064 522996 467070 523048
rect 468570 522996 468576 523048
rect 468628 523036 468634 523048
rect 494054 523036 494060 523048
rect 468628 523008 494060 523036
rect 468628 522996 468634 523008
rect 494054 522996 494060 523008
rect 494112 522996 494118 523048
rect 496078 522996 496084 523048
rect 496136 523036 496142 523048
rect 520918 523036 520924 523048
rect 496136 523008 520924 523036
rect 496136 522996 496142 523008
rect 520918 522996 520924 523008
rect 520976 522996 520982 523048
rect 522298 522996 522304 523048
rect 522356 523036 522362 523048
rect 548058 523036 548064 523048
rect 522356 523008 548064 523036
rect 522356 522996 522362 523008
rect 548058 522996 548064 523008
rect 548116 522996 548122 523048
rect 37918 522248 37924 522300
rect 37976 522288 37982 522300
rect 526438 522288 526444 522300
rect 37976 522260 526444 522288
rect 37976 522248 37982 522260
rect 526438 522248 526444 522260
rect 526496 522248 526502 522300
rect 35618 521704 35624 521756
rect 35676 521744 35682 521756
rect 36630 521744 36636 521756
rect 35676 521716 36636 521744
rect 35676 521704 35682 521716
rect 36630 521704 36636 521716
rect 36688 521704 36694 521756
rect 285766 521364 285772 521416
rect 285824 521404 285830 521416
rect 286134 521404 286140 521416
rect 285824 521376 286140 521404
rect 285824 521364 285830 521376
rect 286134 521364 286140 521376
rect 286192 521364 286198 521416
rect 339586 521296 339592 521348
rect 339644 521336 339650 521348
rect 340138 521336 340144 521348
rect 339644 521308 340144 521336
rect 339644 521296 339650 521308
rect 340138 521296 340144 521308
rect 340196 521296 340202 521348
rect 68922 520412 68928 520464
rect 68980 520452 68986 520464
rect 118694 520452 118700 520464
rect 68980 520424 118700 520452
rect 68980 520412 68986 520424
rect 118694 520412 118700 520424
rect 118752 520412 118758 520464
rect 311802 520412 311808 520464
rect 311860 520452 311866 520464
rect 361574 520452 361580 520464
rect 311860 520424 361580 520452
rect 311860 520412 311866 520424
rect 361574 520412 361580 520424
rect 361632 520412 361638 520464
rect 41322 520344 41328 520396
rect 41380 520384 41386 520396
rect 91094 520384 91100 520396
rect 41380 520356 91100 520384
rect 41380 520344 41386 520356
rect 91094 520344 91100 520356
rect 91152 520344 91158 520396
rect 122742 520344 122748 520396
rect 122800 520384 122806 520396
rect 172514 520384 172520 520396
rect 122800 520356 172520 520384
rect 122800 520344 122806 520356
rect 172514 520344 172520 520356
rect 172572 520344 172578 520396
rect 176562 520344 176568 520396
rect 176620 520384 176626 520396
rect 226334 520384 226340 520396
rect 176620 520356 226340 520384
rect 176620 520344 176626 520356
rect 226334 520344 226340 520356
rect 226392 520344 226398 520396
rect 231854 520344 231860 520396
rect 231912 520384 231918 520396
rect 280154 520384 280160 520396
rect 231912 520356 280160 520384
rect 231912 520344 231918 520356
rect 280154 520344 280160 520356
rect 280212 520344 280218 520396
rect 284202 520344 284208 520396
rect 284260 520384 284266 520396
rect 335354 520384 335360 520396
rect 284260 520356 335360 520384
rect 284260 520344 284266 520356
rect 335354 520344 335360 520356
rect 335412 520344 335418 520396
rect 365622 520344 365628 520396
rect 365680 520384 365686 520396
rect 415394 520384 415400 520396
rect 365680 520356 415400 520384
rect 365680 520344 365686 520356
rect 415394 520344 415400 520356
rect 415452 520344 415458 520396
rect 419442 520344 419448 520396
rect 419500 520384 419506 520396
rect 469214 520384 469220 520396
rect 419500 520356 469220 520384
rect 419500 520344 419506 520356
rect 469214 520344 469220 520356
rect 469272 520344 469278 520396
rect 474826 520344 474832 520396
rect 474884 520384 474890 520396
rect 523034 520384 523040 520396
rect 474884 520356 523040 520384
rect 474884 520344 474890 520356
rect 523034 520344 523040 520356
rect 523092 520344 523098 520396
rect 13722 520276 13728 520328
rect 13780 520316 13786 520328
rect 64874 520316 64880 520328
rect 13780 520288 64880 520316
rect 13780 520276 13786 520288
rect 64874 520276 64880 520288
rect 64932 520276 64938 520328
rect 96890 520276 96896 520328
rect 96948 520316 96954 520328
rect 146294 520316 146300 520328
rect 96948 520288 146300 520316
rect 96948 520276 96954 520288
rect 146294 520276 146300 520288
rect 146352 520276 146358 520328
rect 148962 520276 148968 520328
rect 149020 520316 149026 520328
rect 200114 520316 200120 520328
rect 149020 520288 200120 520316
rect 149020 520276 149026 520288
rect 200114 520276 200120 520288
rect 200172 520276 200178 520328
rect 204898 520276 204904 520328
rect 204956 520316 204962 520328
rect 253934 520316 253940 520328
rect 204956 520288 253940 520316
rect 204956 520276 204962 520288
rect 253934 520276 253940 520288
rect 253992 520276 253998 520328
rect 256602 520276 256608 520328
rect 256660 520316 256666 520328
rect 307754 520316 307760 520328
rect 256660 520288 307760 520316
rect 256660 520276 256666 520288
rect 307754 520276 307760 520288
rect 307812 520276 307818 520328
rect 339862 520276 339868 520328
rect 339920 520316 339926 520328
rect 389174 520316 389180 520328
rect 339920 520288 389180 520316
rect 339920 520276 339926 520288
rect 389174 520276 389180 520288
rect 389232 520276 389238 520328
rect 391842 520276 391848 520328
rect 391900 520316 391906 520328
rect 442994 520316 443000 520328
rect 391900 520288 443000 520316
rect 391900 520276 391906 520288
rect 442994 520276 443000 520288
rect 443052 520276 443058 520328
rect 445662 520276 445668 520328
rect 445720 520316 445726 520328
rect 496814 520316 496820 520328
rect 445720 520288 496820 520316
rect 445720 520276 445726 520288
rect 496814 520276 496820 520288
rect 496872 520276 496878 520328
rect 500862 520276 500868 520328
rect 500920 520316 500926 520328
rect 550634 520316 550640 520328
rect 500920 520288 550640 520316
rect 500920 520276 500926 520288
rect 550634 520276 550640 520288
rect 550692 520276 550698 520328
rect 230382 518848 230388 518900
rect 230440 518888 230446 518900
rect 231854 518888 231860 518900
rect 230440 518860 231860 518888
rect 230440 518848 230446 518860
rect 231854 518848 231860 518860
rect 231912 518848 231918 518900
rect 473262 518848 473268 518900
rect 473320 518888 473326 518900
rect 474826 518888 474832 518900
rect 473320 518860 474832 518888
rect 473320 518848 473326 518860
rect 474826 518848 474832 518860
rect 474884 518848 474890 518900
rect 89714 505588 89720 505640
rect 89772 505628 89778 505640
rect 90450 505628 90456 505640
rect 89772 505600 90456 505628
rect 89772 505588 89778 505600
rect 90450 505588 90456 505600
rect 90508 505588 90514 505640
rect 521746 505588 521752 505640
rect 521804 505628 521810 505640
rect 522390 505628 522396 505640
rect 521804 505600 522396 505628
rect 521804 505588 521810 505600
rect 522390 505588 522396 505600
rect 522448 505588 522454 505640
rect 278682 503616 278688 503668
rect 278740 503656 278746 503668
rect 279510 503656 279516 503668
rect 278740 503628 279516 503656
rect 278740 503616 278746 503628
rect 279510 503616 279516 503628
rect 279568 503616 279574 503668
rect 332502 503616 332508 503668
rect 332560 503656 332566 503668
rect 334618 503656 334624 503668
rect 332560 503628 334624 503656
rect 332560 503616 332566 503628
rect 334618 503616 334624 503628
rect 334676 503616 334682 503668
rect 35618 502256 35624 502308
rect 35676 502296 35682 502308
rect 36814 502296 36820 502308
rect 35676 502268 36820 502296
rect 35676 502256 35682 502268
rect 36814 502256 36820 502268
rect 36872 502256 36878 502308
rect 52730 500896 52736 500948
rect 52788 500936 52794 500948
rect 64138 500936 64144 500948
rect 52788 500908 64144 500936
rect 52788 500896 52794 500908
rect 64138 500896 64144 500908
rect 64196 500896 64202 500948
rect 69106 500896 69112 500948
rect 69164 500936 69170 500948
rect 69164 500908 74534 500936
rect 69164 500896 69170 500908
rect 15194 500828 15200 500880
rect 15252 500868 15258 500880
rect 42978 500868 42984 500880
rect 15252 500840 42984 500868
rect 15252 500828 15258 500840
rect 42978 500828 42984 500840
rect 43036 500828 43042 500880
rect 62758 500828 62764 500880
rect 62816 500868 62822 500880
rect 70026 500868 70032 500880
rect 62816 500840 70032 500868
rect 62816 500828 62822 500840
rect 70026 500828 70032 500840
rect 70084 500828 70090 500880
rect 74506 500868 74534 500908
rect 96706 500896 96712 500948
rect 96764 500936 96770 500948
rect 96764 500908 103514 500936
rect 96764 500896 96770 500908
rect 96982 500868 96988 500880
rect 74506 500840 96988 500868
rect 96982 500828 96988 500840
rect 97040 500828 97046 500880
rect 103486 500868 103514 500908
rect 146938 500896 146944 500948
rect 146996 500936 147002 500948
rect 146996 500908 151814 500936
rect 146996 500896 147002 500908
rect 124030 500868 124036 500880
rect 103486 500840 124036 500868
rect 124030 500828 124036 500840
rect 124088 500828 124094 500880
rect 133690 500828 133696 500880
rect 133748 500868 133754 500880
rect 144270 500868 144276 500880
rect 133748 500840 144276 500868
rect 133748 500828 133754 500840
rect 144270 500828 144276 500840
rect 144328 500828 144334 500880
rect 150986 500868 150992 500880
rect 146588 500840 150992 500868
rect 25682 500760 25688 500812
rect 25740 500800 25746 500812
rect 36538 500800 36544 500812
rect 25740 500772 36544 500800
rect 25740 500760 25746 500772
rect 36538 500760 36544 500772
rect 36596 500760 36602 500812
rect 79686 500760 79692 500812
rect 79744 500800 79750 500812
rect 90358 500800 90364 500812
rect 79744 500772 90364 500800
rect 79744 500760 79750 500772
rect 90358 500760 90364 500772
rect 90416 500760 90422 500812
rect 106642 500760 106648 500812
rect 106700 500800 106706 500812
rect 116578 500800 116584 500812
rect 106700 500772 116584 500800
rect 106700 500760 106706 500772
rect 116578 500760 116584 500772
rect 116636 500760 116642 500812
rect 122926 500760 122932 500812
rect 122984 500800 122990 500812
rect 146588 500800 146616 500840
rect 150986 500828 150992 500840
rect 151044 500828 151050 500880
rect 151786 500868 151814 500908
rect 200758 500896 200764 500948
rect 200816 500936 200822 500948
rect 204990 500936 204996 500948
rect 200816 500908 204996 500936
rect 200816 500896 200822 500908
rect 204990 500896 204996 500908
rect 205048 500896 205054 500948
rect 251818 500896 251824 500948
rect 251876 500936 251882 500948
rect 258994 500936 259000 500948
rect 251876 500908 259000 500936
rect 251876 500896 251882 500908
rect 258994 500896 259000 500908
rect 259052 500896 259058 500948
rect 443638 500896 443644 500948
rect 443696 500936 443702 500948
rect 447962 500936 447968 500948
rect 443696 500908 447968 500936
rect 443696 500896 443702 500908
rect 447962 500896 447968 500908
rect 448020 500896 448026 500948
rect 494698 500896 494704 500948
rect 494756 500936 494762 500948
rect 501966 500936 501972 500948
rect 494756 500908 501972 500936
rect 494756 500896 494762 500908
rect 501966 500896 501972 500908
rect 502024 500896 502030 500948
rect 548334 500868 548340 500880
rect 151786 500840 548340 500868
rect 548334 500828 548340 500840
rect 548392 500828 548398 500880
rect 122984 500772 146616 500800
rect 122984 500760 122990 500772
rect 150526 500760 150532 500812
rect 150584 500800 150590 500812
rect 178034 500800 178040 500812
rect 150584 500772 178040 500800
rect 150584 500760 150590 500772
rect 178034 500760 178040 500772
rect 178092 500760 178098 500812
rect 187694 500760 187700 500812
rect 187752 500800 187758 500812
rect 199378 500800 199384 500812
rect 187752 500772 199384 500800
rect 187752 500760 187758 500772
rect 199378 500760 199384 500772
rect 199436 500760 199442 500812
rect 204346 500760 204352 500812
rect 204404 500800 204410 500812
rect 232038 500800 232044 500812
rect 204404 500772 232044 500800
rect 204404 500760 204410 500772
rect 232038 500760 232044 500772
rect 232096 500760 232102 500812
rect 241698 500760 241704 500812
rect 241756 500800 241762 500812
rect 253198 500800 253204 500812
rect 241756 500772 253204 500800
rect 241756 500760 241762 500772
rect 253198 500760 253204 500772
rect 253256 500760 253262 500812
rect 258166 500760 258172 500812
rect 258224 500800 258230 500812
rect 258224 500772 281764 500800
rect 258224 500760 258230 500772
rect 160646 500692 160652 500744
rect 160704 500732 160710 500744
rect 171778 500732 171784 500744
rect 160704 500704 171784 500732
rect 160704 500692 160710 500704
rect 171778 500692 171784 500704
rect 171836 500692 171842 500744
rect 214650 500692 214656 500744
rect 214708 500732 214714 500744
rect 225598 500732 225604 500744
rect 214708 500704 225604 500732
rect 214708 500692 214714 500704
rect 225598 500692 225604 500704
rect 225656 500692 225662 500744
rect 268654 500692 268660 500744
rect 268712 500732 268718 500744
rect 279418 500732 279424 500744
rect 268712 500704 279424 500732
rect 268712 500692 268718 500704
rect 279418 500692 279424 500704
rect 279476 500692 279482 500744
rect 281736 500732 281764 500772
rect 285766 500760 285772 500812
rect 285824 500800 285830 500812
rect 312998 500800 313004 500812
rect 285824 500772 313004 500800
rect 285824 500760 285830 500772
rect 312998 500760 313004 500772
rect 313056 500760 313062 500812
rect 340046 500800 340052 500812
rect 316006 500772 340052 500800
rect 286042 500732 286048 500744
rect 281736 500704 286048 500732
rect 286042 500692 286048 500704
rect 286100 500692 286106 500744
rect 295702 500692 295708 500744
rect 295760 500732 295766 500744
rect 307018 500732 307024 500744
rect 295760 500704 307024 500732
rect 295760 500692 295766 500704
rect 307018 500692 307024 500704
rect 307076 500692 307082 500744
rect 311986 500692 311992 500744
rect 312044 500732 312050 500744
rect 316006 500732 316034 500772
rect 340046 500760 340052 500772
rect 340104 500760 340110 500812
rect 367002 500800 367008 500812
rect 344986 500772 367008 500800
rect 312044 500704 316034 500732
rect 312044 500692 312050 500704
rect 322658 500692 322664 500744
rect 322716 500732 322722 500744
rect 333238 500732 333244 500744
rect 322716 500704 333244 500732
rect 322716 500692 322722 500704
rect 333238 500692 333244 500704
rect 333296 500692 333302 500744
rect 339586 500692 339592 500744
rect 339644 500732 339650 500744
rect 344986 500732 345014 500772
rect 367002 500760 367008 500772
rect 367060 500760 367066 500812
rect 393958 500800 393964 500812
rect 373966 500772 393964 500800
rect 339644 500704 345014 500732
rect 339644 500692 339650 500704
rect 349706 500692 349712 500744
rect 349764 500732 349770 500744
rect 359550 500732 359556 500744
rect 349764 500704 359556 500732
rect 349764 500692 349770 500704
rect 359550 500692 359556 500704
rect 359608 500692 359614 500744
rect 365806 500692 365812 500744
rect 365864 500732 365870 500744
rect 373966 500732 373994 500772
rect 393958 500760 393964 500772
rect 394016 500760 394022 500812
rect 421006 500800 421012 500812
rect 402946 500772 421012 500800
rect 365864 500704 373994 500732
rect 365864 500692 365870 500704
rect 376662 500692 376668 500744
rect 376720 500732 376726 500744
rect 387058 500732 387064 500744
rect 376720 500704 387064 500732
rect 376720 500692 376726 500704
rect 387058 500692 387064 500704
rect 387116 500692 387122 500744
rect 393406 500692 393412 500744
rect 393464 500732 393470 500744
rect 402946 500732 402974 500772
rect 421006 500760 421012 500772
rect 421064 500760 421070 500812
rect 430666 500760 430672 500812
rect 430724 500800 430730 500812
rect 442258 500800 442264 500812
rect 430724 500772 442264 500800
rect 430724 500760 430730 500772
rect 442258 500760 442264 500772
rect 442316 500760 442322 500812
rect 447226 500760 447232 500812
rect 447284 500800 447290 500812
rect 475010 500800 475016 500812
rect 447284 500772 475016 500800
rect 447284 500760 447290 500772
rect 475010 500760 475016 500772
rect 475068 500760 475074 500812
rect 484670 500760 484676 500812
rect 484728 500800 484734 500812
rect 496078 500800 496084 500812
rect 484728 500772 496084 500800
rect 484728 500760 484734 500772
rect 496078 500760 496084 500772
rect 496136 500760 496142 500812
rect 501046 500760 501052 500812
rect 501104 500800 501110 500812
rect 529014 500800 529020 500812
rect 501104 500772 529020 500800
rect 501104 500760 501110 500772
rect 529014 500760 529020 500772
rect 529072 500760 529078 500812
rect 393464 500704 402974 500732
rect 393464 500692 393470 500704
rect 403710 500692 403716 500744
rect 403768 500732 403774 500744
rect 414658 500732 414664 500744
rect 403768 500704 414664 500732
rect 403768 500692 403774 500704
rect 414658 500692 414664 500704
rect 414716 500692 414722 500744
rect 457714 500692 457720 500744
rect 457772 500732 457778 500744
rect 468570 500732 468576 500744
rect 457772 500704 468576 500732
rect 457772 500692 457778 500704
rect 468570 500692 468576 500704
rect 468628 500692 468634 500744
rect 511718 500692 511724 500744
rect 511776 500732 511782 500744
rect 522298 500732 522304 500744
rect 511776 500704 522304 500732
rect 511776 500692 511782 500704
rect 522298 500692 522304 500704
rect 522356 500692 522362 500744
rect 36722 500624 36728 500676
rect 36780 500664 36786 500676
rect 538674 500664 538680 500676
rect 36780 500636 538680 500664
rect 36780 500624 36786 500636
rect 538674 500624 538680 500636
rect 538732 500624 538738 500676
rect 16022 497428 16028 497480
rect 16080 497468 16086 497480
rect 529014 497468 529020 497480
rect 16080 497440 529020 497468
rect 16080 497428 16086 497440
rect 529014 497428 529020 497440
rect 529072 497428 529078 497480
rect 25682 497088 25688 497140
rect 25740 497128 25746 497140
rect 146938 497128 146944 497140
rect 25740 497100 146944 497128
rect 25740 497088 25746 497100
rect 146938 497088 146944 497100
rect 146996 497088 147002 497140
rect 36722 497020 36728 497072
rect 36780 497060 36786 497072
rect 52638 497060 52644 497072
rect 36780 497032 52644 497060
rect 36780 497020 36786 497032
rect 52638 497020 52644 497032
rect 52696 497020 52702 497072
rect 232038 497020 232044 497072
rect 232096 497060 232102 497072
rect 251818 497060 251824 497072
rect 232096 497032 251824 497060
rect 232096 497020 232102 497032
rect 251818 497020 251824 497032
rect 251876 497020 251882 497072
rect 475010 497020 475016 497072
rect 475068 497060 475074 497072
rect 494698 497060 494704 497072
rect 475068 497032 494704 497060
rect 475068 497020 475074 497032
rect 494698 497020 494704 497032
rect 494756 497020 494762 497072
rect 62482 496952 62488 497004
rect 62540 496992 62546 497004
rect 79686 496992 79692 497004
rect 62540 496964 79692 496992
rect 62540 496952 62546 496964
rect 79686 496952 79692 496964
rect 79744 496952 79750 497004
rect 90358 496952 90364 497004
rect 90416 496992 90422 497004
rect 106642 496992 106648 497004
rect 90416 496964 106648 496992
rect 90416 496952 90422 496964
rect 106642 496952 106648 496964
rect 106700 496952 106706 497004
rect 116486 496952 116492 497004
rect 116544 496992 116550 497004
rect 133690 496992 133696 497004
rect 116544 496964 133696 496992
rect 116544 496952 116550 496964
rect 133690 496952 133696 496964
rect 133748 496952 133754 497004
rect 170490 496952 170496 497004
rect 170548 496992 170554 497004
rect 187694 496992 187700 497004
rect 170548 496964 187700 496992
rect 170548 496952 170554 496964
rect 187694 496952 187700 496964
rect 187752 496952 187758 497004
rect 197446 496952 197452 497004
rect 197504 496992 197510 497004
rect 214650 496992 214656 497004
rect 197504 496964 214656 496992
rect 197504 496952 197510 496964
rect 214650 496952 214656 496964
rect 214708 496952 214714 497004
rect 224494 496952 224500 497004
rect 224552 496992 224558 497004
rect 241698 496992 241704 497004
rect 224552 496964 241704 496992
rect 224552 496952 224558 496964
rect 241698 496952 241704 496964
rect 241756 496952 241762 497004
rect 413462 496952 413468 497004
rect 413520 496992 413526 497004
rect 430666 496992 430672 497004
rect 413520 496964 430672 496992
rect 413520 496952 413526 496964
rect 430666 496952 430672 496964
rect 430724 496952 430730 497004
rect 440510 496952 440516 497004
rect 440568 496992 440574 497004
rect 457622 496992 457628 497004
rect 440568 496964 457628 496992
rect 440568 496952 440574 496964
rect 457622 496952 457628 496964
rect 457680 496952 457686 497004
rect 468570 496952 468576 497004
rect 468628 496992 468634 497004
rect 484670 496992 484676 497004
rect 468628 496964 484676 496992
rect 468628 496952 468634 496964
rect 484670 496952 484676 496964
rect 484728 496952 484734 497004
rect 36814 496884 36820 496936
rect 36872 496924 36878 496936
rect 62298 496924 62304 496936
rect 36872 496896 62304 496924
rect 36872 496884 36878 496896
rect 62298 496884 62304 496896
rect 62356 496884 62362 496936
rect 64138 496884 64144 496936
rect 64196 496924 64202 496936
rect 89346 496924 89352 496936
rect 64196 496896 89352 496924
rect 64196 496884 64202 496896
rect 89346 496884 89352 496896
rect 89404 496884 89410 496936
rect 90450 496884 90456 496936
rect 90508 496924 90514 496936
rect 116302 496924 116308 496936
rect 90508 496896 116308 496924
rect 90508 496884 90514 496896
rect 116302 496884 116308 496896
rect 116360 496884 116366 496936
rect 116578 496884 116584 496936
rect 116636 496924 116642 496936
rect 143350 496924 143356 496936
rect 116636 496896 143356 496924
rect 116636 496884 116642 496896
rect 143350 496884 143356 496896
rect 143408 496884 143414 496936
rect 144270 496884 144276 496936
rect 144328 496924 144334 496936
rect 170306 496924 170312 496936
rect 144328 496896 170312 496924
rect 144328 496884 144334 496896
rect 170306 496884 170312 496896
rect 170364 496884 170370 496936
rect 178034 496884 178040 496936
rect 178092 496924 178098 496936
rect 200758 496924 200764 496936
rect 178092 496896 200764 496924
rect 178092 496884 178098 496896
rect 200758 496884 200764 496896
rect 200816 496884 200822 496936
rect 251450 496884 251456 496936
rect 251508 496924 251514 496936
rect 268654 496924 268660 496936
rect 251508 496896 268660 496924
rect 251508 496884 251514 496896
rect 268654 496884 268660 496896
rect 268712 496884 268718 496936
rect 279510 496884 279516 496936
rect 279568 496924 279574 496936
rect 295702 496924 295708 496936
rect 279568 496896 295708 496924
rect 279568 496884 279574 496896
rect 295702 496884 295708 496896
rect 295760 496884 295766 496936
rect 305454 496884 305460 496936
rect 305512 496924 305518 496936
rect 322658 496924 322664 496936
rect 305512 496896 322664 496924
rect 305512 496884 305518 496896
rect 322658 496884 322664 496896
rect 322716 496884 322722 496936
rect 334618 496884 334624 496936
rect 334676 496924 334682 496936
rect 349706 496924 349712 496936
rect 334676 496896 349712 496924
rect 334676 496884 334682 496896
rect 349706 496884 349712 496896
rect 349764 496884 349770 496936
rect 359458 496884 359464 496936
rect 359516 496924 359522 496936
rect 376662 496924 376668 496936
rect 359516 496896 376668 496924
rect 359516 496884 359522 496896
rect 376662 496884 376668 496896
rect 376720 496884 376726 496936
rect 386506 496884 386512 496936
rect 386564 496924 386570 496936
rect 403618 496924 403624 496936
rect 386564 496896 403624 496924
rect 386564 496884 386570 496896
rect 403618 496884 403624 496896
rect 403676 496884 403682 496936
rect 421006 496884 421012 496936
rect 421064 496924 421070 496936
rect 443638 496924 443644 496936
rect 421064 496896 443644 496924
rect 421064 496884 421070 496896
rect 443638 496884 443644 496896
rect 443696 496884 443702 496936
rect 494514 496884 494520 496936
rect 494572 496924 494578 496936
rect 511626 496924 511632 496936
rect 494572 496896 511632 496924
rect 494572 496884 494578 496896
rect 511626 496884 511632 496896
rect 511684 496884 511690 496936
rect 522390 496884 522396 496936
rect 522448 496924 522454 496936
rect 538674 496924 538680 496936
rect 522448 496896 538680 496924
rect 522448 496884 522454 496896
rect 538674 496884 538680 496896
rect 538732 496884 538738 496936
rect 43070 496816 43076 496868
rect 43128 496856 43134 496868
rect 62758 496856 62764 496868
rect 43128 496828 62764 496856
rect 43128 496816 43134 496828
rect 62758 496816 62764 496828
rect 62816 496816 62822 496868
rect 144178 496816 144184 496868
rect 144236 496856 144242 496868
rect 160646 496856 160652 496868
rect 144236 496828 160652 496856
rect 144236 496816 144242 496828
rect 160646 496816 160652 496828
rect 160704 496816 160710 496868
rect 171778 496816 171784 496868
rect 171836 496856 171842 496868
rect 197354 496856 197360 496868
rect 171836 496828 197360 496856
rect 171836 496816 171842 496828
rect 197354 496816 197360 496828
rect 197412 496816 197418 496868
rect 199378 496816 199384 496868
rect 199436 496856 199442 496868
rect 224310 496856 224316 496868
rect 199436 496828 224316 496856
rect 199436 496816 199442 496828
rect 224310 496816 224316 496828
rect 224368 496816 224374 496868
rect 225598 496816 225604 496868
rect 225656 496856 225662 496868
rect 251358 496856 251364 496868
rect 225656 496828 251364 496856
rect 225656 496816 225662 496828
rect 251358 496816 251364 496828
rect 251416 496816 251422 496868
rect 253198 496816 253204 496868
rect 253256 496856 253262 496868
rect 278314 496856 278320 496868
rect 253256 496828 278320 496856
rect 253256 496816 253262 496828
rect 278314 496816 278320 496828
rect 278372 496816 278378 496868
rect 279418 496816 279424 496868
rect 279476 496856 279482 496868
rect 305362 496856 305368 496868
rect 279476 496828 305368 496856
rect 279476 496816 279482 496828
rect 305362 496816 305368 496828
rect 305420 496816 305426 496868
rect 307018 496816 307024 496868
rect 307076 496856 307082 496868
rect 332318 496856 332324 496868
rect 307076 496828 332324 496856
rect 307076 496816 307082 496828
rect 332318 496816 332324 496828
rect 332376 496816 332382 496868
rect 333238 496816 333244 496868
rect 333296 496856 333302 496868
rect 359366 496856 359372 496868
rect 333296 496828 359372 496856
rect 333296 496816 333302 496828
rect 359366 496816 359372 496828
rect 359424 496816 359430 496868
rect 359550 496816 359556 496868
rect 359608 496856 359614 496868
rect 386322 496856 386328 496868
rect 359608 496828 386328 496856
rect 359608 496816 359614 496828
rect 386322 496816 386328 496828
rect 386380 496816 386386 496868
rect 387058 496816 387064 496868
rect 387116 496856 387122 496868
rect 413278 496856 413284 496868
rect 387116 496828 413284 496856
rect 387116 496816 387122 496828
rect 413278 496816 413284 496828
rect 413336 496816 413342 496868
rect 414658 496816 414664 496868
rect 414716 496856 414722 496868
rect 440326 496856 440332 496868
rect 414716 496828 440332 496856
rect 414716 496816 414722 496828
rect 440326 496816 440332 496828
rect 440384 496816 440390 496868
rect 442258 496816 442264 496868
rect 442316 496856 442322 496868
rect 467282 496856 467288 496868
rect 442316 496828 467288 496856
rect 442316 496816 442322 496828
rect 467282 496816 467288 496828
rect 467340 496816 467346 496868
rect 468478 496816 468484 496868
rect 468536 496856 468542 496868
rect 494330 496856 494336 496868
rect 468536 496828 494336 496856
rect 468536 496816 468542 496828
rect 494330 496816 494336 496828
rect 494388 496816 494394 496868
rect 496078 496816 496084 496868
rect 496136 496856 496142 496868
rect 521286 496856 521292 496868
rect 496136 496828 521292 496856
rect 496136 496816 496142 496828
rect 521286 496816 521292 496828
rect 521344 496816 521350 496868
rect 522298 496816 522304 496868
rect 522356 496856 522362 496868
rect 548334 496856 548340 496868
rect 522356 496828 548340 496856
rect 522356 496816 522362 496828
rect 548334 496816 548340 496828
rect 548392 496816 548398 496868
rect 37918 494708 37924 494760
rect 37976 494748 37982 494760
rect 526438 494748 526444 494760
rect 37976 494720 526444 494748
rect 37976 494708 37982 494720
rect 526438 494708 526444 494720
rect 526496 494708 526502 494760
rect 68922 494096 68928 494148
rect 68980 494136 68986 494148
rect 118694 494136 118700 494148
rect 68980 494108 118700 494136
rect 68980 494096 68986 494108
rect 118694 494096 118700 494108
rect 118752 494096 118758 494148
rect 122742 494096 122748 494148
rect 122800 494136 122806 494148
rect 172514 494136 172520 494148
rect 122800 494108 172520 494136
rect 122800 494096 122806 494108
rect 172514 494096 172520 494108
rect 172572 494096 172578 494148
rect 230382 494096 230388 494148
rect 230440 494136 230446 494148
rect 280154 494136 280160 494148
rect 230440 494108 280160 494136
rect 230440 494096 230446 494108
rect 280154 494096 280160 494108
rect 280212 494096 280218 494148
rect 311802 494096 311808 494148
rect 311860 494136 311866 494148
rect 361574 494136 361580 494148
rect 311860 494108 361580 494136
rect 311860 494096 311866 494108
rect 361574 494096 361580 494108
rect 361632 494096 361638 494148
rect 500862 494096 500868 494148
rect 500920 494136 500926 494148
rect 550634 494136 550640 494148
rect 500920 494108 550640 494136
rect 500920 494096 500926 494108
rect 550634 494096 550640 494108
rect 550692 494096 550698 494148
rect 41322 494028 41328 494080
rect 41380 494068 41386 494080
rect 91094 494068 91100 494080
rect 41380 494040 91100 494068
rect 41380 494028 41386 494040
rect 91094 494028 91100 494040
rect 91152 494028 91158 494080
rect 148962 494028 148968 494080
rect 149020 494068 149026 494080
rect 200114 494068 200120 494080
rect 149020 494040 200120 494068
rect 149020 494028 149026 494040
rect 200114 494028 200120 494040
rect 200172 494028 200178 494080
rect 202782 494028 202788 494080
rect 202840 494068 202846 494080
rect 253934 494068 253940 494080
rect 202840 494040 253940 494068
rect 202840 494028 202846 494040
rect 253934 494028 253940 494040
rect 253992 494028 253998 494080
rect 284202 494028 284208 494080
rect 284260 494068 284266 494080
rect 335354 494068 335360 494080
rect 284260 494040 335360 494068
rect 284260 494028 284266 494040
rect 335354 494028 335360 494040
rect 335412 494028 335418 494080
rect 365622 494028 365628 494080
rect 365680 494068 365686 494080
rect 415394 494068 415400 494080
rect 365680 494040 415400 494068
rect 365680 494028 365686 494040
rect 415394 494028 415400 494040
rect 415452 494028 415458 494080
rect 419442 494028 419448 494080
rect 419500 494068 419506 494080
rect 469214 494068 469220 494080
rect 419500 494040 469220 494068
rect 419500 494028 419506 494040
rect 469214 494028 469220 494040
rect 469272 494028 469278 494080
rect 473262 494028 473268 494080
rect 473320 494068 473326 494080
rect 523034 494068 523040 494080
rect 473320 494040 523040 494068
rect 473320 494028 473326 494040
rect 523034 494028 523040 494040
rect 523092 494028 523098 494080
rect 521746 477640 521752 477692
rect 521804 477680 521810 477692
rect 522390 477680 522396 477692
rect 521804 477652 522396 477680
rect 521804 477640 521810 477652
rect 522390 477640 522396 477652
rect 522448 477640 522454 477692
rect 13722 476008 13728 476060
rect 13780 476048 13786 476060
rect 64874 476048 64880 476060
rect 13780 476020 64880 476048
rect 13780 476008 13786 476020
rect 64874 476008 64880 476020
rect 64932 476008 64938 476060
rect 95142 476008 95148 476060
rect 95200 476048 95206 476060
rect 146294 476048 146300 476060
rect 95200 476020 146300 476048
rect 95200 476008 95206 476020
rect 146294 476008 146300 476020
rect 146352 476008 146358 476060
rect 176562 476008 176568 476060
rect 176620 476048 176626 476060
rect 226334 476048 226340 476060
rect 176620 476020 226340 476048
rect 176620 476008 176626 476020
rect 226334 476008 226340 476020
rect 226392 476008 226398 476060
rect 256602 476008 256608 476060
rect 256660 476048 256666 476060
rect 307754 476048 307760 476060
rect 256660 476020 307760 476048
rect 256660 476008 256666 476020
rect 307754 476008 307760 476020
rect 307812 476008 307818 476060
rect 332502 476008 332508 476060
rect 332560 476048 332566 476060
rect 334618 476048 334624 476060
rect 332560 476020 334624 476048
rect 332560 476008 332566 476020
rect 334618 476008 334624 476020
rect 334676 476008 334682 476060
rect 338022 476008 338028 476060
rect 338080 476048 338086 476060
rect 389174 476048 389180 476060
rect 338080 476020 389180 476048
rect 338080 476008 338086 476020
rect 389174 476008 389180 476020
rect 389232 476008 389238 476060
rect 391842 476008 391848 476060
rect 391900 476048 391906 476060
rect 442994 476048 443000 476060
rect 391900 476020 443000 476048
rect 391900 476008 391906 476020
rect 442994 476008 443000 476020
rect 443052 476008 443058 476060
rect 445662 476008 445668 476060
rect 445720 476048 445726 476060
rect 496814 476048 496820 476060
rect 445720 476020 496820 476048
rect 445720 476008 445726 476020
rect 496814 476008 496820 476020
rect 496872 476008 496878 476060
rect 35618 475940 35624 475992
rect 35676 475980 35682 475992
rect 36722 475980 36728 475992
rect 35676 475952 36728 475980
rect 35676 475940 35682 475952
rect 36722 475940 36728 475952
rect 36780 475940 36786 475992
rect 278682 475940 278688 475992
rect 278740 475980 278746 475992
rect 279510 475980 279516 475992
rect 278740 475952 279516 475980
rect 278740 475940 278746 475952
rect 279510 475940 279516 475952
rect 279568 475940 279574 475992
rect 467650 475940 467656 475992
rect 467708 475980 467714 475992
rect 468570 475980 468576 475992
rect 467708 475952 468576 475980
rect 467708 475940 467714 475952
rect 468570 475940 468576 475952
rect 468628 475940 468634 475992
rect 116210 475600 116216 475652
rect 116268 475640 116274 475652
rect 116486 475640 116492 475652
rect 116268 475612 116492 475640
rect 116268 475600 116274 475612
rect 116486 475600 116492 475612
rect 116544 475600 116550 475652
rect 170214 475600 170220 475652
rect 170272 475640 170278 475652
rect 170490 475640 170496 475652
rect 170272 475612 170496 475640
rect 170272 475600 170278 475612
rect 170490 475600 170496 475612
rect 170548 475600 170554 475652
rect 62758 473288 62764 473340
rect 62816 473328 62822 473340
rect 69750 473328 69756 473340
rect 62816 473300 69756 473328
rect 62816 473288 62822 473300
rect 69750 473288 69756 473300
rect 69808 473288 69814 473340
rect 96706 473288 96712 473340
rect 96764 473328 96770 473340
rect 96764 473300 103514 473328
rect 96764 473288 96770 473300
rect 15194 473220 15200 473272
rect 15252 473260 15258 473272
rect 42794 473260 42800 473272
rect 15252 473232 42800 473260
rect 15252 473220 15258 473232
rect 42794 473220 42800 473232
rect 42852 473220 42858 473272
rect 53098 473220 53104 473272
rect 53156 473260 53162 473272
rect 64138 473260 64144 473272
rect 53156 473232 64144 473260
rect 53156 473220 53162 473232
rect 64138 473220 64144 473232
rect 64196 473220 64202 473272
rect 69106 473220 69112 473272
rect 69164 473260 69170 473272
rect 96798 473260 96804 473272
rect 69164 473232 96804 473260
rect 69164 473220 69170 473232
rect 96798 473220 96804 473232
rect 96856 473220 96862 473272
rect 103486 473260 103514 473300
rect 200758 473288 200764 473340
rect 200816 473328 200822 473340
rect 204622 473328 204628 473340
rect 200816 473300 204628 473328
rect 200816 473288 200822 473300
rect 204622 473288 204628 473300
rect 204680 473288 204686 473340
rect 251818 473288 251824 473340
rect 251876 473328 251882 473340
rect 258718 473328 258724 473340
rect 251876 473300 258724 473328
rect 251876 473288 251882 473300
rect 258718 473288 258724 473300
rect 258776 473288 258782 473340
rect 443638 473288 443644 473340
rect 443696 473328 443702 473340
rect 447686 473328 447692 473340
rect 443696 473300 447692 473328
rect 443696 473288 443702 473300
rect 447686 473288 447692 473300
rect 447744 473288 447750 473340
rect 494698 473288 494704 473340
rect 494756 473328 494762 473340
rect 501598 473328 501604 473340
rect 494756 473300 501604 473328
rect 494756 473288 494762 473300
rect 501598 473288 501604 473300
rect 501656 473288 501662 473340
rect 123662 473260 123668 473272
rect 103486 473232 123668 473260
rect 123662 473220 123668 473232
rect 123720 473220 123726 473272
rect 149698 473220 149704 473272
rect 149756 473260 149762 473272
rect 547966 473260 547972 473272
rect 149756 473232 547972 473260
rect 149756 473220 149762 473232
rect 547966 473220 547972 473232
rect 548024 473220 548030 473272
rect 26050 473152 26056 473204
rect 26108 473192 26114 473204
rect 36814 473192 36820 473204
rect 26108 473164 36820 473192
rect 26108 473152 26114 473164
rect 36814 473152 36820 473164
rect 36872 473152 36878 473204
rect 79962 473152 79968 473204
rect 80020 473192 80026 473204
rect 90450 473192 90456 473204
rect 80020 473164 90456 473192
rect 80020 473152 80026 473164
rect 90450 473152 90456 473164
rect 90508 473152 90514 473204
rect 106550 473152 106556 473204
rect 106608 473192 106614 473204
rect 116578 473192 116584 473204
rect 106608 473164 116584 473192
rect 106608 473152 106614 473164
rect 116578 473152 116584 473164
rect 116636 473152 116642 473204
rect 133782 473152 133788 473204
rect 133840 473192 133846 473204
rect 144270 473192 144276 473204
rect 133840 473164 144276 473192
rect 133840 473152 133846 473164
rect 144270 473152 144276 473164
rect 144328 473152 144334 473204
rect 150526 473152 150532 473204
rect 150584 473192 150590 473204
rect 178126 473192 178132 473204
rect 150584 473164 178132 473192
rect 150584 473152 150590 473164
rect 178126 473152 178132 473164
rect 178184 473152 178190 473204
rect 187970 473152 187976 473204
rect 188028 473192 188034 473204
rect 199378 473192 199384 473204
rect 188028 473164 199384 473192
rect 188028 473152 188034 473164
rect 199378 473152 199384 473164
rect 199436 473152 199442 473204
rect 204346 473152 204352 473204
rect 204404 473192 204410 473204
rect 231854 473192 231860 473204
rect 204404 473164 231860 473192
rect 204404 473152 204410 473164
rect 231854 473152 231860 473164
rect 231912 473152 231918 473204
rect 242066 473152 242072 473204
rect 242124 473192 242130 473204
rect 253198 473192 253204 473204
rect 242124 473164 253204 473192
rect 242124 473152 242130 473164
rect 253198 473152 253204 473164
rect 253256 473152 253262 473204
rect 258166 473152 258172 473204
rect 258224 473192 258230 473204
rect 286134 473192 286140 473204
rect 258224 473164 286140 473192
rect 258224 473152 258230 473164
rect 286134 473152 286140 473164
rect 286192 473152 286198 473204
rect 312630 473192 312636 473204
rect 287026 473164 312636 473192
rect 122926 473084 122932 473136
rect 122984 473124 122990 473136
rect 150710 473124 150716 473136
rect 122984 473096 150716 473124
rect 122984 473084 122990 473096
rect 150710 473084 150716 473096
rect 150768 473084 150774 473136
rect 160554 473084 160560 473136
rect 160612 473124 160618 473136
rect 171778 473124 171784 473136
rect 160612 473096 171784 473124
rect 160612 473084 160618 473096
rect 171778 473084 171784 473096
rect 171836 473084 171842 473136
rect 215018 473084 215024 473136
rect 215076 473124 215082 473136
rect 225598 473124 225604 473136
rect 215076 473096 225604 473124
rect 215076 473084 215082 473096
rect 225598 473084 225604 473096
rect 225656 473084 225662 473136
rect 268930 473084 268936 473136
rect 268988 473124 268994 473136
rect 279418 473124 279424 473136
rect 268988 473096 279424 473124
rect 268988 473084 268994 473096
rect 279418 473084 279424 473096
rect 279476 473084 279482 473136
rect 285766 473084 285772 473136
rect 285824 473124 285830 473136
rect 287026 473124 287054 473164
rect 312630 473152 312636 473164
rect 312688 473152 312694 473204
rect 340138 473192 340144 473204
rect 316006 473164 340144 473192
rect 285824 473096 287054 473124
rect 285824 473084 285830 473096
rect 295978 473084 295984 473136
rect 296036 473124 296042 473136
rect 307018 473124 307024 473136
rect 296036 473096 307024 473124
rect 296036 473084 296042 473096
rect 307018 473084 307024 473096
rect 307076 473084 307082 473136
rect 311986 473084 311992 473136
rect 312044 473124 312050 473136
rect 316006 473124 316034 473164
rect 340138 473152 340144 473164
rect 340196 473152 340202 473204
rect 366726 473192 366732 473204
rect 344986 473164 366732 473192
rect 312044 473096 316034 473124
rect 312044 473084 312050 473096
rect 322842 473084 322848 473136
rect 322900 473124 322906 473136
rect 333238 473124 333244 473136
rect 322900 473096 333244 473124
rect 322900 473084 322906 473096
rect 333238 473084 333244 473096
rect 333296 473084 333302 473136
rect 339586 473084 339592 473136
rect 339644 473124 339650 473136
rect 344986 473124 345014 473164
rect 366726 473152 366732 473164
rect 366784 473152 366790 473204
rect 393590 473192 393596 473204
rect 373966 473164 393596 473192
rect 339644 473096 345014 473124
rect 339644 473084 339650 473096
rect 350074 473084 350080 473136
rect 350132 473124 350138 473136
rect 359550 473124 359556 473136
rect 350132 473096 359556 473124
rect 350132 473084 350138 473096
rect 359550 473084 359556 473096
rect 359608 473084 359614 473136
rect 365806 473084 365812 473136
rect 365864 473124 365870 473136
rect 373966 473124 373994 473164
rect 393590 473152 393596 473164
rect 393648 473152 393654 473204
rect 420914 473192 420920 473204
rect 402946 473164 420920 473192
rect 365864 473096 373994 473124
rect 365864 473084 365870 473096
rect 376570 473084 376576 473136
rect 376628 473124 376634 473136
rect 387058 473124 387064 473136
rect 376628 473096 387064 473124
rect 376628 473084 376634 473096
rect 387058 473084 387064 473096
rect 387116 473084 387122 473136
rect 393406 473084 393412 473136
rect 393464 473124 393470 473136
rect 402946 473124 402974 473164
rect 420914 473152 420920 473164
rect 420972 473152 420978 473204
rect 431034 473152 431040 473204
rect 431092 473192 431098 473204
rect 442258 473192 442264 473204
rect 431092 473164 442264 473192
rect 431092 473152 431098 473164
rect 442258 473152 442264 473164
rect 442316 473152 442322 473204
rect 447226 473152 447232 473204
rect 447284 473192 447290 473204
rect 474734 473192 474740 473204
rect 447284 473164 474740 473192
rect 447284 473152 447290 473164
rect 474734 473152 474740 473164
rect 474792 473152 474798 473204
rect 484946 473152 484952 473204
rect 485004 473192 485010 473204
rect 496078 473192 496084 473204
rect 485004 473164 496084 473192
rect 485004 473152 485010 473164
rect 496078 473152 496084 473164
rect 496136 473152 496142 473204
rect 501046 473152 501052 473204
rect 501104 473192 501110 473204
rect 528646 473192 528652 473204
rect 501104 473164 528652 473192
rect 501104 473152 501110 473164
rect 528646 473152 528652 473164
rect 528704 473152 528710 473204
rect 393464 473096 402974 473124
rect 393464 473084 393470 473096
rect 403986 473084 403992 473136
rect 404044 473124 404050 473136
rect 414658 473124 414664 473136
rect 404044 473096 414664 473124
rect 404044 473084 404050 473096
rect 414658 473084 414664 473096
rect 414716 473084 414722 473136
rect 458082 473084 458088 473136
rect 458140 473124 458146 473136
rect 468478 473124 468484 473136
rect 458140 473096 468484 473124
rect 458140 473084 458146 473096
rect 468478 473084 468484 473096
rect 468536 473084 468542 473136
rect 511902 473084 511908 473136
rect 511960 473124 511966 473136
rect 522298 473124 522304 473136
rect 511960 473096 522304 473124
rect 511960 473084 511966 473096
rect 522298 473084 522304 473096
rect 522356 473084 522362 473136
rect 36630 473016 36636 473068
rect 36688 473056 36694 473068
rect 538398 473056 538404 473068
rect 36688 473028 538404 473056
rect 36688 473016 36694 473028
rect 538398 473016 538404 473028
rect 538456 473016 538462 473068
rect 15286 469820 15292 469872
rect 15344 469860 15350 469872
rect 528738 469860 528744 469872
rect 15344 469832 528744 469860
rect 15344 469820 15350 469832
rect 528738 469820 528744 469832
rect 528796 469820 528802 469872
rect 25958 469480 25964 469532
rect 26016 469520 26022 469532
rect 149698 469520 149704 469532
rect 26016 469492 149704 469520
rect 26016 469480 26022 469492
rect 149698 469480 149704 469492
rect 149756 469480 149762 469532
rect 35710 469412 35716 469464
rect 35768 469452 35774 469464
rect 52454 469452 52460 469464
rect 35768 469424 52460 469452
rect 35768 469412 35774 469424
rect 52454 469412 52460 469424
rect 52512 469412 52518 469464
rect 232314 469412 232320 469464
rect 232372 469452 232378 469464
rect 251818 469452 251824 469464
rect 232372 469424 251824 469452
rect 232372 469412 232378 469424
rect 251818 469412 251824 469424
rect 251876 469412 251882 469464
rect 62482 469344 62488 469396
rect 62540 469384 62546 469396
rect 79318 469384 79324 469396
rect 62540 469356 79324 469384
rect 62540 469344 62546 469356
rect 79318 469344 79324 469356
rect 79376 469344 79382 469396
rect 90450 469344 90456 469396
rect 90508 469384 90514 469396
rect 106366 469384 106372 469396
rect 90508 469356 106372 469384
rect 90508 469344 90514 469356
rect 106366 469344 106372 469356
rect 106424 469344 106430 469396
rect 116486 469344 116492 469396
rect 116544 469384 116550 469396
rect 133414 469384 133420 469396
rect 116544 469356 133420 469384
rect 116544 469344 116550 469356
rect 133414 469344 133420 469356
rect 133472 469344 133478 469396
rect 144270 469344 144276 469396
rect 144328 469384 144334 469396
rect 160278 469384 160284 469396
rect 144328 469356 160284 469384
rect 144328 469344 144334 469356
rect 160278 469344 160284 469356
rect 160336 469344 160342 469396
rect 170490 469344 170496 469396
rect 170548 469384 170554 469396
rect 187786 469384 187792 469396
rect 170548 469356 187792 469384
rect 170548 469344 170554 469356
rect 187786 469344 187792 469356
rect 187844 469344 187850 469396
rect 197538 469344 197544 469396
rect 197596 469384 197602 469396
rect 214374 469384 214380 469396
rect 197596 469356 214380 469384
rect 197596 469344 197602 469356
rect 214374 469344 214380 469356
rect 214432 469344 214438 469396
rect 224494 469344 224500 469396
rect 224552 469384 224558 469396
rect 241514 469384 241520 469396
rect 224552 469356 241520 469384
rect 224552 469344 224558 469356
rect 241514 469344 241520 469356
rect 241572 469344 241578 469396
rect 413462 469344 413468 469396
rect 413520 469384 413526 469396
rect 430574 469384 430580 469396
rect 413520 469356 430580 469384
rect 413520 469344 413526 469356
rect 430574 469344 430580 469356
rect 430632 469344 430638 469396
rect 440510 469344 440516 469396
rect 440568 469384 440574 469396
rect 457254 469384 457260 469396
rect 440568 469356 457260 469384
rect 440568 469344 440574 469356
rect 457254 469344 457260 469356
rect 457312 469344 457318 469396
rect 36722 469276 36728 469328
rect 36780 469316 36786 469328
rect 62114 469316 62120 469328
rect 36780 469288 62120 469316
rect 36780 469276 36786 469288
rect 62114 469276 62120 469288
rect 62172 469276 62178 469328
rect 64138 469276 64144 469328
rect 64196 469316 64202 469328
rect 89070 469316 89076 469328
rect 64196 469288 89076 469316
rect 64196 469276 64202 469288
rect 89070 469276 89076 469288
rect 89128 469276 89134 469328
rect 90358 469276 90364 469328
rect 90416 469316 90422 469328
rect 115934 469316 115940 469328
rect 90416 469288 115940 469316
rect 90416 469276 90422 469288
rect 115934 469276 115940 469288
rect 115992 469276 115998 469328
rect 116578 469276 116584 469328
rect 116636 469316 116642 469328
rect 142982 469316 142988 469328
rect 116636 469288 142988 469316
rect 116636 469276 116642 469288
rect 142982 469276 142988 469288
rect 143040 469276 143046 469328
rect 144178 469276 144184 469328
rect 144236 469316 144242 469328
rect 170030 469316 170036 469328
rect 144236 469288 170036 469316
rect 144236 469276 144242 469288
rect 170030 469276 170036 469288
rect 170088 469276 170094 469328
rect 178402 469276 178408 469328
rect 178460 469316 178466 469328
rect 200758 469316 200764 469328
rect 178460 469288 200764 469316
rect 178460 469276 178466 469288
rect 200758 469276 200764 469288
rect 200816 469276 200822 469328
rect 251450 469276 251456 469328
rect 251508 469316 251514 469328
rect 268286 469316 268292 469328
rect 251508 469288 268292 469316
rect 251508 469276 251514 469288
rect 268286 469276 268292 469288
rect 268344 469276 268350 469328
rect 279510 469276 279516 469328
rect 279568 469316 279574 469328
rect 295794 469316 295800 469328
rect 279568 469288 295800 469316
rect 279568 469276 279574 469288
rect 295794 469276 295800 469288
rect 295852 469276 295858 469328
rect 305546 469276 305552 469328
rect 305604 469316 305610 469328
rect 322382 469316 322388 469328
rect 305604 469288 322388 469316
rect 305604 469276 305610 469288
rect 322382 469276 322388 469288
rect 322440 469276 322446 469328
rect 335998 469276 336004 469328
rect 336056 469316 336062 469328
rect 349798 469316 349804 469328
rect 336056 469288 349804 469316
rect 336056 469276 336062 469288
rect 349798 469276 349804 469288
rect 349856 469276 349862 469328
rect 359550 469276 359556 469328
rect 359608 469316 359614 469328
rect 376294 469316 376300 469328
rect 359608 469288 376300 469316
rect 359608 469276 359614 469288
rect 376294 469276 376300 469288
rect 376352 469276 376358 469328
rect 386506 469276 386512 469328
rect 386564 469316 386570 469328
rect 403342 469316 403348 469328
rect 386564 469288 403348 469316
rect 386564 469276 386570 469288
rect 403342 469276 403348 469288
rect 403400 469276 403406 469328
rect 421282 469276 421288 469328
rect 421340 469316 421346 469328
rect 446398 469316 446404 469328
rect 421340 469288 446404 469316
rect 421340 469276 421346 469288
rect 446398 469276 446404 469288
rect 446456 469276 446462 469328
rect 467466 469276 467472 469328
rect 467524 469316 467530 469328
rect 484394 469316 484400 469328
rect 467524 469288 484400 469316
rect 467524 469276 467530 469288
rect 484394 469276 484400 469288
rect 484452 469276 484458 469328
rect 494514 469276 494520 469328
rect 494572 469316 494578 469328
rect 511350 469316 511356 469328
rect 494572 469288 511356 469316
rect 494572 469276 494578 469288
rect 511350 469276 511356 469288
rect 511408 469276 511414 469328
rect 522298 469276 522304 469328
rect 522356 469316 522362 469328
rect 538398 469316 538404 469328
rect 522356 469288 538404 469316
rect 522356 469276 522362 469288
rect 538398 469276 538404 469288
rect 538456 469276 538462 469328
rect 43346 469208 43352 469260
rect 43404 469248 43410 469260
rect 62758 469248 62764 469260
rect 43404 469220 62764 469248
rect 43404 469208 43410 469220
rect 62758 469208 62764 469220
rect 62816 469208 62822 469260
rect 171778 469208 171784 469260
rect 171836 469248 171842 469260
rect 197446 469248 197452 469260
rect 171836 469220 197452 469248
rect 171836 469208 171842 469220
rect 197446 469208 197452 469220
rect 197504 469208 197510 469260
rect 199378 469208 199384 469260
rect 199436 469248 199442 469260
rect 223942 469248 223948 469260
rect 199436 469220 223948 469248
rect 199436 469208 199442 469220
rect 223942 469208 223948 469220
rect 224000 469208 224006 469260
rect 225598 469208 225604 469260
rect 225656 469248 225662 469260
rect 251174 469248 251180 469260
rect 225656 469220 251180 469248
rect 225656 469208 225662 469220
rect 251174 469208 251180 469220
rect 251232 469208 251238 469260
rect 253198 469208 253204 469260
rect 253256 469248 253262 469260
rect 278038 469248 278044 469260
rect 253256 469220 278044 469248
rect 253256 469208 253262 469220
rect 278038 469208 278044 469220
rect 278096 469208 278102 469260
rect 279418 469208 279424 469260
rect 279476 469248 279482 469260
rect 305454 469248 305460 469260
rect 279476 469220 305460 469248
rect 279476 469208 279482 469220
rect 305454 469208 305460 469220
rect 305512 469208 305518 469260
rect 307018 469208 307024 469260
rect 307076 469248 307082 469260
rect 331950 469248 331956 469260
rect 307076 469220 331956 469248
rect 307076 469208 307082 469220
rect 331950 469208 331956 469220
rect 332008 469208 332014 469260
rect 333238 469208 333244 469260
rect 333296 469248 333302 469260
rect 359458 469248 359464 469260
rect 333296 469220 359464 469248
rect 333296 469208 333302 469220
rect 359458 469208 359464 469220
rect 359516 469208 359522 469260
rect 359734 469208 359740 469260
rect 359792 469248 359798 469260
rect 386046 469248 386052 469260
rect 359792 469220 386052 469248
rect 359792 469208 359798 469220
rect 386046 469208 386052 469220
rect 386104 469208 386110 469260
rect 387058 469208 387064 469260
rect 387116 469248 387122 469260
rect 412910 469248 412916 469260
rect 387116 469220 412916 469248
rect 387116 469208 387122 469220
rect 412910 469208 412916 469220
rect 412968 469208 412974 469260
rect 414658 469208 414664 469260
rect 414716 469248 414722 469260
rect 440234 469248 440240 469260
rect 414716 469220 440240 469248
rect 414716 469208 414722 469220
rect 440234 469208 440240 469220
rect 440292 469208 440298 469260
rect 442258 469208 442264 469260
rect 442316 469248 442322 469260
rect 467006 469248 467012 469260
rect 442316 469220 467012 469248
rect 442316 469208 442322 469220
rect 467006 469208 467012 469220
rect 467064 469208 467070 469260
rect 468478 469208 468484 469260
rect 468536 469248 468542 469260
rect 494054 469248 494060 469260
rect 468536 469220 494060 469248
rect 468536 469208 468542 469220
rect 494054 469208 494060 469220
rect 494112 469208 494118 469260
rect 496078 469208 496084 469260
rect 496136 469248 496142 469260
rect 520918 469248 520924 469260
rect 496136 469220 520924 469248
rect 496136 469208 496142 469220
rect 520918 469208 520924 469220
rect 520976 469208 520982 469260
rect 522390 469208 522396 469260
rect 522448 469248 522454 469260
rect 548058 469248 548064 469260
rect 522448 469220 548064 469248
rect 522448 469208 522454 469220
rect 548058 469208 548064 469220
rect 548116 469208 548122 469260
rect 37918 468460 37924 468512
rect 37976 468500 37982 468512
rect 526438 468500 526444 468512
rect 37976 468472 526444 468500
rect 37976 468460 37982 468472
rect 526438 468460 526444 468472
rect 526496 468460 526502 468512
rect 339586 467304 339592 467356
rect 339644 467344 339650 467356
rect 340138 467344 340144 467356
rect 339644 467316 340144 467344
rect 339644 467304 339650 467316
rect 340138 467304 340144 467316
rect 340196 467304 340202 467356
rect 68922 466556 68928 466608
rect 68980 466596 68986 466608
rect 118694 466596 118700 466608
rect 68980 466568 118700 466596
rect 68980 466556 68986 466568
rect 118694 466556 118700 466568
rect 118752 466556 118758 466608
rect 230382 466556 230388 466608
rect 230440 466596 230446 466608
rect 280154 466596 280160 466608
rect 230440 466568 280160 466596
rect 230440 466556 230446 466568
rect 280154 466556 280160 466568
rect 280212 466556 280218 466608
rect 35618 466488 35624 466540
rect 35676 466528 35682 466540
rect 36630 466528 36636 466540
rect 35676 466500 36636 466528
rect 35676 466488 35682 466500
rect 36630 466488 36636 466500
rect 36688 466488 36694 466540
rect 41322 466488 41328 466540
rect 41380 466528 41386 466540
rect 91094 466528 91100 466540
rect 41380 466500 91100 466528
rect 41380 466488 41386 466500
rect 91094 466488 91100 466500
rect 91152 466488 91158 466540
rect 122742 466488 122748 466540
rect 122800 466528 122806 466540
rect 172514 466528 172520 466540
rect 122800 466500 172520 466528
rect 122800 466488 122806 466500
rect 172514 466488 172520 466500
rect 172572 466488 172578 466540
rect 176562 466488 176568 466540
rect 176620 466528 176626 466540
rect 226334 466528 226340 466540
rect 176620 466500 226340 466528
rect 176620 466488 176626 466500
rect 226334 466488 226340 466500
rect 226392 466488 226398 466540
rect 256602 466488 256608 466540
rect 256660 466528 256666 466540
rect 307754 466528 307760 466540
rect 256660 466500 307760 466528
rect 256660 466488 256666 466500
rect 307754 466488 307760 466500
rect 307812 466488 307818 466540
rect 311802 466488 311808 466540
rect 311860 466528 311866 466540
rect 361574 466528 361580 466540
rect 311860 466500 361580 466528
rect 311860 466488 311866 466500
rect 361574 466488 361580 466500
rect 361632 466488 361638 466540
rect 365622 466488 365628 466540
rect 365680 466528 365686 466540
rect 415394 466528 415400 466540
rect 365680 466500 415400 466528
rect 365680 466488 365686 466500
rect 415394 466488 415400 466500
rect 415452 466488 415458 466540
rect 419442 466488 419448 466540
rect 419500 466528 419506 466540
rect 469214 466528 469220 466540
rect 419500 466500 469220 466528
rect 419500 466488 419506 466500
rect 469214 466488 469220 466500
rect 469272 466488 469278 466540
rect 473262 466488 473268 466540
rect 473320 466528 473326 466540
rect 523034 466528 523040 466540
rect 473320 466500 523040 466528
rect 473320 466488 473326 466500
rect 523034 466488 523040 466500
rect 523092 466488 523098 466540
rect 13722 466420 13728 466472
rect 13780 466460 13786 466472
rect 64874 466460 64880 466472
rect 13780 466432 64880 466460
rect 13780 466420 13786 466432
rect 64874 466420 64880 466432
rect 64932 466420 64938 466472
rect 95142 466420 95148 466472
rect 95200 466460 95206 466472
rect 146294 466460 146300 466472
rect 95200 466432 146300 466460
rect 95200 466420 95206 466432
rect 146294 466420 146300 466432
rect 146352 466420 146358 466472
rect 148962 466420 148968 466472
rect 149020 466460 149026 466472
rect 200114 466460 200120 466472
rect 149020 466432 200120 466460
rect 149020 466420 149026 466432
rect 200114 466420 200120 466432
rect 200172 466420 200178 466472
rect 202782 466420 202788 466472
rect 202840 466460 202846 466472
rect 253934 466460 253940 466472
rect 202840 466432 253940 466460
rect 202840 466420 202846 466432
rect 253934 466420 253940 466432
rect 253992 466420 253998 466472
rect 284202 466420 284208 466472
rect 284260 466460 284266 466472
rect 335354 466460 335360 466472
rect 284260 466432 335360 466460
rect 284260 466420 284266 466432
rect 335354 466420 335360 466432
rect 335412 466420 335418 466472
rect 338022 466420 338028 466472
rect 338080 466460 338086 466472
rect 389174 466460 389180 466472
rect 338080 466432 389180 466460
rect 338080 466420 338086 466432
rect 389174 466420 389180 466432
rect 389232 466420 389238 466472
rect 391842 466420 391848 466472
rect 391900 466460 391906 466472
rect 442994 466460 443000 466472
rect 391900 466432 443000 466460
rect 391900 466420 391906 466432
rect 442994 466420 443000 466432
rect 443052 466420 443058 466472
rect 445662 466420 445668 466472
rect 445720 466460 445726 466472
rect 496814 466460 496820 466472
rect 445720 466432 496820 466460
rect 445720 466420 445726 466432
rect 496814 466420 496820 466432
rect 496872 466420 496878 466472
rect 500862 466420 500868 466472
rect 500920 466460 500926 466472
rect 550634 466460 550640 466472
rect 500920 466432 550640 466460
rect 500920 466420 500926 466432
rect 550634 466420 550640 466432
rect 550692 466420 550698 466472
rect 143626 449624 143632 449676
rect 143684 449664 143690 449676
rect 144270 449664 144276 449676
rect 143684 449636 144276 449664
rect 143684 449624 143690 449636
rect 144270 449624 144276 449636
rect 144328 449624 144334 449676
rect 89714 448468 89720 448520
rect 89772 448508 89778 448520
rect 90450 448508 90456 448520
rect 89772 448480 90456 448508
rect 89772 448468 89778 448480
rect 90450 448468 90456 448480
rect 90508 448468 90514 448520
rect 200758 448468 200764 448520
rect 200816 448508 200822 448520
rect 204622 448508 204628 448520
rect 200816 448480 204628 448508
rect 200816 448468 200822 448480
rect 204622 448468 204628 448480
rect 204680 448468 204686 448520
rect 278682 448468 278688 448520
rect 278740 448508 278746 448520
rect 279510 448508 279516 448520
rect 278740 448480 279516 448508
rect 278740 448468 278746 448480
rect 279510 448468 279516 448480
rect 279568 448468 279574 448520
rect 332594 448468 332600 448520
rect 332652 448508 332658 448520
rect 335998 448508 336004 448520
rect 332652 448480 336004 448508
rect 332652 448468 332658 448480
rect 335998 448468 336004 448480
rect 336056 448468 336062 448520
rect 446398 448468 446404 448520
rect 446456 448508 446462 448520
rect 447686 448508 447692 448520
rect 446456 448480 447692 448508
rect 446456 448468 446462 448480
rect 447686 448468 447692 448480
rect 447744 448468 447750 448520
rect 25682 445680 25688 445732
rect 25740 445720 25746 445732
rect 36722 445720 36728 445732
rect 25740 445692 36728 445720
rect 25740 445680 25746 445692
rect 36722 445680 36728 445692
rect 36780 445680 36786 445732
rect 62758 445680 62764 445732
rect 62816 445720 62822 445732
rect 70026 445720 70032 445732
rect 62816 445692 70032 445720
rect 62816 445680 62822 445692
rect 70026 445680 70032 445692
rect 70084 445680 70090 445732
rect 96706 445680 96712 445732
rect 96764 445720 96770 445732
rect 96764 445692 103514 445720
rect 96764 445680 96770 445692
rect 15194 445612 15200 445664
rect 15252 445652 15258 445664
rect 42978 445652 42984 445664
rect 15252 445624 42984 445652
rect 15252 445612 15258 445624
rect 42978 445612 42984 445624
rect 43036 445612 43042 445664
rect 52730 445612 52736 445664
rect 52788 445652 52794 445664
rect 64138 445652 64144 445664
rect 52788 445624 64144 445652
rect 52788 445612 52794 445624
rect 64138 445612 64144 445624
rect 64196 445612 64202 445664
rect 69106 445612 69112 445664
rect 69164 445652 69170 445664
rect 96982 445652 96988 445664
rect 69164 445624 96988 445652
rect 69164 445612 69170 445624
rect 96982 445612 96988 445624
rect 97040 445612 97046 445664
rect 103486 445652 103514 445692
rect 146938 445680 146944 445732
rect 146996 445720 147002 445732
rect 146996 445692 151814 445720
rect 146996 445680 147002 445692
rect 124030 445652 124036 445664
rect 103486 445624 124036 445652
rect 124030 445612 124036 445624
rect 124088 445612 124094 445664
rect 133690 445612 133696 445664
rect 133748 445652 133754 445664
rect 144178 445652 144184 445664
rect 133748 445624 144184 445652
rect 133748 445612 133754 445624
rect 144178 445612 144184 445624
rect 144236 445612 144242 445664
rect 150986 445652 150992 445664
rect 146588 445624 150992 445652
rect 79686 445544 79692 445596
rect 79744 445584 79750 445596
rect 90358 445584 90364 445596
rect 79744 445556 90364 445584
rect 79744 445544 79750 445556
rect 90358 445544 90364 445556
rect 90416 445544 90422 445596
rect 106642 445544 106648 445596
rect 106700 445584 106706 445596
rect 116578 445584 116584 445596
rect 106700 445556 116584 445584
rect 106700 445544 106706 445556
rect 116578 445544 116584 445556
rect 116636 445544 116642 445596
rect 122926 445544 122932 445596
rect 122984 445584 122990 445596
rect 146588 445584 146616 445624
rect 150986 445612 150992 445624
rect 151044 445612 151050 445664
rect 151786 445652 151814 445692
rect 251818 445680 251824 445732
rect 251876 445720 251882 445732
rect 258994 445720 259000 445732
rect 251876 445692 259000 445720
rect 251876 445680 251882 445692
rect 258994 445680 259000 445692
rect 259052 445680 259058 445732
rect 548334 445652 548340 445664
rect 151786 445624 548340 445652
rect 548334 445612 548340 445624
rect 548392 445612 548398 445664
rect 122984 445556 146616 445584
rect 122984 445544 122990 445556
rect 150526 445544 150532 445596
rect 150584 445584 150590 445596
rect 178034 445584 178040 445596
rect 150584 445556 178040 445584
rect 150584 445544 150590 445556
rect 178034 445544 178040 445556
rect 178092 445544 178098 445596
rect 187694 445544 187700 445596
rect 187752 445584 187758 445596
rect 199378 445584 199384 445596
rect 187752 445556 199384 445584
rect 187752 445544 187758 445556
rect 199378 445544 199384 445556
rect 199436 445544 199442 445596
rect 204346 445544 204352 445596
rect 204404 445584 204410 445596
rect 232038 445584 232044 445596
rect 204404 445556 232044 445584
rect 204404 445544 204410 445556
rect 232038 445544 232044 445556
rect 232096 445544 232102 445596
rect 241698 445544 241704 445596
rect 241756 445584 241762 445596
rect 253198 445584 253204 445596
rect 241756 445556 253204 445584
rect 241756 445544 241762 445556
rect 253198 445544 253204 445556
rect 253256 445544 253262 445596
rect 258166 445544 258172 445596
rect 258224 445584 258230 445596
rect 258224 445556 281764 445584
rect 258224 445544 258230 445556
rect 160646 445476 160652 445528
rect 160704 445516 160710 445528
rect 171778 445516 171784 445528
rect 160704 445488 171784 445516
rect 160704 445476 160710 445488
rect 171778 445476 171784 445488
rect 171836 445476 171842 445528
rect 214650 445476 214656 445528
rect 214708 445516 214714 445528
rect 225598 445516 225604 445528
rect 214708 445488 225604 445516
rect 214708 445476 214714 445488
rect 225598 445476 225604 445488
rect 225656 445476 225662 445528
rect 268654 445476 268660 445528
rect 268712 445516 268718 445528
rect 279418 445516 279424 445528
rect 268712 445488 279424 445516
rect 268712 445476 268718 445488
rect 279418 445476 279424 445488
rect 279476 445476 279482 445528
rect 281736 445516 281764 445556
rect 285766 445544 285772 445596
rect 285824 445584 285830 445596
rect 312998 445584 313004 445596
rect 285824 445556 313004 445584
rect 285824 445544 285830 445556
rect 312998 445544 313004 445556
rect 313056 445544 313062 445596
rect 340046 445584 340052 445596
rect 316006 445556 340052 445584
rect 286042 445516 286048 445528
rect 281736 445488 286048 445516
rect 286042 445476 286048 445488
rect 286100 445476 286106 445528
rect 295702 445476 295708 445528
rect 295760 445516 295766 445528
rect 307018 445516 307024 445528
rect 295760 445488 307024 445516
rect 295760 445476 295766 445488
rect 307018 445476 307024 445488
rect 307076 445476 307082 445528
rect 311986 445476 311992 445528
rect 312044 445516 312050 445528
rect 316006 445516 316034 445556
rect 340046 445544 340052 445556
rect 340104 445544 340110 445596
rect 344986 445556 364334 445584
rect 312044 445488 316034 445516
rect 312044 445476 312050 445488
rect 322658 445476 322664 445528
rect 322716 445516 322722 445528
rect 333238 445516 333244 445528
rect 322716 445488 333244 445516
rect 322716 445476 322722 445488
rect 333238 445476 333244 445488
rect 333296 445476 333302 445528
rect 339586 445476 339592 445528
rect 339644 445516 339650 445528
rect 344986 445516 345014 445556
rect 339644 445488 345014 445516
rect 339644 445476 339650 445488
rect 349706 445476 349712 445528
rect 349764 445516 349770 445528
rect 359550 445516 359556 445528
rect 349764 445488 359556 445516
rect 349764 445476 349770 445488
rect 359550 445476 359556 445488
rect 359608 445476 359614 445528
rect 364306 445516 364334 445556
rect 365806 445544 365812 445596
rect 365864 445584 365870 445596
rect 393958 445584 393964 445596
rect 365864 445556 393964 445584
rect 365864 445544 365870 445556
rect 393958 445544 393964 445556
rect 394016 445544 394022 445596
rect 421006 445584 421012 445596
rect 402946 445556 421012 445584
rect 367002 445516 367008 445528
rect 364306 445488 367008 445516
rect 367002 445476 367008 445488
rect 367060 445476 367066 445528
rect 376662 445476 376668 445528
rect 376720 445516 376726 445528
rect 387058 445516 387064 445528
rect 376720 445488 387064 445516
rect 376720 445476 376726 445488
rect 387058 445476 387064 445488
rect 387116 445476 387122 445528
rect 393406 445476 393412 445528
rect 393464 445516 393470 445528
rect 402946 445516 402974 445556
rect 421006 445544 421012 445556
rect 421064 445544 421070 445596
rect 430666 445544 430672 445596
rect 430724 445584 430730 445596
rect 442258 445584 442264 445596
rect 430724 445556 442264 445584
rect 430724 445544 430730 445556
rect 442258 445544 442264 445556
rect 442316 445544 442322 445596
rect 447226 445544 447232 445596
rect 447284 445584 447290 445596
rect 475010 445584 475016 445596
rect 447284 445556 475016 445584
rect 447284 445544 447290 445556
rect 475010 445544 475016 445556
rect 475068 445544 475074 445596
rect 480226 445556 499574 445584
rect 393464 445488 402974 445516
rect 393464 445476 393470 445488
rect 403710 445476 403716 445528
rect 403768 445516 403774 445528
rect 414658 445516 414664 445528
rect 403768 445488 414664 445516
rect 403768 445476 403774 445488
rect 414658 445476 414664 445488
rect 414716 445476 414722 445528
rect 457714 445476 457720 445528
rect 457772 445516 457778 445528
rect 468478 445516 468484 445528
rect 457772 445488 468484 445516
rect 457772 445476 457778 445488
rect 468478 445476 468484 445488
rect 468536 445476 468542 445528
rect 474826 445476 474832 445528
rect 474884 445516 474890 445528
rect 480226 445516 480254 445556
rect 474884 445488 480254 445516
rect 474884 445476 474890 445488
rect 484670 445476 484676 445528
rect 484728 445516 484734 445528
rect 496078 445516 496084 445528
rect 484728 445488 496084 445516
rect 484728 445476 484734 445488
rect 496078 445476 496084 445488
rect 496136 445476 496142 445528
rect 499546 445516 499574 445556
rect 501046 445544 501052 445596
rect 501104 445584 501110 445596
rect 529014 445584 529020 445596
rect 501104 445556 529020 445584
rect 501104 445544 501110 445556
rect 529014 445544 529020 445556
rect 529072 445544 529078 445596
rect 501966 445516 501972 445528
rect 499546 445488 501972 445516
rect 501966 445476 501972 445488
rect 502024 445476 502030 445528
rect 511718 445476 511724 445528
rect 511776 445516 511782 445528
rect 522390 445516 522396 445528
rect 511776 445488 522396 445516
rect 511776 445476 511782 445488
rect 522390 445476 522396 445488
rect 522448 445476 522454 445528
rect 36538 445408 36544 445460
rect 36596 445448 36602 445460
rect 538674 445448 538680 445460
rect 36596 445420 538680 445448
rect 36596 445408 36602 445420
rect 538674 445408 538680 445420
rect 538732 445408 538738 445460
rect 16022 443640 16028 443692
rect 16080 443680 16086 443692
rect 529014 443680 529020 443692
rect 16080 443652 529020 443680
rect 16080 443640 16086 443652
rect 529014 443640 529020 443652
rect 529072 443640 529078 443692
rect 25682 443232 25688 443284
rect 25740 443272 25746 443284
rect 146938 443272 146944 443284
rect 25740 443244 146944 443272
rect 25740 443232 25746 443244
rect 146938 443232 146944 443244
rect 146996 443232 147002 443284
rect 36722 443164 36728 443216
rect 36780 443204 36786 443216
rect 52638 443204 52644 443216
rect 36780 443176 52644 443204
rect 36780 443164 36786 443176
rect 52638 443164 52644 443176
rect 52696 443164 52702 443216
rect 232038 443164 232044 443216
rect 232096 443204 232102 443216
rect 251818 443204 251824 443216
rect 232096 443176 251824 443204
rect 232096 443164 232102 443176
rect 251818 443164 251824 443176
rect 251876 443164 251882 443216
rect 502058 443164 502064 443216
rect 502116 443204 502122 443216
rect 522482 443204 522488 443216
rect 502116 443176 522488 443204
rect 502116 443164 502122 443176
rect 522482 443164 522488 443176
rect 522540 443164 522546 443216
rect 62482 443096 62488 443148
rect 62540 443136 62546 443148
rect 79686 443136 79692 443148
rect 62540 443108 79692 443136
rect 62540 443096 62546 443108
rect 79686 443096 79692 443108
rect 79744 443096 79750 443148
rect 90450 443096 90456 443148
rect 90508 443136 90514 443148
rect 106642 443136 106648 443148
rect 90508 443108 106648 443136
rect 90508 443096 90514 443108
rect 106642 443096 106648 443108
rect 106700 443096 106706 443148
rect 116486 443096 116492 443148
rect 116544 443136 116550 443148
rect 133690 443136 133696 443148
rect 116544 443108 133696 443136
rect 116544 443096 116550 443108
rect 133690 443096 133696 443108
rect 133748 443096 133754 443148
rect 170490 443096 170496 443148
rect 170548 443136 170554 443148
rect 187694 443136 187700 443148
rect 170548 443108 187700 443136
rect 170548 443096 170554 443108
rect 187694 443096 187700 443108
rect 187752 443096 187758 443148
rect 197446 443096 197452 443148
rect 197504 443136 197510 443148
rect 214650 443136 214656 443148
rect 197504 443108 214656 443136
rect 197504 443096 197510 443108
rect 214650 443096 214656 443108
rect 214708 443096 214714 443148
rect 224494 443096 224500 443148
rect 224552 443136 224558 443148
rect 241698 443136 241704 443148
rect 224552 443108 241704 443136
rect 224552 443096 224558 443108
rect 241698 443096 241704 443108
rect 241756 443096 241762 443148
rect 305454 443096 305460 443148
rect 305512 443136 305518 443148
rect 322658 443136 322664 443148
rect 305512 443108 322664 443136
rect 305512 443096 305518 443108
rect 322658 443096 322664 443108
rect 322716 443096 322722 443148
rect 413462 443096 413468 443148
rect 413520 443136 413526 443148
rect 430666 443136 430672 443148
rect 413520 443108 430672 443136
rect 413520 443096 413526 443108
rect 430666 443096 430672 443108
rect 430724 443096 430730 443148
rect 440510 443096 440516 443148
rect 440568 443136 440574 443148
rect 457254 443136 457260 443148
rect 440568 443108 457260 443136
rect 440568 443096 440574 443108
rect 457254 443096 457260 443108
rect 457312 443096 457318 443148
rect 468570 443096 468576 443148
rect 468628 443136 468634 443148
rect 484670 443136 484676 443148
rect 468628 443108 484676 443136
rect 468628 443096 468634 443108
rect 484670 443096 484676 443108
rect 484728 443096 484734 443148
rect 494514 443096 494520 443148
rect 494572 443136 494578 443148
rect 511626 443136 511632 443148
rect 494572 443108 511632 443136
rect 494572 443096 494578 443108
rect 511626 443096 511632 443108
rect 511684 443096 511690 443148
rect 36814 443028 36820 443080
rect 36872 443068 36878 443080
rect 62298 443068 62304 443080
rect 36872 443040 62304 443068
rect 36872 443028 36878 443040
rect 62298 443028 62304 443040
rect 62356 443028 62362 443080
rect 64138 443028 64144 443080
rect 64196 443068 64202 443080
rect 89346 443068 89352 443080
rect 64196 443040 89352 443068
rect 64196 443028 64202 443040
rect 89346 443028 89352 443040
rect 89404 443028 89410 443080
rect 90358 443028 90364 443080
rect 90416 443068 90422 443080
rect 116302 443068 116308 443080
rect 90416 443040 116308 443068
rect 90416 443028 90422 443040
rect 116302 443028 116308 443040
rect 116360 443028 116366 443080
rect 116578 443028 116584 443080
rect 116636 443068 116642 443080
rect 143350 443068 143356 443080
rect 116636 443040 143356 443068
rect 116636 443028 116642 443040
rect 143350 443028 143356 443040
rect 143408 443028 143414 443080
rect 144270 443028 144276 443080
rect 144328 443068 144334 443080
rect 170306 443068 170312 443080
rect 144328 443040 170312 443068
rect 144328 443028 144334 443040
rect 170306 443028 170312 443040
rect 170364 443028 170370 443080
rect 178034 443028 178040 443080
rect 178092 443068 178098 443080
rect 200758 443068 200764 443080
rect 178092 443040 200764 443068
rect 178092 443028 178098 443040
rect 200758 443028 200764 443040
rect 200816 443028 200822 443080
rect 251450 443028 251456 443080
rect 251508 443068 251514 443080
rect 268654 443068 268660 443080
rect 251508 443040 268660 443068
rect 251508 443028 251514 443040
rect 268654 443028 268660 443040
rect 268712 443028 268718 443080
rect 279510 443028 279516 443080
rect 279568 443068 279574 443080
rect 295702 443068 295708 443080
rect 279568 443040 295708 443068
rect 279568 443028 279574 443040
rect 295702 443028 295708 443040
rect 295760 443028 295766 443080
rect 312998 443028 313004 443080
rect 313056 443068 313062 443080
rect 333330 443068 333336 443080
rect 313056 443040 333336 443068
rect 313056 443028 313062 443040
rect 333330 443028 333336 443040
rect 333388 443028 333394 443080
rect 334618 443028 334624 443080
rect 334676 443068 334682 443080
rect 349706 443068 349712 443080
rect 334676 443040 349712 443068
rect 334676 443028 334682 443040
rect 349706 443028 349712 443040
rect 349764 443028 349770 443080
rect 359458 443028 359464 443080
rect 359516 443068 359522 443080
rect 376662 443068 376668 443080
rect 359516 443040 376668 443068
rect 359516 443028 359522 443040
rect 376662 443028 376668 443040
rect 376720 443028 376726 443080
rect 386506 443028 386512 443080
rect 386564 443068 386570 443080
rect 403342 443068 403348 443080
rect 386564 443040 403348 443068
rect 386564 443028 386570 443040
rect 403342 443028 403348 443040
rect 403400 443028 403406 443080
rect 421006 443028 421012 443080
rect 421064 443068 421070 443080
rect 443638 443068 443644 443080
rect 421064 443040 443644 443068
rect 421064 443028 421070 443040
rect 443638 443028 443644 443040
rect 443696 443028 443702 443080
rect 475010 443028 475016 443080
rect 475068 443068 475074 443080
rect 494698 443068 494704 443080
rect 475068 443040 494704 443068
rect 475068 443028 475074 443040
rect 494698 443028 494704 443040
rect 494756 443028 494762 443080
rect 522298 443028 522304 443080
rect 522356 443068 522362 443080
rect 538674 443068 538680 443080
rect 522356 443040 538680 443068
rect 522356 443028 522362 443040
rect 538674 443028 538680 443040
rect 538732 443028 538738 443080
rect 43346 442960 43352 443012
rect 43404 443000 43410 443012
rect 62758 443000 62764 443012
rect 43404 442972 62764 443000
rect 43404 442960 43410 442972
rect 62758 442960 62764 442972
rect 62816 442960 62822 443012
rect 144178 442960 144184 443012
rect 144236 443000 144242 443012
rect 160646 443000 160652 443012
rect 144236 442972 160652 443000
rect 144236 442960 144242 442972
rect 160646 442960 160652 442972
rect 160704 442960 160710 443012
rect 171778 442960 171784 443012
rect 171836 443000 171842 443012
rect 197354 443000 197360 443012
rect 171836 442972 197360 443000
rect 171836 442960 171842 442972
rect 197354 442960 197360 442972
rect 197412 442960 197418 443012
rect 199378 442960 199384 443012
rect 199436 443000 199442 443012
rect 224310 443000 224316 443012
rect 199436 442972 224316 443000
rect 199436 442960 199442 442972
rect 224310 442960 224316 442972
rect 224368 442960 224374 443012
rect 225598 442960 225604 443012
rect 225656 443000 225662 443012
rect 251358 443000 251364 443012
rect 225656 442972 251364 443000
rect 225656 442960 225662 442972
rect 251358 442960 251364 442972
rect 251416 442960 251422 443012
rect 253198 442960 253204 443012
rect 253256 443000 253262 443012
rect 278314 443000 278320 443012
rect 253256 442972 278320 443000
rect 253256 442960 253262 442972
rect 278314 442960 278320 442972
rect 278372 442960 278378 443012
rect 279418 442960 279424 443012
rect 279476 443000 279482 443012
rect 305362 443000 305368 443012
rect 279476 442972 305368 443000
rect 279476 442960 279482 442972
rect 305362 442960 305368 442972
rect 305420 442960 305426 443012
rect 307018 442960 307024 443012
rect 307076 443000 307082 443012
rect 332318 443000 332324 443012
rect 307076 442972 332324 443000
rect 307076 442960 307082 442972
rect 332318 442960 332324 442972
rect 332376 442960 332382 443012
rect 333238 442960 333244 443012
rect 333296 443000 333302 443012
rect 359366 443000 359372 443012
rect 333296 442972 359372 443000
rect 333296 442960 333302 442972
rect 359366 442960 359372 442972
rect 359424 442960 359430 443012
rect 359550 442960 359556 443012
rect 359608 443000 359614 443012
rect 386322 443000 386328 443012
rect 359608 442972 386328 443000
rect 359608 442960 359614 442972
rect 386322 442960 386328 442972
rect 386380 442960 386386 443012
rect 387058 442960 387064 443012
rect 387116 443000 387122 443012
rect 412910 443000 412916 443012
rect 387116 442972 412916 443000
rect 387116 442960 387122 442972
rect 412910 442960 412916 442972
rect 412968 442960 412974 443012
rect 414658 442960 414664 443012
rect 414716 443000 414722 443012
rect 440326 443000 440332 443012
rect 414716 442972 440332 443000
rect 414716 442960 414722 442972
rect 440326 442960 440332 442972
rect 440384 442960 440390 443012
rect 442258 442960 442264 443012
rect 442316 443000 442322 443012
rect 467006 443000 467012 443012
rect 442316 442972 467012 443000
rect 442316 442960 442322 442972
rect 467006 442960 467012 442972
rect 467064 442960 467070 443012
rect 468478 442960 468484 443012
rect 468536 443000 468542 443012
rect 494330 443000 494336 443012
rect 468536 442972 494336 443000
rect 468536 442960 468542 442972
rect 494330 442960 494336 442972
rect 494388 442960 494394 443012
rect 496078 442960 496084 443012
rect 496136 443000 496142 443012
rect 521286 443000 521292 443012
rect 496136 442972 521292 443000
rect 496136 442960 496142 442972
rect 521286 442960 521292 442972
rect 521344 442960 521350 443012
rect 522390 442960 522396 443012
rect 522448 443000 522454 443012
rect 548334 443000 548340 443012
rect 522448 442972 548340 443000
rect 522448 442960 522454 442972
rect 548334 442960 548340 442972
rect 548392 442960 548398 443012
rect 37918 440852 37924 440904
rect 37976 440892 37982 440904
rect 526438 440892 526444 440904
rect 37976 440864 526444 440892
rect 37976 440852 37982 440864
rect 526438 440852 526444 440864
rect 526496 440852 526502 440904
rect 68922 440376 68928 440428
rect 68980 440416 68986 440428
rect 118694 440416 118700 440428
rect 68980 440388 118700 440416
rect 68980 440376 68986 440388
rect 118694 440376 118700 440388
rect 118752 440376 118758 440428
rect 311802 440376 311808 440428
rect 311860 440416 311866 440428
rect 361574 440416 361580 440428
rect 311860 440388 361580 440416
rect 311860 440376 311866 440388
rect 361574 440376 361580 440388
rect 361632 440376 361638 440428
rect 41322 440308 41328 440360
rect 41380 440348 41386 440360
rect 91094 440348 91100 440360
rect 41380 440320 91100 440348
rect 41380 440308 41386 440320
rect 91094 440308 91100 440320
rect 91152 440308 91158 440360
rect 122742 440308 122748 440360
rect 122800 440348 122806 440360
rect 172514 440348 172520 440360
rect 122800 440320 172520 440348
rect 122800 440308 122806 440320
rect 172514 440308 172520 440320
rect 172572 440308 172578 440360
rect 176562 440308 176568 440360
rect 176620 440348 176626 440360
rect 226334 440348 226340 440360
rect 176620 440320 226340 440348
rect 176620 440308 176626 440320
rect 226334 440308 226340 440320
rect 226392 440308 226398 440360
rect 230382 440308 230388 440360
rect 230440 440348 230446 440360
rect 280154 440348 280160 440360
rect 230440 440320 280160 440348
rect 230440 440308 230446 440320
rect 280154 440308 280160 440320
rect 280212 440308 280218 440360
rect 284202 440308 284208 440360
rect 284260 440348 284266 440360
rect 335354 440348 335360 440360
rect 284260 440320 335360 440348
rect 284260 440308 284266 440320
rect 335354 440308 335360 440320
rect 335412 440308 335418 440360
rect 338022 440308 338028 440360
rect 338080 440348 338086 440360
rect 338080 440320 345014 440348
rect 338080 440308 338086 440320
rect 13722 440240 13728 440292
rect 13780 440280 13786 440292
rect 64874 440280 64880 440292
rect 13780 440252 64880 440280
rect 13780 440240 13786 440252
rect 64874 440240 64880 440252
rect 64932 440240 64938 440292
rect 95142 440240 95148 440292
rect 95200 440280 95206 440292
rect 146294 440280 146300 440292
rect 95200 440252 146300 440280
rect 95200 440240 95206 440252
rect 146294 440240 146300 440252
rect 146352 440240 146358 440292
rect 148962 440240 148968 440292
rect 149020 440280 149026 440292
rect 200114 440280 200120 440292
rect 149020 440252 200120 440280
rect 149020 440240 149026 440252
rect 200114 440240 200120 440252
rect 200172 440240 200178 440292
rect 202782 440240 202788 440292
rect 202840 440280 202846 440292
rect 253934 440280 253940 440292
rect 202840 440252 253940 440280
rect 202840 440240 202846 440252
rect 253934 440240 253940 440252
rect 253992 440240 253998 440292
rect 256602 440240 256608 440292
rect 256660 440280 256666 440292
rect 307754 440280 307760 440292
rect 256660 440252 307760 440280
rect 256660 440240 256666 440252
rect 307754 440240 307760 440252
rect 307812 440240 307818 440292
rect 339586 440240 339592 440292
rect 339644 440280 339650 440292
rect 340138 440280 340144 440292
rect 339644 440252 340144 440280
rect 339644 440240 339650 440252
rect 340138 440240 340144 440252
rect 340196 440240 340202 440292
rect 344986 440280 345014 440320
rect 365622 440308 365628 440360
rect 365680 440348 365686 440360
rect 415394 440348 415400 440360
rect 365680 440320 415400 440348
rect 365680 440308 365686 440320
rect 415394 440308 415400 440320
rect 415452 440308 415458 440360
rect 419442 440308 419448 440360
rect 419500 440348 419506 440360
rect 469214 440348 469220 440360
rect 419500 440320 469220 440348
rect 419500 440308 419506 440320
rect 469214 440308 469220 440320
rect 469272 440308 469278 440360
rect 473262 440308 473268 440360
rect 473320 440348 473326 440360
rect 523034 440348 523040 440360
rect 473320 440320 523040 440348
rect 473320 440308 473326 440320
rect 523034 440308 523040 440320
rect 523092 440308 523098 440360
rect 389174 440280 389180 440292
rect 344986 440252 389180 440280
rect 389174 440240 389180 440252
rect 389232 440240 389238 440292
rect 391842 440240 391848 440292
rect 391900 440280 391906 440292
rect 442994 440280 443000 440292
rect 391900 440252 443000 440280
rect 391900 440240 391906 440252
rect 442994 440240 443000 440252
rect 443052 440240 443058 440292
rect 445662 440240 445668 440292
rect 445720 440280 445726 440292
rect 496814 440280 496820 440292
rect 445720 440252 496820 440280
rect 445720 440240 445726 440252
rect 496814 440240 496820 440252
rect 496872 440240 496878 440292
rect 500862 440240 500868 440292
rect 500920 440280 500926 440292
rect 550634 440280 550640 440292
rect 500920 440252 550640 440280
rect 500920 440240 500926 440252
rect 550634 440240 550640 440252
rect 550692 440240 550698 440292
rect 89714 423784 89720 423836
rect 89772 423824 89778 423836
rect 90450 423824 90456 423836
rect 89772 423796 90456 423824
rect 89772 423784 89778 423796
rect 90450 423784 90456 423796
rect 90508 423784 90514 423836
rect 522482 423036 522488 423088
rect 522540 423076 522546 423088
rect 528646 423076 528652 423088
rect 522540 423048 528652 423076
rect 522540 423036 522546 423048
rect 528646 423036 528652 423048
rect 528704 423036 528710 423088
rect 333330 422900 333336 422952
rect 333388 422940 333394 422952
rect 339862 422940 339868 422952
rect 333388 422912 339868 422940
rect 333388 422900 333394 422912
rect 339862 422900 339868 422912
rect 339920 422900 339926 422952
rect 35618 422220 35624 422272
rect 35676 422260 35682 422272
rect 36722 422260 36728 422272
rect 35676 422232 36728 422260
rect 35676 422220 35682 422232
rect 36722 422220 36728 422232
rect 36780 422220 36786 422272
rect 278682 421676 278688 421728
rect 278740 421716 278746 421728
rect 279510 421716 279516 421728
rect 278740 421688 279516 421716
rect 278740 421676 278746 421688
rect 279510 421676 279516 421688
rect 279568 421676 279574 421728
rect 332502 421676 332508 421728
rect 332560 421716 332566 421728
rect 334618 421716 334624 421728
rect 332560 421688 334624 421716
rect 332560 421676 332566 421688
rect 334618 421676 334624 421688
rect 334676 421676 334682 421728
rect 467650 421676 467656 421728
rect 467708 421716 467714 421728
rect 468570 421716 468576 421728
rect 467708 421688 468576 421716
rect 467708 421676 467714 421688
rect 468570 421676 468576 421688
rect 468628 421676 468634 421728
rect 170214 421608 170220 421660
rect 170272 421648 170278 421660
rect 170490 421648 170496 421660
rect 170272 421620 170496 421648
rect 170272 421608 170278 421620
rect 170490 421608 170496 421620
rect 170548 421608 170554 421660
rect 53098 419432 53104 419484
rect 53156 419472 53162 419484
rect 64138 419472 64144 419484
rect 53156 419444 64144 419472
rect 53156 419432 53162 419444
rect 64138 419432 64144 419444
rect 64196 419432 64202 419484
rect 69106 419432 69112 419484
rect 69164 419472 69170 419484
rect 69164 419444 74534 419472
rect 69164 419432 69170 419444
rect 15194 419364 15200 419416
rect 15252 419404 15258 419416
rect 42794 419404 42800 419416
rect 15252 419376 42800 419404
rect 15252 419364 15258 419376
rect 42794 419364 42800 419376
rect 42852 419364 42858 419416
rect 62758 419364 62764 419416
rect 62816 419404 62822 419416
rect 69750 419404 69756 419416
rect 62816 419376 69756 419404
rect 62816 419364 62822 419376
rect 69750 419364 69756 419376
rect 69808 419364 69814 419416
rect 74506 419404 74534 419444
rect 96706 419432 96712 419484
rect 96764 419472 96770 419484
rect 96764 419444 103514 419472
rect 96764 419432 96770 419444
rect 96798 419404 96804 419416
rect 74506 419376 96804 419404
rect 96798 419364 96804 419376
rect 96856 419364 96862 419416
rect 103486 419404 103514 419444
rect 200758 419432 200764 419484
rect 200816 419472 200822 419484
rect 204622 419472 204628 419484
rect 200816 419444 204628 419472
rect 200816 419432 200822 419444
rect 204622 419432 204628 419444
rect 204680 419432 204686 419484
rect 251818 419432 251824 419484
rect 251876 419472 251882 419484
rect 258718 419472 258724 419484
rect 251876 419444 258724 419472
rect 251876 419432 251882 419444
rect 258718 419432 258724 419444
rect 258776 419432 258782 419484
rect 443638 419432 443644 419484
rect 443696 419472 443702 419484
rect 447686 419472 447692 419484
rect 443696 419444 447692 419472
rect 443696 419432 443702 419444
rect 447686 419432 447692 419444
rect 447744 419432 447750 419484
rect 494698 419432 494704 419484
rect 494756 419472 494762 419484
rect 501598 419472 501604 419484
rect 494756 419444 501604 419472
rect 494756 419432 494762 419444
rect 501598 419432 501604 419444
rect 501656 419432 501662 419484
rect 123662 419404 123668 419416
rect 103486 419376 123668 419404
rect 123662 419364 123668 419376
rect 123720 419364 123726 419416
rect 149698 419364 149704 419416
rect 149756 419404 149762 419416
rect 547966 419404 547972 419416
rect 149756 419376 547972 419404
rect 149756 419364 149762 419376
rect 547966 419364 547972 419376
rect 548024 419364 548030 419416
rect 26050 419296 26056 419348
rect 26108 419336 26114 419348
rect 36814 419336 36820 419348
rect 26108 419308 36820 419336
rect 26108 419296 26114 419308
rect 36814 419296 36820 419308
rect 36872 419296 36878 419348
rect 79962 419296 79968 419348
rect 80020 419336 80026 419348
rect 90358 419336 90364 419348
rect 80020 419308 90364 419336
rect 80020 419296 80026 419308
rect 90358 419296 90364 419308
rect 90416 419296 90422 419348
rect 106550 419296 106556 419348
rect 106608 419336 106614 419348
rect 116578 419336 116584 419348
rect 106608 419308 116584 419336
rect 106608 419296 106614 419308
rect 116578 419296 116584 419308
rect 116636 419296 116642 419348
rect 133782 419296 133788 419348
rect 133840 419336 133846 419348
rect 144270 419336 144276 419348
rect 133840 419308 144276 419336
rect 133840 419296 133846 419308
rect 144270 419296 144276 419308
rect 144328 419296 144334 419348
rect 150526 419296 150532 419348
rect 150584 419336 150590 419348
rect 178126 419336 178132 419348
rect 150584 419308 178132 419336
rect 150584 419296 150590 419308
rect 178126 419296 178132 419308
rect 178184 419296 178190 419348
rect 187970 419296 187976 419348
rect 188028 419336 188034 419348
rect 199378 419336 199384 419348
rect 188028 419308 199384 419336
rect 188028 419296 188034 419308
rect 199378 419296 199384 419308
rect 199436 419296 199442 419348
rect 204346 419296 204352 419348
rect 204404 419336 204410 419348
rect 231854 419336 231860 419348
rect 204404 419308 231860 419336
rect 204404 419296 204410 419308
rect 231854 419296 231860 419308
rect 231912 419296 231918 419348
rect 242066 419296 242072 419348
rect 242124 419336 242130 419348
rect 253198 419336 253204 419348
rect 242124 419308 253204 419336
rect 242124 419296 242130 419308
rect 253198 419296 253204 419308
rect 253256 419296 253262 419348
rect 258166 419296 258172 419348
rect 258224 419336 258230 419348
rect 258224 419308 281764 419336
rect 258224 419296 258230 419308
rect 122926 419228 122932 419280
rect 122984 419268 122990 419280
rect 150710 419268 150716 419280
rect 122984 419240 150716 419268
rect 122984 419228 122990 419240
rect 150710 419228 150716 419240
rect 150768 419228 150774 419280
rect 160554 419228 160560 419280
rect 160612 419268 160618 419280
rect 171778 419268 171784 419280
rect 160612 419240 171784 419268
rect 160612 419228 160618 419240
rect 171778 419228 171784 419240
rect 171836 419228 171842 419280
rect 215018 419228 215024 419280
rect 215076 419268 215082 419280
rect 225598 419268 225604 419280
rect 215076 419240 225604 419268
rect 215076 419228 215082 419240
rect 225598 419228 225604 419240
rect 225656 419228 225662 419280
rect 268930 419228 268936 419280
rect 268988 419268 268994 419280
rect 279418 419268 279424 419280
rect 268988 419240 279424 419268
rect 268988 419228 268994 419240
rect 279418 419228 279424 419240
rect 279476 419228 279482 419280
rect 281736 419268 281764 419308
rect 285766 419296 285772 419348
rect 285824 419336 285830 419348
rect 312630 419336 312636 419348
rect 285824 419308 312636 419336
rect 285824 419296 285830 419308
rect 312630 419296 312636 419308
rect 312688 419296 312694 419348
rect 322842 419296 322848 419348
rect 322900 419336 322906 419348
rect 333238 419336 333244 419348
rect 322900 419308 333244 419336
rect 322900 419296 322906 419308
rect 333238 419296 333244 419308
rect 333296 419296 333302 419348
rect 339586 419296 339592 419348
rect 339644 419336 339650 419348
rect 339644 419308 364334 419336
rect 339644 419296 339650 419308
rect 286134 419268 286140 419280
rect 281736 419240 286140 419268
rect 286134 419228 286140 419240
rect 286192 419228 286198 419280
rect 295978 419228 295984 419280
rect 296036 419268 296042 419280
rect 307018 419268 307024 419280
rect 296036 419240 307024 419268
rect 296036 419228 296042 419240
rect 307018 419228 307024 419240
rect 307076 419228 307082 419280
rect 350074 419228 350080 419280
rect 350132 419268 350138 419280
rect 359550 419268 359556 419280
rect 350132 419240 359556 419268
rect 350132 419228 350138 419240
rect 359550 419228 359556 419240
rect 359608 419228 359614 419280
rect 364306 419268 364334 419308
rect 365806 419296 365812 419348
rect 365864 419336 365870 419348
rect 393590 419336 393596 419348
rect 365864 419308 393596 419336
rect 365864 419296 365870 419308
rect 393590 419296 393596 419308
rect 393648 419296 393654 419348
rect 420914 419336 420920 419348
rect 402946 419308 420920 419336
rect 366726 419268 366732 419280
rect 364306 419240 366732 419268
rect 366726 419228 366732 419240
rect 366784 419228 366790 419280
rect 376570 419228 376576 419280
rect 376628 419268 376634 419280
rect 387058 419268 387064 419280
rect 376628 419240 387064 419268
rect 376628 419228 376634 419240
rect 387058 419228 387064 419240
rect 387116 419228 387122 419280
rect 393406 419228 393412 419280
rect 393464 419268 393470 419280
rect 402946 419268 402974 419308
rect 420914 419296 420920 419308
rect 420972 419296 420978 419348
rect 431034 419296 431040 419348
rect 431092 419336 431098 419348
rect 442258 419336 442264 419348
rect 431092 419308 442264 419336
rect 431092 419296 431098 419308
rect 442258 419296 442264 419308
rect 442316 419296 442322 419348
rect 447226 419296 447232 419348
rect 447284 419336 447290 419348
rect 474734 419336 474740 419348
rect 447284 419308 474740 419336
rect 447284 419296 447290 419308
rect 474734 419296 474740 419308
rect 474792 419296 474798 419348
rect 484946 419296 484952 419348
rect 485004 419336 485010 419348
rect 496078 419336 496084 419348
rect 485004 419308 496084 419336
rect 485004 419296 485010 419308
rect 496078 419296 496084 419308
rect 496136 419296 496142 419348
rect 511902 419296 511908 419348
rect 511960 419336 511966 419348
rect 522390 419336 522396 419348
rect 511960 419308 522396 419336
rect 511960 419296 511966 419308
rect 522390 419296 522396 419308
rect 522448 419296 522454 419348
rect 393464 419240 402974 419268
rect 393464 419228 393470 419240
rect 403986 419228 403992 419280
rect 404044 419268 404050 419280
rect 414658 419268 414664 419280
rect 404044 419240 414664 419268
rect 404044 419228 404050 419240
rect 414658 419228 414664 419240
rect 414716 419228 414722 419280
rect 458082 419228 458088 419280
rect 458140 419268 458146 419280
rect 468478 419268 468484 419280
rect 458140 419240 468484 419268
rect 458140 419228 458146 419240
rect 468478 419228 468484 419240
rect 468536 419228 468542 419280
rect 36630 419160 36636 419212
rect 36688 419200 36694 419212
rect 538398 419200 538404 419212
rect 36688 419172 538404 419200
rect 36688 419160 36694 419172
rect 538398 419160 538404 419172
rect 538456 419160 538462 419212
rect 16298 416032 16304 416084
rect 16356 416072 16362 416084
rect 528738 416072 528744 416084
rect 16356 416044 528744 416072
rect 16356 416032 16362 416044
rect 528738 416032 528744 416044
rect 528796 416032 528802 416084
rect 25958 415692 25964 415744
rect 26016 415732 26022 415744
rect 149698 415732 149704 415744
rect 26016 415704 149704 415732
rect 26016 415692 26022 415704
rect 149698 415692 149704 415704
rect 149756 415692 149762 415744
rect 36722 415624 36728 415676
rect 36780 415664 36786 415676
rect 52454 415664 52460 415676
rect 36780 415636 52460 415664
rect 36780 415624 36786 415636
rect 52454 415624 52460 415636
rect 52512 415624 52518 415676
rect 475378 415624 475384 415676
rect 475436 415664 475442 415676
rect 494698 415664 494704 415676
rect 475436 415636 494704 415664
rect 475436 415624 475442 415636
rect 494698 415624 494704 415636
rect 494756 415624 494762 415676
rect 43346 415556 43352 415608
rect 43404 415596 43410 415608
rect 62758 415596 62764 415608
rect 43404 415568 62764 415596
rect 43404 415556 43410 415568
rect 62758 415556 62764 415568
rect 62816 415556 62822 415608
rect 90450 415556 90456 415608
rect 90508 415596 90514 415608
rect 106366 415596 106372 415608
rect 90508 415568 106372 415596
rect 90508 415556 90514 415568
rect 106366 415556 106372 415568
rect 106424 415556 106430 415608
rect 116486 415556 116492 415608
rect 116544 415596 116550 415608
rect 133414 415596 133420 415608
rect 116544 415568 133420 415596
rect 116544 415556 116550 415568
rect 133414 415556 133420 415568
rect 133472 415556 133478 415608
rect 144270 415556 144276 415608
rect 144328 415596 144334 415608
rect 160278 415596 160284 415608
rect 144328 415568 160284 415596
rect 144328 415556 144334 415568
rect 160278 415556 160284 415568
rect 160336 415556 160342 415608
rect 170490 415556 170496 415608
rect 170548 415596 170554 415608
rect 187786 415596 187792 415608
rect 170548 415568 187792 415596
rect 170548 415556 170554 415568
rect 187786 415556 187792 415568
rect 187844 415556 187850 415608
rect 197538 415556 197544 415608
rect 197596 415596 197602 415608
rect 214374 415596 214380 415608
rect 197596 415568 214380 415596
rect 197596 415556 197602 415568
rect 214374 415556 214380 415568
rect 214432 415556 214438 415608
rect 224494 415556 224500 415608
rect 224552 415596 224558 415608
rect 241514 415596 241520 415608
rect 224552 415568 241520 415596
rect 224552 415556 224558 415568
rect 241514 415556 241520 415568
rect 241572 415556 241578 415608
rect 251450 415556 251456 415608
rect 251508 415596 251514 415608
rect 268286 415596 268292 415608
rect 251508 415568 268292 415596
rect 251508 415556 251514 415568
rect 268286 415556 268292 415568
rect 268344 415556 268350 415608
rect 413462 415556 413468 415608
rect 413520 415596 413526 415608
rect 430574 415596 430580 415608
rect 413520 415568 430580 415596
rect 413520 415556 413526 415568
rect 430574 415556 430580 415568
rect 430632 415556 430638 415608
rect 440510 415556 440516 415608
rect 440568 415596 440574 415608
rect 457254 415596 457260 415608
rect 440568 415568 457260 415596
rect 440568 415556 440574 415568
rect 457254 415556 457260 415568
rect 457312 415556 457318 415608
rect 468570 415556 468576 415608
rect 468628 415596 468634 415608
rect 484394 415596 484400 415608
rect 468628 415568 484400 415596
rect 468628 415556 468634 415568
rect 484394 415556 484400 415568
rect 484452 415556 484458 415608
rect 36814 415488 36820 415540
rect 36872 415528 36878 415540
rect 62114 415528 62120 415540
rect 36872 415500 62120 415528
rect 36872 415488 36878 415500
rect 62114 415488 62120 415500
rect 62172 415488 62178 415540
rect 64138 415488 64144 415540
rect 64196 415528 64202 415540
rect 89070 415528 89076 415540
rect 64196 415500 89076 415528
rect 64196 415488 64202 415500
rect 89070 415488 89076 415500
rect 89128 415488 89134 415540
rect 90358 415488 90364 415540
rect 90416 415528 90422 415540
rect 115934 415528 115940 415540
rect 90416 415500 115940 415528
rect 90416 415488 90422 415500
rect 115934 415488 115940 415500
rect 115992 415488 115998 415540
rect 116578 415488 116584 415540
rect 116636 415528 116642 415540
rect 142982 415528 142988 415540
rect 116636 415500 142988 415528
rect 116636 415488 116642 415500
rect 142982 415488 142988 415500
rect 143040 415488 143046 415540
rect 144178 415488 144184 415540
rect 144236 415528 144242 415540
rect 170030 415528 170036 415540
rect 144236 415500 170036 415528
rect 144236 415488 144242 415500
rect 170030 415488 170036 415500
rect 170088 415488 170094 415540
rect 178402 415488 178408 415540
rect 178460 415528 178466 415540
rect 200758 415528 200764 415540
rect 178460 415500 200764 415528
rect 178460 415488 178466 415500
rect 200758 415488 200764 415500
rect 200816 415488 200822 415540
rect 232314 415488 232320 415540
rect 232372 415528 232378 415540
rect 251818 415528 251824 415540
rect 232372 415500 251824 415528
rect 232372 415488 232378 415500
rect 251818 415488 251824 415500
rect 251876 415488 251882 415540
rect 279510 415488 279516 415540
rect 279568 415528 279574 415540
rect 295794 415528 295800 415540
rect 279568 415500 295800 415528
rect 279568 415488 279574 415500
rect 295794 415488 295800 415500
rect 295852 415488 295858 415540
rect 305638 415488 305644 415540
rect 305696 415528 305702 415540
rect 322382 415528 322388 415540
rect 305696 415500 322388 415528
rect 305696 415488 305702 415500
rect 322382 415488 322388 415500
rect 322440 415488 322446 415540
rect 335998 415488 336004 415540
rect 336056 415528 336062 415540
rect 349798 415528 349804 415540
rect 336056 415500 349804 415528
rect 336056 415488 336062 415500
rect 349798 415488 349804 415500
rect 349856 415488 349862 415540
rect 359642 415488 359648 415540
rect 359700 415528 359706 415540
rect 376294 415528 376300 415540
rect 359700 415500 376300 415528
rect 359700 415488 359706 415500
rect 376294 415488 376300 415500
rect 376352 415488 376358 415540
rect 386506 415488 386512 415540
rect 386564 415528 386570 415540
rect 403342 415528 403348 415540
rect 386564 415500 403348 415528
rect 386564 415488 386570 415500
rect 403342 415488 403348 415500
rect 403400 415488 403406 415540
rect 421282 415488 421288 415540
rect 421340 415528 421346 415540
rect 445018 415528 445024 415540
rect 421340 415500 445024 415528
rect 421340 415488 421346 415500
rect 445018 415488 445024 415500
rect 445076 415488 445082 415540
rect 494514 415488 494520 415540
rect 494572 415528 494578 415540
rect 511350 415528 511356 415540
rect 494572 415500 511356 415528
rect 494572 415488 494578 415500
rect 511350 415488 511356 415500
rect 511408 415488 511414 415540
rect 522298 415488 522304 415540
rect 522356 415528 522362 415540
rect 538398 415528 538404 415540
rect 522356 415500 538404 415528
rect 522356 415488 522362 415500
rect 538398 415488 538404 415500
rect 538456 415488 538462 415540
rect 62482 415420 62488 415472
rect 62540 415460 62546 415472
rect 79318 415460 79324 415472
rect 62540 415432 79324 415460
rect 62540 415420 62546 415432
rect 79318 415420 79324 415432
rect 79376 415420 79382 415472
rect 171778 415420 171784 415472
rect 171836 415460 171842 415472
rect 197446 415460 197452 415472
rect 171836 415432 197452 415460
rect 171836 415420 171842 415432
rect 197446 415420 197452 415432
rect 197504 415420 197510 415472
rect 199378 415420 199384 415472
rect 199436 415460 199442 415472
rect 223942 415460 223948 415472
rect 199436 415432 223948 415460
rect 199436 415420 199442 415432
rect 223942 415420 223948 415432
rect 224000 415420 224006 415472
rect 225598 415420 225604 415472
rect 225656 415460 225662 415472
rect 251174 415460 251180 415472
rect 225656 415432 251180 415460
rect 225656 415420 225662 415432
rect 251174 415420 251180 415432
rect 251232 415420 251238 415472
rect 253198 415420 253204 415472
rect 253256 415460 253262 415472
rect 278038 415460 278044 415472
rect 253256 415432 278044 415460
rect 253256 415420 253262 415432
rect 278038 415420 278044 415432
rect 278096 415420 278102 415472
rect 279418 415420 279424 415472
rect 279476 415460 279482 415472
rect 305546 415460 305552 415472
rect 279476 415432 305552 415460
rect 279476 415420 279482 415432
rect 305546 415420 305552 415432
rect 305604 415420 305610 415472
rect 307018 415420 307024 415472
rect 307076 415460 307082 415472
rect 331950 415460 331956 415472
rect 307076 415432 331956 415460
rect 307076 415420 307082 415432
rect 331950 415420 331956 415432
rect 332008 415420 332014 415472
rect 333238 415420 333244 415472
rect 333296 415460 333302 415472
rect 359458 415460 359464 415472
rect 333296 415432 359464 415460
rect 333296 415420 333302 415432
rect 359458 415420 359464 415432
rect 359516 415420 359522 415472
rect 359734 415420 359740 415472
rect 359792 415460 359798 415472
rect 386046 415460 386052 415472
rect 359792 415432 386052 415460
rect 359792 415420 359798 415432
rect 386046 415420 386052 415432
rect 386104 415420 386110 415472
rect 387058 415420 387064 415472
rect 387116 415460 387122 415472
rect 412910 415460 412916 415472
rect 387116 415432 412916 415460
rect 387116 415420 387122 415432
rect 412910 415420 412916 415432
rect 412968 415420 412974 415472
rect 414658 415420 414664 415472
rect 414716 415460 414722 415472
rect 440234 415460 440240 415472
rect 414716 415432 440240 415460
rect 414716 415420 414722 415432
rect 440234 415420 440240 415432
rect 440292 415420 440298 415472
rect 442258 415420 442264 415472
rect 442316 415460 442322 415472
rect 467006 415460 467012 415472
rect 442316 415432 467012 415460
rect 442316 415420 442322 415432
rect 467006 415420 467012 415432
rect 467064 415420 467070 415472
rect 468478 415420 468484 415472
rect 468536 415460 468542 415472
rect 494054 415460 494060 415472
rect 468536 415432 494060 415460
rect 468536 415420 468542 415432
rect 494054 415420 494060 415432
rect 494112 415420 494118 415472
rect 496078 415420 496084 415472
rect 496136 415460 496142 415472
rect 520918 415460 520924 415472
rect 496136 415432 520924 415460
rect 496136 415420 496142 415432
rect 520918 415420 520924 415432
rect 520976 415420 520982 415472
rect 522390 415420 522396 415472
rect 522448 415460 522454 415472
rect 548058 415460 548064 415472
rect 522448 415432 548064 415460
rect 522448 415420 522454 415432
rect 548058 415420 548064 415432
rect 548116 415420 548122 415472
rect 37918 414672 37924 414724
rect 37976 414712 37982 414724
rect 526438 414712 526444 414724
rect 37976 414684 526444 414712
rect 37976 414672 37982 414684
rect 526438 414672 526444 414684
rect 526496 414672 526502 414724
rect 339586 413312 339592 413364
rect 339644 413352 339650 413364
rect 340138 413352 340144 413364
rect 339644 413324 340144 413352
rect 339644 413312 339650 413324
rect 340138 413312 340144 413324
rect 340196 413312 340202 413364
rect 35618 412632 35624 412684
rect 35676 412672 35682 412684
rect 36630 412672 36636 412684
rect 35676 412644 36636 412672
rect 35676 412632 35682 412644
rect 36630 412632 36636 412644
rect 36688 412632 36694 412684
rect 143552 394692 144408 394720
rect 13722 394612 13728 394664
rect 13780 394652 13786 394664
rect 64874 394652 64880 394664
rect 13780 394624 64880 394652
rect 13780 394612 13786 394624
rect 64874 394612 64880 394624
rect 64932 394612 64938 394664
rect 89714 394612 89720 394664
rect 89772 394652 89778 394664
rect 90450 394652 90456 394664
rect 89772 394624 90456 394652
rect 89772 394612 89778 394624
rect 90450 394612 90456 394624
rect 90508 394612 90514 394664
rect 95142 394612 95148 394664
rect 95200 394652 95206 394664
rect 143552 394652 143580 394692
rect 95200 394624 143580 394652
rect 95200 394612 95206 394624
rect 143626 394612 143632 394664
rect 143684 394652 143690 394664
rect 144270 394652 144276 394664
rect 143684 394624 144276 394652
rect 143684 394612 143690 394624
rect 144270 394612 144276 394624
rect 144328 394612 144334 394664
rect 144380 394652 144408 394692
rect 445018 394680 445024 394732
rect 445076 394720 445082 394732
rect 447686 394720 447692 394732
rect 445076 394692 447692 394720
rect 445076 394680 445082 394692
rect 447686 394680 447692 394692
rect 447744 394680 447750 394732
rect 146294 394652 146300 394664
rect 144380 394624 146300 394652
rect 146294 394612 146300 394624
rect 146352 394612 146358 394664
rect 148962 394612 148968 394664
rect 149020 394652 149026 394664
rect 200114 394652 200120 394664
rect 149020 394624 200120 394652
rect 149020 394612 149026 394624
rect 200114 394612 200120 394624
rect 200172 394612 200178 394664
rect 202782 394612 202788 394664
rect 202840 394652 202846 394664
rect 253934 394652 253940 394664
rect 202840 394624 253940 394652
rect 202840 394612 202846 394624
rect 253934 394612 253940 394624
rect 253992 394612 253998 394664
rect 278682 394612 278688 394664
rect 278740 394652 278746 394664
rect 279510 394652 279516 394664
rect 278740 394624 279516 394652
rect 278740 394612 278746 394624
rect 279510 394612 279516 394624
rect 279568 394612 279574 394664
rect 284202 394612 284208 394664
rect 284260 394652 284266 394664
rect 335354 394652 335360 394664
rect 284260 394624 335360 394652
rect 284260 394612 284266 394624
rect 335354 394612 335360 394624
rect 335412 394612 335418 394664
rect 338022 394612 338028 394664
rect 338080 394652 338086 394664
rect 389174 394652 389180 394664
rect 338080 394624 389180 394652
rect 338080 394612 338086 394624
rect 389174 394612 389180 394624
rect 389232 394612 389238 394664
rect 391842 394612 391848 394664
rect 391900 394652 391906 394664
rect 442994 394652 443000 394664
rect 391900 394624 443000 394652
rect 391900 394612 391906 394624
rect 442994 394612 443000 394624
rect 443052 394612 443058 394664
rect 445662 394612 445668 394664
rect 445720 394652 445726 394664
rect 496814 394652 496820 394664
rect 445720 394624 496820 394652
rect 445720 394612 445726 394624
rect 496814 394612 496820 394624
rect 496872 394612 496878 394664
rect 500862 394612 500868 394664
rect 500920 394652 500926 394664
rect 550634 394652 550640 394664
rect 500920 394624 550640 394652
rect 500920 394612 500926 394624
rect 550634 394612 550640 394624
rect 550692 394612 550698 394664
rect 35618 394544 35624 394596
rect 35676 394584 35682 394596
rect 36722 394584 36728 394596
rect 35676 394556 36728 394584
rect 35676 394544 35682 394556
rect 36722 394544 36728 394556
rect 36780 394544 36786 394596
rect 41322 394544 41328 394596
rect 41380 394584 41386 394596
rect 91094 394584 91100 394596
rect 41380 394556 91100 394584
rect 41380 394544 41386 394556
rect 91094 394544 91100 394556
rect 91152 394544 91158 394596
rect 122742 394544 122748 394596
rect 122800 394584 122806 394596
rect 172514 394584 172520 394596
rect 122800 394556 172520 394584
rect 122800 394544 122806 394556
rect 172514 394544 172520 394556
rect 172572 394544 172578 394596
rect 176562 394544 176568 394596
rect 176620 394584 176626 394596
rect 226334 394584 226340 394596
rect 176620 394556 226340 394584
rect 176620 394544 176626 394556
rect 226334 394544 226340 394556
rect 226392 394544 226398 394596
rect 256602 394544 256608 394596
rect 256660 394584 256666 394596
rect 307754 394584 307760 394596
rect 256660 394556 307760 394584
rect 256660 394544 256666 394556
rect 307754 394544 307760 394556
rect 307812 394544 307818 394596
rect 311802 394544 311808 394596
rect 311860 394584 311866 394596
rect 361574 394584 361580 394596
rect 311860 394556 361580 394584
rect 311860 394544 311866 394556
rect 361574 394544 361580 394556
rect 361632 394544 361638 394596
rect 365622 394544 365628 394596
rect 365680 394584 365686 394596
rect 415394 394584 415400 394596
rect 365680 394556 415400 394584
rect 365680 394544 365686 394556
rect 415394 394544 415400 394556
rect 415452 394544 415458 394596
rect 419442 394544 419448 394596
rect 419500 394584 419506 394596
rect 419500 394556 451274 394584
rect 419500 394544 419506 394556
rect 68922 394476 68928 394528
rect 68980 394516 68986 394528
rect 118694 394516 118700 394528
rect 68980 394488 118700 394516
rect 68980 394476 68986 394488
rect 118694 394476 118700 394488
rect 118752 394476 118758 394528
rect 230382 394476 230388 394528
rect 230440 394516 230446 394528
rect 280154 394516 280160 394528
rect 230440 394488 280160 394516
rect 230440 394476 230446 394488
rect 280154 394476 280160 394488
rect 280212 394476 280218 394528
rect 332594 394476 332600 394528
rect 332652 394516 332658 394528
rect 335998 394516 336004 394528
rect 332652 394488 336004 394516
rect 332652 394476 332658 394488
rect 335998 394476 336004 394488
rect 336056 394476 336062 394528
rect 451246 394516 451274 394556
rect 467650 394544 467656 394596
rect 467708 394584 467714 394596
rect 468570 394584 468576 394596
rect 467708 394556 468576 394584
rect 467708 394544 467714 394556
rect 468570 394544 468576 394556
rect 468628 394544 468634 394596
rect 473262 394544 473268 394596
rect 473320 394584 473326 394596
rect 523034 394584 523040 394596
rect 473320 394556 523040 394584
rect 473320 394544 473326 394556
rect 523034 394544 523040 394556
rect 523092 394544 523098 394596
rect 469214 394516 469220 394528
rect 451246 394488 469220 394516
rect 469214 394476 469220 394488
rect 469272 394476 469278 394528
rect 52730 391892 52736 391944
rect 52788 391932 52794 391944
rect 64138 391932 64144 391944
rect 52788 391904 64144 391932
rect 52788 391892 52794 391904
rect 64138 391892 64144 391904
rect 64196 391892 64202 391944
rect 69106 391892 69112 391944
rect 69164 391932 69170 391944
rect 69164 391904 74534 391932
rect 69164 391892 69170 391904
rect 15194 391824 15200 391876
rect 15252 391864 15258 391876
rect 42978 391864 42984 391876
rect 15252 391836 42984 391864
rect 15252 391824 15258 391836
rect 42978 391824 42984 391836
rect 43036 391824 43042 391876
rect 62758 391824 62764 391876
rect 62816 391864 62822 391876
rect 70026 391864 70032 391876
rect 62816 391836 70032 391864
rect 62816 391824 62822 391836
rect 70026 391824 70032 391836
rect 70084 391824 70090 391876
rect 74506 391864 74534 391904
rect 96706 391892 96712 391944
rect 96764 391932 96770 391944
rect 96764 391904 103514 391932
rect 96764 391892 96770 391904
rect 96982 391864 96988 391876
rect 74506 391836 96988 391864
rect 96982 391824 96988 391836
rect 97040 391824 97046 391876
rect 103486 391864 103514 391904
rect 200758 391892 200764 391944
rect 200816 391932 200822 391944
rect 204990 391932 204996 391944
rect 200816 391904 204996 391932
rect 200816 391892 200822 391904
rect 204990 391892 204996 391904
rect 205048 391892 205054 391944
rect 251818 391892 251824 391944
rect 251876 391932 251882 391944
rect 258994 391932 259000 391944
rect 251876 391904 259000 391932
rect 251876 391892 251882 391904
rect 258994 391892 259000 391904
rect 259052 391892 259058 391944
rect 494698 391892 494704 391944
rect 494756 391932 494762 391944
rect 501966 391932 501972 391944
rect 494756 391904 501972 391932
rect 494756 391892 494762 391904
rect 501966 391892 501972 391904
rect 502024 391892 502030 391944
rect 124030 391864 124036 391876
rect 103486 391836 124036 391864
rect 124030 391824 124036 391836
rect 124088 391824 124094 391876
rect 133690 391824 133696 391876
rect 133748 391864 133754 391876
rect 144178 391864 144184 391876
rect 133748 391836 144184 391864
rect 133748 391824 133754 391836
rect 144178 391824 144184 391836
rect 144236 391824 144242 391876
rect 146938 391824 146944 391876
rect 146996 391864 147002 391876
rect 548334 391864 548340 391876
rect 146996 391836 548340 391864
rect 146996 391824 147002 391836
rect 548334 391824 548340 391836
rect 548392 391824 548398 391876
rect 25682 391756 25688 391808
rect 25740 391796 25746 391808
rect 36814 391796 36820 391808
rect 25740 391768 36820 391796
rect 25740 391756 25746 391768
rect 36814 391756 36820 391768
rect 36872 391756 36878 391808
rect 79686 391756 79692 391808
rect 79744 391796 79750 391808
rect 90358 391796 90364 391808
rect 79744 391768 90364 391796
rect 79744 391756 79750 391768
rect 90358 391756 90364 391768
rect 90416 391756 90422 391808
rect 106642 391756 106648 391808
rect 106700 391796 106706 391808
rect 116578 391796 116584 391808
rect 106700 391768 116584 391796
rect 106700 391756 106706 391768
rect 116578 391756 116584 391768
rect 116636 391756 116642 391808
rect 122926 391756 122932 391808
rect 122984 391796 122990 391808
rect 122984 391768 142154 391796
rect 122984 391756 122990 391768
rect 142126 391728 142154 391768
rect 150526 391756 150532 391808
rect 150584 391796 150590 391808
rect 178034 391796 178040 391808
rect 150584 391768 178040 391796
rect 150584 391756 150590 391768
rect 178034 391756 178040 391768
rect 178092 391756 178098 391808
rect 187694 391756 187700 391808
rect 187752 391796 187758 391808
rect 199378 391796 199384 391808
rect 187752 391768 199384 391796
rect 187752 391756 187758 391768
rect 199378 391756 199384 391768
rect 199436 391756 199442 391808
rect 204346 391756 204352 391808
rect 204404 391796 204410 391808
rect 232038 391796 232044 391808
rect 204404 391768 232044 391796
rect 204404 391756 204410 391768
rect 232038 391756 232044 391768
rect 232096 391756 232102 391808
rect 241698 391756 241704 391808
rect 241756 391796 241762 391808
rect 253198 391796 253204 391808
rect 241756 391768 253204 391796
rect 241756 391756 241762 391768
rect 253198 391756 253204 391768
rect 253256 391756 253262 391808
rect 258166 391756 258172 391808
rect 258224 391796 258230 391808
rect 258224 391768 281764 391796
rect 258224 391756 258230 391768
rect 150986 391728 150992 391740
rect 142126 391700 150992 391728
rect 150986 391688 150992 391700
rect 151044 391688 151050 391740
rect 160646 391688 160652 391740
rect 160704 391728 160710 391740
rect 171778 391728 171784 391740
rect 160704 391700 171784 391728
rect 160704 391688 160710 391700
rect 171778 391688 171784 391700
rect 171836 391688 171842 391740
rect 214650 391688 214656 391740
rect 214708 391728 214714 391740
rect 225598 391728 225604 391740
rect 214708 391700 225604 391728
rect 214708 391688 214714 391700
rect 225598 391688 225604 391700
rect 225656 391688 225662 391740
rect 268654 391688 268660 391740
rect 268712 391728 268718 391740
rect 279418 391728 279424 391740
rect 268712 391700 279424 391728
rect 268712 391688 268718 391700
rect 279418 391688 279424 391700
rect 279476 391688 279482 391740
rect 281736 391728 281764 391768
rect 285766 391756 285772 391808
rect 285824 391796 285830 391808
rect 312998 391796 313004 391808
rect 285824 391768 313004 391796
rect 285824 391756 285830 391768
rect 312998 391756 313004 391768
rect 313056 391756 313062 391808
rect 340046 391796 340052 391808
rect 316006 391768 340052 391796
rect 286042 391728 286048 391740
rect 281736 391700 286048 391728
rect 286042 391688 286048 391700
rect 286100 391688 286106 391740
rect 295702 391688 295708 391740
rect 295760 391728 295766 391740
rect 307018 391728 307024 391740
rect 295760 391700 307024 391728
rect 295760 391688 295766 391700
rect 307018 391688 307024 391700
rect 307076 391688 307082 391740
rect 311986 391688 311992 391740
rect 312044 391728 312050 391740
rect 316006 391728 316034 391768
rect 340046 391756 340052 391768
rect 340104 391756 340110 391808
rect 366726 391796 366732 391808
rect 344986 391768 366732 391796
rect 312044 391700 316034 391728
rect 312044 391688 312050 391700
rect 322658 391688 322664 391740
rect 322716 391728 322722 391740
rect 333238 391728 333244 391740
rect 322716 391700 333244 391728
rect 322716 391688 322722 391700
rect 333238 391688 333244 391700
rect 333296 391688 333302 391740
rect 339586 391688 339592 391740
rect 339644 391728 339650 391740
rect 344986 391728 345014 391768
rect 366726 391756 366732 391768
rect 366784 391756 366790 391808
rect 393958 391796 393964 391808
rect 373966 391768 393964 391796
rect 339644 391700 345014 391728
rect 339644 391688 339650 391700
rect 349706 391688 349712 391740
rect 349764 391728 349770 391740
rect 359550 391728 359556 391740
rect 349764 391700 359556 391728
rect 349764 391688 349770 391700
rect 359550 391688 359556 391700
rect 359608 391688 359614 391740
rect 365806 391688 365812 391740
rect 365864 391728 365870 391740
rect 373966 391728 373994 391768
rect 393958 391756 393964 391768
rect 394016 391756 394022 391808
rect 421006 391796 421012 391808
rect 402946 391768 421012 391796
rect 365864 391700 373994 391728
rect 365864 391688 365870 391700
rect 376662 391688 376668 391740
rect 376720 391728 376726 391740
rect 387058 391728 387064 391740
rect 376720 391700 387064 391728
rect 376720 391688 376726 391700
rect 387058 391688 387064 391700
rect 387116 391688 387122 391740
rect 393406 391688 393412 391740
rect 393464 391728 393470 391740
rect 402946 391728 402974 391768
rect 421006 391756 421012 391768
rect 421064 391756 421070 391808
rect 430666 391756 430672 391808
rect 430724 391796 430730 391808
rect 442258 391796 442264 391808
rect 430724 391768 442264 391796
rect 430724 391756 430730 391768
rect 442258 391756 442264 391768
rect 442316 391756 442322 391808
rect 447226 391756 447232 391808
rect 447284 391796 447290 391808
rect 475010 391796 475016 391808
rect 447284 391768 475016 391796
rect 447284 391756 447290 391768
rect 475010 391756 475016 391768
rect 475068 391756 475074 391808
rect 484670 391756 484676 391808
rect 484728 391796 484734 391808
rect 496078 391796 496084 391808
rect 484728 391768 496084 391796
rect 484728 391756 484734 391768
rect 496078 391756 496084 391768
rect 496136 391756 496142 391808
rect 501046 391756 501052 391808
rect 501104 391796 501110 391808
rect 529014 391796 529020 391808
rect 501104 391768 529020 391796
rect 501104 391756 501110 391768
rect 529014 391756 529020 391768
rect 529072 391756 529078 391808
rect 393464 391700 402974 391728
rect 393464 391688 393470 391700
rect 403710 391688 403716 391740
rect 403768 391728 403774 391740
rect 414658 391728 414664 391740
rect 403768 391700 414664 391728
rect 403768 391688 403774 391700
rect 414658 391688 414664 391700
rect 414716 391688 414722 391740
rect 457714 391688 457720 391740
rect 457772 391728 457778 391740
rect 468478 391728 468484 391740
rect 457772 391700 468484 391728
rect 457772 391688 457778 391700
rect 468478 391688 468484 391700
rect 468536 391688 468542 391740
rect 511718 391688 511724 391740
rect 511776 391728 511782 391740
rect 522390 391728 522396 391740
rect 511776 391700 522396 391728
rect 511776 391688 511782 391700
rect 522390 391688 522396 391700
rect 522448 391688 522454 391740
rect 36538 391620 36544 391672
rect 36596 391660 36602 391672
rect 538674 391660 538680 391672
rect 36596 391632 538680 391660
rect 36596 391620 36602 391632
rect 538674 391620 538680 391632
rect 538732 391620 538738 391672
rect 16022 389784 16028 389836
rect 16080 389824 16086 389836
rect 528738 389824 528744 389836
rect 16080 389796 528744 389824
rect 16080 389784 16086 389796
rect 528738 389784 528744 389796
rect 528796 389784 528802 389836
rect 25958 389444 25964 389496
rect 26016 389484 26022 389496
rect 146938 389484 146944 389496
rect 26016 389456 146944 389484
rect 26016 389444 26022 389456
rect 146938 389444 146944 389456
rect 146996 389444 147002 389496
rect 36814 389376 36820 389428
rect 36872 389416 36878 389428
rect 52454 389416 52460 389428
rect 36872 389388 52460 389416
rect 36872 389376 36878 389388
rect 52454 389376 52460 389388
rect 52512 389376 52518 389428
rect 232314 389376 232320 389428
rect 232372 389416 232378 389428
rect 251818 389416 251824 389428
rect 232372 389388 251824 389416
rect 232372 389376 232378 389388
rect 251818 389376 251824 389388
rect 251876 389376 251882 389428
rect 475378 389376 475384 389428
rect 475436 389416 475442 389428
rect 494698 389416 494704 389428
rect 475436 389388 494704 389416
rect 475436 389376 475442 389388
rect 494698 389376 494704 389388
rect 494756 389376 494762 389428
rect 43346 389308 43352 389360
rect 43404 389348 43410 389360
rect 62758 389348 62764 389360
rect 43404 389320 62764 389348
rect 43404 389308 43410 389320
rect 62758 389308 62764 389320
rect 62816 389308 62822 389360
rect 90450 389308 90456 389360
rect 90508 389348 90514 389360
rect 106366 389348 106372 389360
rect 90508 389320 106372 389348
rect 90508 389308 90514 389320
rect 106366 389308 106372 389320
rect 106424 389308 106430 389360
rect 116486 389308 116492 389360
rect 116544 389348 116550 389360
rect 133414 389348 133420 389360
rect 116544 389320 133420 389348
rect 116544 389308 116550 389320
rect 133414 389308 133420 389320
rect 133472 389308 133478 389360
rect 170490 389308 170496 389360
rect 170548 389348 170554 389360
rect 187786 389348 187792 389360
rect 170548 389320 187792 389348
rect 170548 389308 170554 389320
rect 187786 389308 187792 389320
rect 187844 389308 187850 389360
rect 197538 389308 197544 389360
rect 197596 389348 197602 389360
rect 214374 389348 214380 389360
rect 197596 389320 214380 389348
rect 197596 389308 197602 389320
rect 214374 389308 214380 389320
rect 214432 389308 214438 389360
rect 224494 389308 224500 389360
rect 224552 389348 224558 389360
rect 241514 389348 241520 389360
rect 224552 389320 241520 389348
rect 224552 389308 224558 389320
rect 241514 389308 241520 389320
rect 241572 389308 241578 389360
rect 413462 389308 413468 389360
rect 413520 389348 413526 389360
rect 430574 389348 430580 389360
rect 413520 389320 430580 389348
rect 413520 389308 413526 389320
rect 430574 389308 430580 389320
rect 430632 389308 430638 389360
rect 440510 389308 440516 389360
rect 440568 389348 440574 389360
rect 457254 389348 457260 389360
rect 440568 389320 457260 389348
rect 440568 389308 440574 389320
rect 457254 389308 457260 389320
rect 457312 389308 457318 389360
rect 468570 389308 468576 389360
rect 468628 389348 468634 389360
rect 484394 389348 484400 389360
rect 468628 389320 484400 389348
rect 468628 389308 468634 389320
rect 484394 389308 484400 389320
rect 484452 389308 484458 389360
rect 36722 389240 36728 389292
rect 36780 389280 36786 389292
rect 62114 389280 62120 389292
rect 36780 389252 62120 389280
rect 36780 389240 36786 389252
rect 62114 389240 62120 389252
rect 62172 389240 62178 389292
rect 64138 389240 64144 389292
rect 64196 389280 64202 389292
rect 89070 389280 89076 389292
rect 64196 389252 89076 389280
rect 64196 389240 64202 389252
rect 89070 389240 89076 389252
rect 89128 389240 89134 389292
rect 90358 389240 90364 389292
rect 90416 389280 90422 389292
rect 115934 389280 115940 389292
rect 90416 389252 115940 389280
rect 90416 389240 90422 389252
rect 115934 389240 115940 389252
rect 115992 389240 115998 389292
rect 116578 389240 116584 389292
rect 116636 389280 116642 389292
rect 142982 389280 142988 389292
rect 116636 389252 142988 389280
rect 116636 389240 116642 389252
rect 142982 389240 142988 389252
rect 143040 389240 143046 389292
rect 144270 389240 144276 389292
rect 144328 389280 144334 389292
rect 170030 389280 170036 389292
rect 144328 389252 170036 389280
rect 144328 389240 144334 389252
rect 170030 389240 170036 389252
rect 170088 389240 170094 389292
rect 178402 389240 178408 389292
rect 178460 389280 178466 389292
rect 200758 389280 200764 389292
rect 178460 389252 200764 389280
rect 178460 389240 178466 389252
rect 200758 389240 200764 389252
rect 200816 389240 200822 389292
rect 251450 389240 251456 389292
rect 251508 389280 251514 389292
rect 268286 389280 268292 389292
rect 251508 389252 268292 389280
rect 251508 389240 251514 389252
rect 268286 389240 268292 389252
rect 268344 389240 268350 389292
rect 279418 389240 279424 389292
rect 279476 389280 279482 389292
rect 295794 389280 295800 389292
rect 279476 389252 295800 389280
rect 279476 389240 279482 389252
rect 295794 389240 295800 389252
rect 295852 389240 295858 389292
rect 305638 389240 305644 389292
rect 305696 389280 305702 389292
rect 322382 389280 322388 389292
rect 305696 389252 322388 389280
rect 305696 389240 305702 389252
rect 322382 389240 322388 389252
rect 322440 389240 322446 389292
rect 335998 389240 336004 389292
rect 336056 389280 336062 389292
rect 349798 389280 349804 389292
rect 336056 389252 349804 389280
rect 336056 389240 336062 389252
rect 349798 389240 349804 389252
rect 349856 389240 349862 389292
rect 359550 389240 359556 389292
rect 359608 389280 359614 389292
rect 376294 389280 376300 389292
rect 359608 389252 376300 389280
rect 359608 389240 359614 389252
rect 376294 389240 376300 389252
rect 376352 389240 376358 389292
rect 386506 389240 386512 389292
rect 386564 389280 386570 389292
rect 403342 389280 403348 389292
rect 386564 389252 403348 389280
rect 386564 389240 386570 389252
rect 403342 389240 403348 389252
rect 403400 389240 403406 389292
rect 421282 389240 421288 389292
rect 421340 389280 421346 389292
rect 446398 389280 446404 389292
rect 421340 389252 446404 389280
rect 421340 389240 421346 389252
rect 446398 389240 446404 389252
rect 446456 389240 446462 389292
rect 494514 389240 494520 389292
rect 494572 389280 494578 389292
rect 511350 389280 511356 389292
rect 494572 389252 511356 389280
rect 494572 389240 494578 389252
rect 511350 389240 511356 389252
rect 511408 389240 511414 389292
rect 522298 389240 522304 389292
rect 522356 389280 522362 389292
rect 538398 389280 538404 389292
rect 522356 389252 538404 389280
rect 522356 389240 522362 389252
rect 538398 389240 538404 389252
rect 538456 389240 538462 389292
rect 62482 389172 62488 389224
rect 62540 389212 62546 389224
rect 79318 389212 79324 389224
rect 62540 389184 79324 389212
rect 62540 389172 62546 389184
rect 79318 389172 79324 389184
rect 79376 389172 79382 389224
rect 144178 389172 144184 389224
rect 144236 389212 144242 389224
rect 160278 389212 160284 389224
rect 144236 389184 160284 389212
rect 144236 389172 144242 389184
rect 160278 389172 160284 389184
rect 160336 389172 160342 389224
rect 171778 389172 171784 389224
rect 171836 389212 171842 389224
rect 197446 389212 197452 389224
rect 171836 389184 197452 389212
rect 171836 389172 171842 389184
rect 197446 389172 197452 389184
rect 197504 389172 197510 389224
rect 199378 389172 199384 389224
rect 199436 389212 199442 389224
rect 223942 389212 223948 389224
rect 199436 389184 223948 389212
rect 199436 389172 199442 389184
rect 223942 389172 223948 389184
rect 224000 389172 224006 389224
rect 225598 389172 225604 389224
rect 225656 389212 225662 389224
rect 251174 389212 251180 389224
rect 225656 389184 251180 389212
rect 225656 389172 225662 389184
rect 251174 389172 251180 389184
rect 251232 389172 251238 389224
rect 253198 389172 253204 389224
rect 253256 389212 253262 389224
rect 278038 389212 278044 389224
rect 253256 389184 278044 389212
rect 253256 389172 253262 389184
rect 278038 389172 278044 389184
rect 278096 389172 278102 389224
rect 279510 389172 279516 389224
rect 279568 389212 279574 389224
rect 305546 389212 305552 389224
rect 279568 389184 305552 389212
rect 279568 389172 279574 389184
rect 305546 389172 305552 389184
rect 305604 389172 305610 389224
rect 307018 389172 307024 389224
rect 307076 389212 307082 389224
rect 331950 389212 331956 389224
rect 307076 389184 331956 389212
rect 307076 389172 307082 389184
rect 331950 389172 331956 389184
rect 332008 389172 332014 389224
rect 333238 389172 333244 389224
rect 333296 389212 333302 389224
rect 359458 389212 359464 389224
rect 333296 389184 359464 389212
rect 333296 389172 333302 389184
rect 359458 389172 359464 389184
rect 359516 389172 359522 389224
rect 359734 389172 359740 389224
rect 359792 389212 359798 389224
rect 386046 389212 386052 389224
rect 359792 389184 386052 389212
rect 359792 389172 359798 389184
rect 386046 389172 386052 389184
rect 386104 389172 386110 389224
rect 387058 389172 387064 389224
rect 387116 389212 387122 389224
rect 412910 389212 412916 389224
rect 387116 389184 412916 389212
rect 387116 389172 387122 389184
rect 412910 389172 412916 389184
rect 412968 389172 412974 389224
rect 414658 389172 414664 389224
rect 414716 389212 414722 389224
rect 440234 389212 440240 389224
rect 414716 389184 440240 389212
rect 414716 389172 414722 389184
rect 440234 389172 440240 389184
rect 440292 389172 440298 389224
rect 442258 389172 442264 389224
rect 442316 389212 442322 389224
rect 467006 389212 467012 389224
rect 442316 389184 467012 389212
rect 442316 389172 442322 389184
rect 467006 389172 467012 389184
rect 467064 389172 467070 389224
rect 468478 389172 468484 389224
rect 468536 389212 468542 389224
rect 494054 389212 494060 389224
rect 468536 389184 494060 389212
rect 468536 389172 468542 389184
rect 494054 389172 494060 389184
rect 494112 389172 494118 389224
rect 496078 389172 496084 389224
rect 496136 389212 496142 389224
rect 520918 389212 520924 389224
rect 496136 389184 520924 389212
rect 496136 389172 496142 389184
rect 520918 389172 520924 389184
rect 520976 389172 520982 389224
rect 522390 389172 522396 389224
rect 522448 389212 522454 389224
rect 548058 389212 548064 389224
rect 522448 389184 548064 389212
rect 522448 389172 522454 389184
rect 548058 389172 548064 389184
rect 548116 389172 548122 389224
rect 37918 387064 37924 387116
rect 37976 387104 37982 387116
rect 526438 387104 526444 387116
rect 37976 387076 526444 387104
rect 37976 387064 37982 387076
rect 526438 387064 526444 387076
rect 526496 387064 526502 387116
rect 285766 386248 285772 386300
rect 285824 386288 285830 386300
rect 286134 386288 286140 386300
rect 285824 386260 286140 386288
rect 285824 386248 285830 386260
rect 286134 386248 286140 386260
rect 286192 386248 286198 386300
rect 339586 386248 339592 386300
rect 339644 386288 339650 386300
rect 340138 386288 340144 386300
rect 339644 386260 340144 386288
rect 339644 386248 339650 386260
rect 340138 386248 340144 386260
rect 340196 386248 340202 386300
rect 89714 370540 89720 370592
rect 89772 370580 89778 370592
rect 90450 370580 90456 370592
rect 89772 370552 90456 370580
rect 89772 370540 89778 370552
rect 90450 370540 90456 370552
rect 90508 370540 90514 370592
rect 13722 368432 13728 368484
rect 13780 368472 13786 368484
rect 64874 368472 64880 368484
rect 13780 368444 64880 368472
rect 13780 368432 13786 368444
rect 64874 368432 64880 368444
rect 64932 368432 64938 368484
rect 95142 368432 95148 368484
rect 95200 368472 95206 368484
rect 144822 368472 144828 368484
rect 95200 368444 144828 368472
rect 95200 368432 95206 368444
rect 144822 368432 144828 368444
rect 144880 368432 144886 368484
rect 148962 368432 148968 368484
rect 149020 368472 149026 368484
rect 200114 368472 200120 368484
rect 149020 368444 200120 368472
rect 149020 368432 149026 368444
rect 200114 368432 200120 368444
rect 200172 368432 200178 368484
rect 202782 368432 202788 368484
rect 202840 368472 202846 368484
rect 253934 368472 253940 368484
rect 202840 368444 253940 368472
rect 202840 368432 202846 368444
rect 253934 368432 253940 368444
rect 253992 368432 253998 368484
rect 284202 368432 284208 368484
rect 284260 368472 284266 368484
rect 335354 368472 335360 368484
rect 284260 368444 335360 368472
rect 284260 368432 284266 368444
rect 335354 368432 335360 368444
rect 335412 368432 335418 368484
rect 338022 368432 338028 368484
rect 338080 368472 338086 368484
rect 389174 368472 389180 368484
rect 338080 368444 389180 368472
rect 338080 368432 338086 368444
rect 389174 368432 389180 368444
rect 389232 368432 389238 368484
rect 391842 368432 391848 368484
rect 391900 368472 391906 368484
rect 442994 368472 443000 368484
rect 391900 368444 443000 368472
rect 391900 368432 391906 368444
rect 442994 368432 443000 368444
rect 443052 368432 443058 368484
rect 446398 368432 446404 368484
rect 446456 368472 446462 368484
rect 447686 368472 447692 368484
rect 446456 368444 447692 368472
rect 446456 368432 446462 368444
rect 447686 368432 447692 368444
rect 447744 368432 447750 368484
rect 496814 368472 496820 368484
rect 448532 368444 496820 368472
rect 41322 368364 41328 368416
rect 41380 368404 41386 368416
rect 91094 368404 91100 368416
rect 41380 368376 91100 368404
rect 41380 368364 41386 368376
rect 91094 368364 91100 368376
rect 91152 368364 91158 368416
rect 122742 368364 122748 368416
rect 122800 368404 122806 368416
rect 172514 368404 172520 368416
rect 122800 368376 172520 368404
rect 122800 368364 122806 368376
rect 172514 368364 172520 368376
rect 172572 368364 172578 368416
rect 176562 368364 176568 368416
rect 176620 368404 176626 368416
rect 226334 368404 226340 368416
rect 176620 368376 226340 368404
rect 176620 368364 176626 368376
rect 226334 368364 226340 368376
rect 226392 368364 226398 368416
rect 256602 368364 256608 368416
rect 256660 368404 256666 368416
rect 307754 368404 307760 368416
rect 256660 368376 307760 368404
rect 256660 368364 256666 368376
rect 307754 368364 307760 368376
rect 307812 368364 307818 368416
rect 311802 368364 311808 368416
rect 311860 368404 311866 368416
rect 361574 368404 361580 368416
rect 311860 368376 361580 368404
rect 311860 368364 311866 368376
rect 361574 368364 361580 368376
rect 361632 368364 361638 368416
rect 365622 368364 365628 368416
rect 365680 368404 365686 368416
rect 415394 368404 415400 368416
rect 365680 368376 415400 368404
rect 365680 368364 365686 368376
rect 415394 368364 415400 368376
rect 415452 368364 415458 368416
rect 419442 368364 419448 368416
rect 419500 368404 419506 368416
rect 419500 368376 431954 368404
rect 419500 368364 419506 368376
rect 68922 368296 68928 368348
rect 68980 368336 68986 368348
rect 118694 368336 118700 368348
rect 68980 368308 118700 368336
rect 68980 368296 68986 368308
rect 118694 368296 118700 368308
rect 118752 368296 118758 368348
rect 230382 368296 230388 368348
rect 230440 368336 230446 368348
rect 280154 368336 280160 368348
rect 230440 368308 280160 368336
rect 230440 368296 230446 368308
rect 280154 368296 280160 368308
rect 280212 368296 280218 368348
rect 431926 368268 431954 368376
rect 445662 368296 445668 368348
rect 445720 368336 445726 368348
rect 448532 368336 448560 368444
rect 496814 368432 496820 368444
rect 496872 368432 496878 368484
rect 500862 368432 500868 368484
rect 500920 368472 500926 368484
rect 550634 368472 550640 368484
rect 500920 368444 550640 368472
rect 500920 368432 500926 368444
rect 550634 368432 550640 368444
rect 550692 368432 550698 368484
rect 469214 368404 469220 368416
rect 445720 368308 448560 368336
rect 451246 368376 469220 368404
rect 445720 368296 445726 368308
rect 451246 368268 451274 368376
rect 469214 368364 469220 368376
rect 469272 368364 469278 368416
rect 473262 368364 473268 368416
rect 473320 368404 473326 368416
rect 523034 368404 523040 368416
rect 473320 368376 523040 368404
rect 473320 368364 473326 368376
rect 523034 368364 523040 368376
rect 523092 368364 523098 368416
rect 467650 368296 467656 368348
rect 467708 368336 467714 368348
rect 468570 368336 468576 368348
rect 467708 368308 468576 368336
rect 467708 368296 467714 368308
rect 468570 368296 468576 368308
rect 468628 368296 468634 368348
rect 431926 368240 451274 368268
rect 170214 367616 170220 367668
rect 170272 367656 170278 367668
rect 170490 367656 170496 367668
rect 170272 367628 170496 367656
rect 170272 367616 170278 367628
rect 170490 367616 170496 367628
rect 170548 367616 170554 367668
rect 35618 367004 35624 367056
rect 35676 367044 35682 367056
rect 36814 367044 36820 367056
rect 35676 367016 36820 367044
rect 35676 367004 35682 367016
rect 36814 367004 36820 367016
rect 36872 367004 36878 367056
rect 53098 365644 53104 365696
rect 53156 365684 53162 365696
rect 64138 365684 64144 365696
rect 53156 365656 64144 365684
rect 53156 365644 53162 365656
rect 64138 365644 64144 365656
rect 64196 365644 64202 365696
rect 69106 365644 69112 365696
rect 69164 365684 69170 365696
rect 69164 365656 74534 365684
rect 69164 365644 69170 365656
rect 15194 365576 15200 365628
rect 15252 365616 15258 365628
rect 42794 365616 42800 365628
rect 15252 365588 42800 365616
rect 15252 365576 15258 365588
rect 42794 365576 42800 365588
rect 42852 365576 42858 365628
rect 62758 365576 62764 365628
rect 62816 365616 62822 365628
rect 69750 365616 69756 365628
rect 62816 365588 69756 365616
rect 62816 365576 62822 365588
rect 69750 365576 69756 365588
rect 69808 365576 69814 365628
rect 74506 365616 74534 365656
rect 96706 365644 96712 365696
rect 96764 365684 96770 365696
rect 96764 365656 103514 365684
rect 96764 365644 96770 365656
rect 96798 365616 96804 365628
rect 74506 365588 96804 365616
rect 96798 365576 96804 365588
rect 96856 365576 96862 365628
rect 103486 365616 103514 365656
rect 200758 365644 200764 365696
rect 200816 365684 200822 365696
rect 204622 365684 204628 365696
rect 200816 365656 204628 365684
rect 200816 365644 200822 365656
rect 204622 365644 204628 365656
rect 204680 365644 204686 365696
rect 251818 365644 251824 365696
rect 251876 365684 251882 365696
rect 258718 365684 258724 365696
rect 251876 365656 258724 365684
rect 251876 365644 251882 365656
rect 258718 365644 258724 365656
rect 258776 365644 258782 365696
rect 332502 365644 332508 365696
rect 332560 365684 332566 365696
rect 335998 365684 336004 365696
rect 332560 365656 336004 365684
rect 332560 365644 332566 365656
rect 335998 365644 336004 365656
rect 336056 365644 336062 365696
rect 494698 365644 494704 365696
rect 494756 365684 494762 365696
rect 501598 365684 501604 365696
rect 494756 365656 501604 365684
rect 494756 365644 494762 365656
rect 501598 365644 501604 365656
rect 501656 365644 501662 365696
rect 123662 365616 123668 365628
rect 103486 365588 123668 365616
rect 123662 365576 123668 365588
rect 123720 365576 123726 365628
rect 149698 365576 149704 365628
rect 149756 365616 149762 365628
rect 548058 365616 548064 365628
rect 149756 365588 548064 365616
rect 149756 365576 149762 365588
rect 548058 365576 548064 365588
rect 548116 365576 548122 365628
rect 26050 365508 26056 365560
rect 26108 365548 26114 365560
rect 36722 365548 36728 365560
rect 26108 365520 36728 365548
rect 26108 365508 26114 365520
rect 36722 365508 36728 365520
rect 36780 365508 36786 365560
rect 79962 365508 79968 365560
rect 80020 365548 80026 365560
rect 90358 365548 90364 365560
rect 80020 365520 90364 365548
rect 80020 365508 80026 365520
rect 90358 365508 90364 365520
rect 90416 365508 90422 365560
rect 106550 365508 106556 365560
rect 106608 365548 106614 365560
rect 116578 365548 116584 365560
rect 106608 365520 116584 365548
rect 106608 365508 106614 365520
rect 116578 365508 116584 365520
rect 116636 365508 116642 365560
rect 133782 365508 133788 365560
rect 133840 365548 133846 365560
rect 144270 365548 144276 365560
rect 133840 365520 144276 365548
rect 133840 365508 133846 365520
rect 144270 365508 144276 365520
rect 144328 365508 144334 365560
rect 150526 365508 150532 365560
rect 150584 365548 150590 365560
rect 178126 365548 178132 365560
rect 150584 365520 178132 365548
rect 150584 365508 150590 365520
rect 178126 365508 178132 365520
rect 178184 365508 178190 365560
rect 187970 365508 187976 365560
rect 188028 365548 188034 365560
rect 199378 365548 199384 365560
rect 188028 365520 199384 365548
rect 188028 365508 188034 365520
rect 199378 365508 199384 365520
rect 199436 365508 199442 365560
rect 204346 365508 204352 365560
rect 204404 365548 204410 365560
rect 231854 365548 231860 365560
rect 204404 365520 231860 365548
rect 204404 365508 204410 365520
rect 231854 365508 231860 365520
rect 231912 365508 231918 365560
rect 242066 365508 242072 365560
rect 242124 365548 242130 365560
rect 253198 365548 253204 365560
rect 242124 365520 253204 365548
rect 242124 365508 242130 365520
rect 253198 365508 253204 365520
rect 253256 365508 253262 365560
rect 258166 365508 258172 365560
rect 258224 365548 258230 365560
rect 286134 365548 286140 365560
rect 258224 365520 286140 365548
rect 258224 365508 258230 365520
rect 286134 365508 286140 365520
rect 286192 365508 286198 365560
rect 312630 365548 312636 365560
rect 287026 365520 312636 365548
rect 122926 365440 122932 365492
rect 122984 365480 122990 365492
rect 150710 365480 150716 365492
rect 122984 365452 150716 365480
rect 122984 365440 122990 365452
rect 150710 365440 150716 365452
rect 150768 365440 150774 365492
rect 160554 365440 160560 365492
rect 160612 365480 160618 365492
rect 171778 365480 171784 365492
rect 160612 365452 171784 365480
rect 160612 365440 160618 365452
rect 171778 365440 171784 365452
rect 171836 365440 171842 365492
rect 215018 365440 215024 365492
rect 215076 365480 215082 365492
rect 225598 365480 225604 365492
rect 215076 365452 225604 365480
rect 215076 365440 215082 365452
rect 225598 365440 225604 365452
rect 225656 365440 225662 365492
rect 268930 365440 268936 365492
rect 268988 365480 268994 365492
rect 279510 365480 279516 365492
rect 268988 365452 279516 365480
rect 268988 365440 268994 365452
rect 279510 365440 279516 365452
rect 279568 365440 279574 365492
rect 285766 365440 285772 365492
rect 285824 365480 285830 365492
rect 287026 365480 287054 365520
rect 312630 365508 312636 365520
rect 312688 365508 312694 365560
rect 340138 365548 340144 365560
rect 316006 365520 340144 365548
rect 285824 365452 287054 365480
rect 285824 365440 285830 365452
rect 295978 365440 295984 365492
rect 296036 365480 296042 365492
rect 307018 365480 307024 365492
rect 296036 365452 307024 365480
rect 296036 365440 296042 365452
rect 307018 365440 307024 365452
rect 307076 365440 307082 365492
rect 311986 365440 311992 365492
rect 312044 365480 312050 365492
rect 316006 365480 316034 365520
rect 340138 365508 340144 365520
rect 340196 365508 340202 365560
rect 366726 365548 366732 365560
rect 344986 365520 366732 365548
rect 312044 365452 316034 365480
rect 312044 365440 312050 365452
rect 322842 365440 322848 365492
rect 322900 365480 322906 365492
rect 333238 365480 333244 365492
rect 322900 365452 333244 365480
rect 322900 365440 322906 365452
rect 333238 365440 333244 365452
rect 333296 365440 333302 365492
rect 339586 365440 339592 365492
rect 339644 365480 339650 365492
rect 344986 365480 345014 365520
rect 366726 365508 366732 365520
rect 366784 365508 366790 365560
rect 393590 365548 393596 365560
rect 373966 365520 393596 365548
rect 339644 365452 345014 365480
rect 339644 365440 339650 365452
rect 350074 365440 350080 365492
rect 350132 365480 350138 365492
rect 359550 365480 359556 365492
rect 350132 365452 359556 365480
rect 350132 365440 350138 365452
rect 359550 365440 359556 365452
rect 359608 365440 359614 365492
rect 365806 365440 365812 365492
rect 365864 365480 365870 365492
rect 373966 365480 373994 365520
rect 393590 365508 393596 365520
rect 393648 365508 393654 365560
rect 420914 365548 420920 365560
rect 402946 365520 420920 365548
rect 365864 365452 373994 365480
rect 365864 365440 365870 365452
rect 376570 365440 376576 365492
rect 376628 365480 376634 365492
rect 387058 365480 387064 365492
rect 376628 365452 387064 365480
rect 376628 365440 376634 365452
rect 387058 365440 387064 365452
rect 387116 365440 387122 365492
rect 393406 365440 393412 365492
rect 393464 365480 393470 365492
rect 402946 365480 402974 365520
rect 420914 365508 420920 365520
rect 420972 365508 420978 365560
rect 431034 365508 431040 365560
rect 431092 365548 431098 365560
rect 442258 365548 442264 365560
rect 431092 365520 442264 365548
rect 431092 365508 431098 365520
rect 442258 365508 442264 365520
rect 442316 365508 442322 365560
rect 447226 365508 447232 365560
rect 447284 365548 447290 365560
rect 474734 365548 474740 365560
rect 447284 365520 474740 365548
rect 447284 365508 447290 365520
rect 474734 365508 474740 365520
rect 474792 365508 474798 365560
rect 484946 365508 484952 365560
rect 485004 365548 485010 365560
rect 496078 365548 496084 365560
rect 485004 365520 496084 365548
rect 485004 365508 485010 365520
rect 496078 365508 496084 365520
rect 496136 365508 496142 365560
rect 501046 365508 501052 365560
rect 501104 365548 501110 365560
rect 528646 365548 528652 365560
rect 501104 365520 528652 365548
rect 501104 365508 501110 365520
rect 528646 365508 528652 365520
rect 528704 365508 528710 365560
rect 393464 365452 402974 365480
rect 393464 365440 393470 365452
rect 403986 365440 403992 365492
rect 404044 365480 404050 365492
rect 414658 365480 414664 365492
rect 404044 365452 414664 365480
rect 404044 365440 404050 365452
rect 414658 365440 414664 365452
rect 414716 365440 414722 365492
rect 458082 365440 458088 365492
rect 458140 365480 458146 365492
rect 468478 365480 468484 365492
rect 458140 365452 468484 365480
rect 458140 365440 458146 365452
rect 468478 365440 468484 365452
rect 468536 365440 468542 365492
rect 511902 365440 511908 365492
rect 511960 365480 511966 365492
rect 522390 365480 522396 365492
rect 511960 365452 522396 365480
rect 511960 365440 511966 365452
rect 522390 365440 522396 365452
rect 522448 365440 522454 365492
rect 36630 365372 36636 365424
rect 36688 365412 36694 365424
rect 538398 365412 538404 365424
rect 36688 365384 538404 365412
rect 36688 365372 36694 365384
rect 538398 365372 538404 365384
rect 538456 365372 538462 365424
rect 16114 362176 16120 362228
rect 16172 362216 16178 362228
rect 529014 362216 529020 362228
rect 16172 362188 529020 362216
rect 16172 362176 16178 362188
rect 529014 362176 529020 362188
rect 529072 362176 529078 362228
rect 25682 361836 25688 361888
rect 25740 361876 25746 361888
rect 149698 361876 149704 361888
rect 25740 361848 149704 361876
rect 25740 361836 25746 361848
rect 149698 361836 149704 361848
rect 149756 361836 149762 361888
rect 36814 361768 36820 361820
rect 36872 361808 36878 361820
rect 52638 361808 52644 361820
rect 36872 361780 52644 361808
rect 36872 361768 36878 361780
rect 52638 361768 52644 361780
rect 52696 361768 52702 361820
rect 232038 361768 232044 361820
rect 232096 361808 232102 361820
rect 251818 361808 251824 361820
rect 232096 361780 251824 361808
rect 232096 361768 232102 361780
rect 251818 361768 251824 361780
rect 251876 361768 251882 361820
rect 475010 361768 475016 361820
rect 475068 361808 475074 361820
rect 494698 361808 494704 361820
rect 475068 361780 494704 361808
rect 475068 361768 475074 361780
rect 494698 361768 494704 361780
rect 494756 361768 494762 361820
rect 62482 361700 62488 361752
rect 62540 361740 62546 361752
rect 79686 361740 79692 361752
rect 62540 361712 79692 361740
rect 62540 361700 62546 361712
rect 79686 361700 79692 361712
rect 79744 361700 79750 361752
rect 90358 361700 90364 361752
rect 90416 361740 90422 361752
rect 106642 361740 106648 361752
rect 90416 361712 106648 361740
rect 90416 361700 90422 361712
rect 106642 361700 106648 361712
rect 106700 361700 106706 361752
rect 116486 361700 116492 361752
rect 116544 361740 116550 361752
rect 133690 361740 133696 361752
rect 116544 361712 133696 361740
rect 116544 361700 116550 361712
rect 133690 361700 133696 361712
rect 133748 361700 133754 361752
rect 144270 361700 144276 361752
rect 144328 361740 144334 361752
rect 160646 361740 160652 361752
rect 144328 361712 160652 361740
rect 144328 361700 144334 361712
rect 160646 361700 160652 361712
rect 160704 361700 160710 361752
rect 170490 361700 170496 361752
rect 170548 361740 170554 361752
rect 187694 361740 187700 361752
rect 170548 361712 187700 361740
rect 170548 361700 170554 361712
rect 187694 361700 187700 361712
rect 187752 361700 187758 361752
rect 197446 361700 197452 361752
rect 197504 361740 197510 361752
rect 214650 361740 214656 361752
rect 197504 361712 214656 361740
rect 197504 361700 197510 361712
rect 214650 361700 214656 361712
rect 214708 361700 214714 361752
rect 224494 361700 224500 361752
rect 224552 361740 224558 361752
rect 241698 361740 241704 361752
rect 224552 361712 241704 361740
rect 224552 361700 224558 361712
rect 241698 361700 241704 361712
rect 241756 361700 241762 361752
rect 413462 361700 413468 361752
rect 413520 361740 413526 361752
rect 430666 361740 430672 361752
rect 413520 361712 430672 361740
rect 413520 361700 413526 361712
rect 430666 361700 430672 361712
rect 430724 361700 430730 361752
rect 440510 361700 440516 361752
rect 440568 361740 440574 361752
rect 457622 361740 457628 361752
rect 440568 361712 457628 361740
rect 440568 361700 440574 361712
rect 457622 361700 457628 361712
rect 457680 361700 457686 361752
rect 468570 361700 468576 361752
rect 468628 361740 468634 361752
rect 484670 361740 484676 361752
rect 468628 361712 484676 361740
rect 468628 361700 468634 361712
rect 484670 361700 484676 361712
rect 484728 361700 484734 361752
rect 36630 361632 36636 361684
rect 36688 361672 36694 361684
rect 62298 361672 62304 361684
rect 36688 361644 62304 361672
rect 36688 361632 36694 361644
rect 62298 361632 62304 361644
rect 62356 361632 62362 361684
rect 64138 361632 64144 361684
rect 64196 361672 64202 361684
rect 89346 361672 89352 361684
rect 64196 361644 89352 361672
rect 64196 361632 64202 361644
rect 89346 361632 89352 361644
rect 89404 361632 89410 361684
rect 90450 361632 90456 361684
rect 90508 361672 90514 361684
rect 116302 361672 116308 361684
rect 90508 361644 116308 361672
rect 90508 361632 90514 361644
rect 116302 361632 116308 361644
rect 116360 361632 116366 361684
rect 116578 361632 116584 361684
rect 116636 361672 116642 361684
rect 143350 361672 143356 361684
rect 116636 361644 143356 361672
rect 116636 361632 116642 361644
rect 143350 361632 143356 361644
rect 143408 361632 143414 361684
rect 144178 361632 144184 361684
rect 144236 361672 144242 361684
rect 170306 361672 170312 361684
rect 144236 361644 170312 361672
rect 144236 361632 144242 361644
rect 170306 361632 170312 361644
rect 170364 361632 170370 361684
rect 178034 361632 178040 361684
rect 178092 361672 178098 361684
rect 200758 361672 200764 361684
rect 178092 361644 200764 361672
rect 178092 361632 178098 361644
rect 200758 361632 200764 361644
rect 200816 361632 200822 361684
rect 251450 361632 251456 361684
rect 251508 361672 251514 361684
rect 268654 361672 268660 361684
rect 251508 361644 268660 361672
rect 251508 361632 251514 361644
rect 268654 361632 268660 361644
rect 268712 361632 268718 361684
rect 279510 361632 279516 361684
rect 279568 361672 279574 361684
rect 295702 361672 295708 361684
rect 279568 361644 295708 361672
rect 279568 361632 279574 361644
rect 295702 361632 295708 361644
rect 295760 361632 295766 361684
rect 305454 361632 305460 361684
rect 305512 361672 305518 361684
rect 322658 361672 322664 361684
rect 305512 361644 322664 361672
rect 305512 361632 305518 361644
rect 322658 361632 322664 361644
rect 322716 361632 322722 361684
rect 334618 361632 334624 361684
rect 334676 361672 334682 361684
rect 349706 361672 349712 361684
rect 334676 361644 349712 361672
rect 334676 361632 334682 361644
rect 349706 361632 349712 361644
rect 349764 361632 349770 361684
rect 359458 361632 359464 361684
rect 359516 361672 359522 361684
rect 376662 361672 376668 361684
rect 359516 361644 376668 361672
rect 359516 361632 359522 361644
rect 376662 361632 376668 361644
rect 376720 361632 376726 361684
rect 386506 361632 386512 361684
rect 386564 361672 386570 361684
rect 403618 361672 403624 361684
rect 386564 361644 403624 361672
rect 386564 361632 386570 361644
rect 403618 361632 403624 361644
rect 403676 361632 403682 361684
rect 421006 361632 421012 361684
rect 421064 361672 421070 361684
rect 443638 361672 443644 361684
rect 421064 361644 443644 361672
rect 421064 361632 421070 361644
rect 443638 361632 443644 361644
rect 443696 361632 443702 361684
rect 494514 361632 494520 361684
rect 494572 361672 494578 361684
rect 511626 361672 511632 361684
rect 494572 361644 511632 361672
rect 494572 361632 494578 361644
rect 511626 361632 511632 361644
rect 511684 361632 511690 361684
rect 522298 361632 522304 361684
rect 522356 361672 522362 361684
rect 538674 361672 538680 361684
rect 522356 361644 538680 361672
rect 522356 361632 522362 361644
rect 538674 361632 538680 361644
rect 538732 361632 538738 361684
rect 43070 361564 43076 361616
rect 43128 361604 43134 361616
rect 62758 361604 62764 361616
rect 43128 361576 62764 361604
rect 43128 361564 43134 361576
rect 62758 361564 62764 361576
rect 62816 361564 62822 361616
rect 171778 361564 171784 361616
rect 171836 361604 171842 361616
rect 197354 361604 197360 361616
rect 171836 361576 197360 361604
rect 171836 361564 171842 361576
rect 197354 361564 197360 361576
rect 197412 361564 197418 361616
rect 199378 361564 199384 361616
rect 199436 361604 199442 361616
rect 224310 361604 224316 361616
rect 199436 361576 224316 361604
rect 199436 361564 199442 361576
rect 224310 361564 224316 361576
rect 224368 361564 224374 361616
rect 225598 361564 225604 361616
rect 225656 361604 225662 361616
rect 251358 361604 251364 361616
rect 225656 361576 251364 361604
rect 225656 361564 225662 361576
rect 251358 361564 251364 361576
rect 251416 361564 251422 361616
rect 253198 361564 253204 361616
rect 253256 361604 253262 361616
rect 278314 361604 278320 361616
rect 253256 361576 278320 361604
rect 253256 361564 253262 361576
rect 278314 361564 278320 361576
rect 278372 361564 278378 361616
rect 279418 361564 279424 361616
rect 279476 361604 279482 361616
rect 305362 361604 305368 361616
rect 279476 361576 305368 361604
rect 279476 361564 279482 361576
rect 305362 361564 305368 361576
rect 305420 361564 305426 361616
rect 307018 361564 307024 361616
rect 307076 361604 307082 361616
rect 332318 361604 332324 361616
rect 307076 361576 332324 361604
rect 307076 361564 307082 361576
rect 332318 361564 332324 361576
rect 332376 361564 332382 361616
rect 333238 361564 333244 361616
rect 333296 361604 333302 361616
rect 359366 361604 359372 361616
rect 333296 361576 359372 361604
rect 333296 361564 333302 361576
rect 359366 361564 359372 361576
rect 359424 361564 359430 361616
rect 359550 361564 359556 361616
rect 359608 361604 359614 361616
rect 386322 361604 386328 361616
rect 359608 361576 386328 361604
rect 359608 361564 359614 361576
rect 386322 361564 386328 361576
rect 386380 361564 386386 361616
rect 387058 361564 387064 361616
rect 387116 361604 387122 361616
rect 413278 361604 413284 361616
rect 387116 361576 413284 361604
rect 387116 361564 387122 361576
rect 413278 361564 413284 361576
rect 413336 361564 413342 361616
rect 414658 361564 414664 361616
rect 414716 361604 414722 361616
rect 440326 361604 440332 361616
rect 414716 361576 440332 361604
rect 414716 361564 414722 361576
rect 440326 361564 440332 361576
rect 440384 361564 440390 361616
rect 442258 361564 442264 361616
rect 442316 361604 442322 361616
rect 467282 361604 467288 361616
rect 442316 361576 467288 361604
rect 442316 361564 442322 361576
rect 467282 361564 467288 361576
rect 467340 361564 467346 361616
rect 468478 361564 468484 361616
rect 468536 361604 468542 361616
rect 494330 361604 494336 361616
rect 468536 361576 494336 361604
rect 468536 361564 468542 361576
rect 494330 361564 494336 361576
rect 494388 361564 494394 361616
rect 496078 361564 496084 361616
rect 496136 361604 496142 361616
rect 521286 361604 521292 361616
rect 496136 361576 521292 361604
rect 496136 361564 496142 361576
rect 521286 361564 521292 361576
rect 521344 361564 521350 361616
rect 522390 361564 522396 361616
rect 522448 361604 522454 361616
rect 548334 361604 548340 361616
rect 522448 361576 548340 361604
rect 522448 361564 522454 361576
rect 548334 361564 548340 361576
rect 548392 361564 548398 361616
rect 37918 359456 37924 359508
rect 37976 359496 37982 359508
rect 526438 359496 526444 359508
rect 37976 359468 526444 359496
rect 37976 359456 37982 359468
rect 526438 359456 526444 359468
rect 526496 359456 526502 359508
rect 35618 358776 35624 358828
rect 35676 358816 35682 358828
rect 36722 358816 36728 358828
rect 35676 358788 36728 358816
rect 35676 358776 35682 358788
rect 36722 358776 36728 358788
rect 36780 358776 36786 358828
rect 143626 342524 143632 342576
rect 143684 342564 143690 342576
rect 144270 342564 144276 342576
rect 143684 342536 144276 342564
rect 143684 342524 143690 342536
rect 144270 342524 144276 342536
rect 144328 342524 144334 342576
rect 443638 340892 443644 340944
rect 443696 340932 443702 340944
rect 447686 340932 447692 340944
rect 443696 340904 447692 340932
rect 443696 340892 443702 340904
rect 447686 340892 447692 340904
rect 447744 340892 447750 340944
rect 13722 340824 13728 340876
rect 13780 340864 13786 340876
rect 64874 340864 64880 340876
rect 13780 340836 64880 340864
rect 13780 340824 13786 340836
rect 64874 340824 64880 340836
rect 64932 340824 64938 340876
rect 95142 340824 95148 340876
rect 95200 340864 95206 340876
rect 146294 340864 146300 340876
rect 95200 340836 146300 340864
rect 95200 340824 95206 340836
rect 146294 340824 146300 340836
rect 146352 340824 146358 340876
rect 148962 340824 148968 340876
rect 149020 340864 149026 340876
rect 200114 340864 200120 340876
rect 149020 340836 200120 340864
rect 149020 340824 149026 340836
rect 200114 340824 200120 340836
rect 200172 340824 200178 340876
rect 202782 340824 202788 340876
rect 202840 340864 202846 340876
rect 253934 340864 253940 340876
rect 202840 340836 253940 340864
rect 202840 340824 202846 340836
rect 253934 340824 253940 340836
rect 253992 340824 253998 340876
rect 256602 340824 256608 340876
rect 256660 340864 256666 340876
rect 307754 340864 307760 340876
rect 256660 340836 307760 340864
rect 256660 340824 256666 340836
rect 307754 340824 307760 340836
rect 307812 340824 307818 340876
rect 332502 340824 332508 340876
rect 332560 340864 332566 340876
rect 334618 340864 334624 340876
rect 332560 340836 334624 340864
rect 332560 340824 332566 340836
rect 334618 340824 334624 340836
rect 334676 340824 334682 340876
rect 338022 340824 338028 340876
rect 338080 340864 338086 340876
rect 389174 340864 389180 340876
rect 338080 340836 389180 340864
rect 338080 340824 338086 340836
rect 389174 340824 389180 340836
rect 389232 340824 389238 340876
rect 391842 340824 391848 340876
rect 391900 340864 391906 340876
rect 442994 340864 443000 340876
rect 391900 340836 443000 340864
rect 391900 340824 391906 340836
rect 442994 340824 443000 340836
rect 443052 340824 443058 340876
rect 445662 340824 445668 340876
rect 445720 340864 445726 340876
rect 496814 340864 496820 340876
rect 445720 340836 496820 340864
rect 445720 340824 445726 340836
rect 496814 340824 496820 340836
rect 496872 340824 496878 340876
rect 500862 340824 500868 340876
rect 500920 340864 500926 340876
rect 550634 340864 550640 340876
rect 500920 340836 550640 340864
rect 500920 340824 500926 340836
rect 550634 340824 550640 340836
rect 550692 340824 550698 340876
rect 35618 340756 35624 340808
rect 35676 340796 35682 340808
rect 36814 340796 36820 340808
rect 35676 340768 36820 340796
rect 35676 340756 35682 340768
rect 36814 340756 36820 340768
rect 36872 340756 36878 340808
rect 41322 340756 41328 340808
rect 41380 340796 41386 340808
rect 91094 340796 91100 340808
rect 41380 340768 91100 340796
rect 41380 340756 41386 340768
rect 91094 340756 91100 340768
rect 91152 340756 91158 340808
rect 122742 340756 122748 340808
rect 122800 340796 122806 340808
rect 172514 340796 172520 340808
rect 122800 340768 172520 340796
rect 122800 340756 122806 340768
rect 172514 340756 172520 340768
rect 172572 340756 172578 340808
rect 176562 340756 176568 340808
rect 176620 340796 176626 340808
rect 226334 340796 226340 340808
rect 176620 340768 226340 340796
rect 176620 340756 176626 340768
rect 226334 340756 226340 340768
rect 226392 340756 226398 340808
rect 230382 340756 230388 340808
rect 230440 340796 230446 340808
rect 280154 340796 280160 340808
rect 230440 340768 280160 340796
rect 230440 340756 230446 340768
rect 280154 340756 280160 340768
rect 280212 340756 280218 340808
rect 284202 340756 284208 340808
rect 284260 340796 284266 340808
rect 335354 340796 335360 340808
rect 284260 340768 335360 340796
rect 284260 340756 284266 340768
rect 335354 340756 335360 340768
rect 335412 340756 335418 340808
rect 365622 340756 365628 340808
rect 365680 340796 365686 340808
rect 415394 340796 415400 340808
rect 365680 340768 415400 340796
rect 365680 340756 365686 340768
rect 415394 340756 415400 340768
rect 415452 340756 415458 340808
rect 419442 340756 419448 340808
rect 419500 340796 419506 340808
rect 469214 340796 469220 340808
rect 419500 340768 469220 340796
rect 419500 340756 419506 340768
rect 469214 340756 469220 340768
rect 469272 340756 469278 340808
rect 473262 340756 473268 340808
rect 473320 340796 473326 340808
rect 523034 340796 523040 340808
rect 473320 340768 523040 340796
rect 473320 340756 473326 340768
rect 523034 340756 523040 340768
rect 523092 340756 523098 340808
rect 68922 340688 68928 340740
rect 68980 340728 68986 340740
rect 118694 340728 118700 340740
rect 68980 340700 118700 340728
rect 68980 340688 68986 340700
rect 118694 340688 118700 340700
rect 118752 340688 118758 340740
rect 200758 340688 200764 340740
rect 200816 340728 200822 340740
rect 204622 340728 204628 340740
rect 200816 340700 204628 340728
rect 200816 340688 200822 340700
rect 204622 340688 204628 340700
rect 204680 340688 204686 340740
rect 278682 340688 278688 340740
rect 278740 340728 278746 340740
rect 279510 340728 279516 340740
rect 278740 340700 279516 340728
rect 278740 340688 278746 340700
rect 279510 340688 279516 340700
rect 279568 340688 279574 340740
rect 311802 340688 311808 340740
rect 311860 340728 311866 340740
rect 361574 340728 361580 340740
rect 311860 340700 361580 340728
rect 311860 340688 311866 340700
rect 361574 340688 361580 340700
rect 361632 340688 361638 340740
rect 467650 340688 467656 340740
rect 467708 340728 467714 340740
rect 468570 340728 468576 340740
rect 467708 340700 468576 340728
rect 467708 340688 467714 340700
rect 468570 340688 468576 340700
rect 468628 340688 468634 340740
rect 25682 338036 25688 338088
rect 25740 338076 25746 338088
rect 36630 338076 36636 338088
rect 25740 338048 36636 338076
rect 25740 338036 25746 338048
rect 36630 338036 36636 338048
rect 36688 338036 36694 338088
rect 52730 338036 52736 338088
rect 52788 338076 52794 338088
rect 64138 338076 64144 338088
rect 52788 338048 64144 338076
rect 52788 338036 52794 338048
rect 64138 338036 64144 338048
rect 64196 338036 64202 338088
rect 69106 338036 69112 338088
rect 69164 338076 69170 338088
rect 69164 338048 74534 338076
rect 69164 338036 69170 338048
rect 15194 337968 15200 338020
rect 15252 338008 15258 338020
rect 42978 338008 42984 338020
rect 15252 337980 42984 338008
rect 15252 337968 15258 337980
rect 42978 337968 42984 337980
rect 43036 337968 43042 338020
rect 62758 337968 62764 338020
rect 62816 338008 62822 338020
rect 70026 338008 70032 338020
rect 62816 337980 70032 338008
rect 62816 337968 62822 337980
rect 70026 337968 70032 337980
rect 70084 337968 70090 338020
rect 74506 338008 74534 338048
rect 96706 338036 96712 338088
rect 96764 338076 96770 338088
rect 96764 338048 103514 338076
rect 96764 338036 96770 338048
rect 96982 338008 96988 338020
rect 74506 337980 96988 338008
rect 96982 337968 96988 337980
rect 97040 337968 97046 338020
rect 103486 338008 103514 338048
rect 146938 338036 146944 338088
rect 146996 338076 147002 338088
rect 146996 338048 151814 338076
rect 146996 338036 147002 338048
rect 124030 338008 124036 338020
rect 103486 337980 124036 338008
rect 124030 337968 124036 337980
rect 124088 337968 124094 338020
rect 133690 337968 133696 338020
rect 133748 338008 133754 338020
rect 144178 338008 144184 338020
rect 133748 337980 144184 338008
rect 133748 337968 133754 337980
rect 144178 337968 144184 337980
rect 144236 337968 144242 338020
rect 150526 337968 150532 338020
rect 150584 338008 150590 338020
rect 151786 338008 151814 338048
rect 251818 338036 251824 338088
rect 251876 338076 251882 338088
rect 258994 338076 259000 338088
rect 251876 338048 259000 338076
rect 251876 338036 251882 338048
rect 258994 338036 259000 338048
rect 259052 338036 259058 338088
rect 494698 338036 494704 338088
rect 494756 338076 494762 338088
rect 501966 338076 501972 338088
rect 494756 338048 501972 338076
rect 494756 338036 494762 338048
rect 501966 338036 501972 338048
rect 502024 338036 502030 338088
rect 548334 338008 548340 338020
rect 150584 337980 151124 338008
rect 151786 337980 548340 338008
rect 150584 337968 150590 337980
rect 79686 337900 79692 337952
rect 79744 337940 79750 337952
rect 90450 337940 90456 337952
rect 79744 337912 90456 337940
rect 79744 337900 79750 337912
rect 90450 337900 90456 337912
rect 90508 337900 90514 337952
rect 106642 337900 106648 337952
rect 106700 337940 106706 337952
rect 116578 337940 116584 337952
rect 106700 337912 116584 337940
rect 106700 337900 106706 337912
rect 116578 337900 116584 337912
rect 116636 337900 116642 337952
rect 122926 337900 122932 337952
rect 122984 337940 122990 337952
rect 150986 337940 150992 337952
rect 122984 337912 150992 337940
rect 122984 337900 122990 337912
rect 150986 337900 150992 337912
rect 151044 337900 151050 337952
rect 151096 337940 151124 337980
rect 548334 337968 548340 337980
rect 548392 337968 548398 338020
rect 178034 337940 178040 337952
rect 151096 337912 178040 337940
rect 178034 337900 178040 337912
rect 178092 337900 178098 337952
rect 187694 337900 187700 337952
rect 187752 337940 187758 337952
rect 199378 337940 199384 337952
rect 187752 337912 199384 337940
rect 187752 337900 187758 337912
rect 199378 337900 199384 337912
rect 199436 337900 199442 337952
rect 204346 337900 204352 337952
rect 204404 337940 204410 337952
rect 232038 337940 232044 337952
rect 204404 337912 232044 337940
rect 204404 337900 204410 337912
rect 232038 337900 232044 337912
rect 232096 337900 232102 337952
rect 241698 337900 241704 337952
rect 241756 337940 241762 337952
rect 253198 337940 253204 337952
rect 241756 337912 253204 337940
rect 241756 337900 241762 337912
rect 253198 337900 253204 337912
rect 253256 337900 253262 337952
rect 258166 337900 258172 337952
rect 258224 337940 258230 337952
rect 286042 337940 286048 337952
rect 258224 337912 286048 337940
rect 258224 337900 258230 337912
rect 286042 337900 286048 337912
rect 286100 337900 286106 337952
rect 312998 337940 313004 337952
rect 287026 337912 313004 337940
rect 160646 337832 160652 337884
rect 160704 337872 160710 337884
rect 171778 337872 171784 337884
rect 160704 337844 171784 337872
rect 160704 337832 160710 337844
rect 171778 337832 171784 337844
rect 171836 337832 171842 337884
rect 214650 337832 214656 337884
rect 214708 337872 214714 337884
rect 225598 337872 225604 337884
rect 214708 337844 225604 337872
rect 214708 337832 214714 337844
rect 225598 337832 225604 337844
rect 225656 337832 225662 337884
rect 268654 337832 268660 337884
rect 268712 337872 268718 337884
rect 279418 337872 279424 337884
rect 268712 337844 279424 337872
rect 268712 337832 268718 337844
rect 279418 337832 279424 337844
rect 279476 337832 279482 337884
rect 285766 337832 285772 337884
rect 285824 337872 285830 337884
rect 287026 337872 287054 337912
rect 312998 337900 313004 337912
rect 313056 337900 313062 337952
rect 340046 337940 340052 337952
rect 316006 337912 340052 337940
rect 285824 337844 287054 337872
rect 285824 337832 285830 337844
rect 295702 337832 295708 337884
rect 295760 337872 295766 337884
rect 307018 337872 307024 337884
rect 295760 337844 307024 337872
rect 295760 337832 295766 337844
rect 307018 337832 307024 337844
rect 307076 337832 307082 337884
rect 311986 337832 311992 337884
rect 312044 337872 312050 337884
rect 316006 337872 316034 337912
rect 340046 337900 340052 337912
rect 340104 337900 340110 337952
rect 367002 337940 367008 337952
rect 344986 337912 367008 337940
rect 312044 337844 316034 337872
rect 312044 337832 312050 337844
rect 322658 337832 322664 337884
rect 322716 337872 322722 337884
rect 333238 337872 333244 337884
rect 322716 337844 333244 337872
rect 322716 337832 322722 337844
rect 333238 337832 333244 337844
rect 333296 337832 333302 337884
rect 339586 337832 339592 337884
rect 339644 337872 339650 337884
rect 344986 337872 345014 337912
rect 367002 337900 367008 337912
rect 367060 337900 367066 337952
rect 393958 337940 393964 337952
rect 373966 337912 393964 337940
rect 339644 337844 345014 337872
rect 339644 337832 339650 337844
rect 349706 337832 349712 337884
rect 349764 337872 349770 337884
rect 359550 337872 359556 337884
rect 349764 337844 359556 337872
rect 349764 337832 349770 337844
rect 359550 337832 359556 337844
rect 359608 337832 359614 337884
rect 365806 337832 365812 337884
rect 365864 337872 365870 337884
rect 373966 337872 373994 337912
rect 393958 337900 393964 337912
rect 394016 337900 394022 337952
rect 421006 337940 421012 337952
rect 402946 337912 421012 337940
rect 365864 337844 373994 337872
rect 365864 337832 365870 337844
rect 376662 337832 376668 337884
rect 376720 337872 376726 337884
rect 387058 337872 387064 337884
rect 376720 337844 387064 337872
rect 376720 337832 376726 337844
rect 387058 337832 387064 337844
rect 387116 337832 387122 337884
rect 393406 337832 393412 337884
rect 393464 337872 393470 337884
rect 402946 337872 402974 337912
rect 421006 337900 421012 337912
rect 421064 337900 421070 337952
rect 430666 337900 430672 337952
rect 430724 337940 430730 337952
rect 442258 337940 442264 337952
rect 430724 337912 442264 337940
rect 430724 337900 430730 337912
rect 442258 337900 442264 337912
rect 442316 337900 442322 337952
rect 447226 337900 447232 337952
rect 447284 337940 447290 337952
rect 475010 337940 475016 337952
rect 447284 337912 475016 337940
rect 447284 337900 447290 337912
rect 475010 337900 475016 337912
rect 475068 337900 475074 337952
rect 484670 337900 484676 337952
rect 484728 337940 484734 337952
rect 496078 337940 496084 337952
rect 484728 337912 496084 337940
rect 484728 337900 484734 337912
rect 496078 337900 496084 337912
rect 496136 337900 496142 337952
rect 501046 337900 501052 337952
rect 501104 337940 501110 337952
rect 529014 337940 529020 337952
rect 501104 337912 529020 337940
rect 501104 337900 501110 337912
rect 529014 337900 529020 337912
rect 529072 337900 529078 337952
rect 393464 337844 402974 337872
rect 393464 337832 393470 337844
rect 403710 337832 403716 337884
rect 403768 337872 403774 337884
rect 414658 337872 414664 337884
rect 403768 337844 414664 337872
rect 403768 337832 403774 337844
rect 414658 337832 414664 337844
rect 414716 337832 414722 337884
rect 457714 337832 457720 337884
rect 457772 337872 457778 337884
rect 468478 337872 468484 337884
rect 457772 337844 468484 337872
rect 457772 337832 457778 337844
rect 468478 337832 468484 337844
rect 468536 337832 468542 337884
rect 511718 337832 511724 337884
rect 511776 337872 511782 337884
rect 522390 337872 522396 337884
rect 511776 337844 522396 337872
rect 511776 337832 511782 337844
rect 522390 337832 522396 337844
rect 522448 337832 522454 337884
rect 36538 337764 36544 337816
rect 36596 337804 36602 337816
rect 538674 337804 538680 337816
rect 36596 337776 538680 337804
rect 36596 337764 36602 337776
rect 538674 337764 538680 337776
rect 538732 337764 538738 337816
rect 16022 335996 16028 336048
rect 16080 336036 16086 336048
rect 528646 336036 528652 336048
rect 16080 336008 528652 336036
rect 16080 335996 16086 336008
rect 528646 335996 528652 336008
rect 528704 335996 528710 336048
rect 26050 335588 26056 335640
rect 26108 335628 26114 335640
rect 146938 335628 146944 335640
rect 26108 335600 146944 335628
rect 26108 335588 26114 335600
rect 146938 335588 146944 335600
rect 146996 335588 147002 335640
rect 36538 335520 36544 335572
rect 36596 335560 36602 335572
rect 52454 335560 52460 335572
rect 36596 335532 52460 335560
rect 36596 335520 36602 335532
rect 52454 335520 52460 335532
rect 52512 335520 52518 335572
rect 232314 335520 232320 335572
rect 232372 335560 232378 335572
rect 251818 335560 251824 335572
rect 232372 335532 251824 335560
rect 232372 335520 232378 335532
rect 251818 335520 251824 335532
rect 251876 335520 251882 335572
rect 475378 335520 475384 335572
rect 475436 335560 475442 335572
rect 494698 335560 494704 335572
rect 475436 335532 494704 335560
rect 475436 335520 475442 335532
rect 494698 335520 494704 335532
rect 494756 335520 494762 335572
rect 62482 335452 62488 335504
rect 62540 335492 62546 335504
rect 79318 335492 79324 335504
rect 62540 335464 79324 335492
rect 62540 335452 62546 335464
rect 79318 335452 79324 335464
rect 79376 335452 79382 335504
rect 90450 335452 90456 335504
rect 90508 335492 90514 335504
rect 106458 335492 106464 335504
rect 90508 335464 106464 335492
rect 90508 335452 90514 335464
rect 106458 335452 106464 335464
rect 106516 335452 106522 335504
rect 116486 335452 116492 335504
rect 116544 335492 116550 335504
rect 133414 335492 133420 335504
rect 116544 335464 133420 335492
rect 116544 335452 116550 335464
rect 133414 335452 133420 335464
rect 133472 335452 133478 335504
rect 170490 335452 170496 335504
rect 170548 335492 170554 335504
rect 187786 335492 187792 335504
rect 170548 335464 187792 335492
rect 170548 335452 170554 335464
rect 187786 335452 187792 335464
rect 187844 335452 187850 335504
rect 197538 335452 197544 335504
rect 197596 335492 197602 335504
rect 214374 335492 214380 335504
rect 197596 335464 214380 335492
rect 197596 335452 197602 335464
rect 214374 335452 214380 335464
rect 214432 335452 214438 335504
rect 224494 335452 224500 335504
rect 224552 335492 224558 335504
rect 241606 335492 241612 335504
rect 224552 335464 241612 335492
rect 224552 335452 224558 335464
rect 241606 335452 241612 335464
rect 241664 335452 241670 335504
rect 413462 335452 413468 335504
rect 413520 335492 413526 335504
rect 430574 335492 430580 335504
rect 413520 335464 430580 335492
rect 413520 335452 413526 335464
rect 430574 335452 430580 335464
rect 430632 335452 430638 335504
rect 440510 335452 440516 335504
rect 440568 335492 440574 335504
rect 457254 335492 457260 335504
rect 440568 335464 457260 335492
rect 440568 335452 440574 335464
rect 457254 335452 457260 335464
rect 457312 335452 457318 335504
rect 468478 335452 468484 335504
rect 468536 335492 468542 335504
rect 484394 335492 484400 335504
rect 468536 335464 484400 335492
rect 468536 335452 468542 335464
rect 484394 335452 484400 335464
rect 484452 335452 484458 335504
rect 36814 335384 36820 335436
rect 36872 335424 36878 335436
rect 62114 335424 62120 335436
rect 36872 335396 62120 335424
rect 36872 335384 36878 335396
rect 62114 335384 62120 335396
rect 62172 335384 62178 335436
rect 64138 335384 64144 335436
rect 64196 335424 64202 335436
rect 89070 335424 89076 335436
rect 64196 335396 89076 335424
rect 64196 335384 64202 335396
rect 89070 335384 89076 335396
rect 89128 335384 89134 335436
rect 90358 335384 90364 335436
rect 90416 335424 90422 335436
rect 116118 335424 116124 335436
rect 90416 335396 116124 335424
rect 90416 335384 90422 335396
rect 116118 335384 116124 335396
rect 116176 335384 116182 335436
rect 116578 335384 116584 335436
rect 116636 335424 116642 335436
rect 142982 335424 142988 335436
rect 116636 335396 142988 335424
rect 116636 335384 116642 335396
rect 142982 335384 142988 335396
rect 143040 335384 143046 335436
rect 144270 335384 144276 335436
rect 144328 335424 144334 335436
rect 170030 335424 170036 335436
rect 144328 335396 170036 335424
rect 144328 335384 144334 335396
rect 170030 335384 170036 335396
rect 170088 335384 170094 335436
rect 178402 335384 178408 335436
rect 178460 335424 178466 335436
rect 200758 335424 200764 335436
rect 178460 335396 200764 335424
rect 178460 335384 178466 335396
rect 200758 335384 200764 335396
rect 200816 335384 200822 335436
rect 251450 335384 251456 335436
rect 251508 335424 251514 335436
rect 268286 335424 268292 335436
rect 251508 335396 268292 335424
rect 251508 335384 251514 335396
rect 268286 335384 268292 335396
rect 268344 335384 268350 335436
rect 279510 335384 279516 335436
rect 279568 335424 279574 335436
rect 295794 335424 295800 335436
rect 279568 335396 295800 335424
rect 279568 335384 279574 335396
rect 295794 335384 295800 335396
rect 295852 335384 295858 335436
rect 305546 335384 305552 335436
rect 305604 335424 305610 335436
rect 322382 335424 322388 335436
rect 305604 335396 322388 335424
rect 305604 335384 305610 335396
rect 322382 335384 322388 335396
rect 322440 335384 322446 335436
rect 335998 335384 336004 335436
rect 336056 335424 336062 335436
rect 349798 335424 349804 335436
rect 336056 335396 349804 335424
rect 336056 335384 336062 335396
rect 349798 335384 349804 335396
rect 349856 335384 349862 335436
rect 359642 335384 359648 335436
rect 359700 335424 359706 335436
rect 376294 335424 376300 335436
rect 359700 335396 376300 335424
rect 359700 335384 359706 335396
rect 376294 335384 376300 335396
rect 376352 335384 376358 335436
rect 386506 335384 386512 335436
rect 386564 335424 386570 335436
rect 403342 335424 403348 335436
rect 386564 335396 403348 335424
rect 386564 335384 386570 335396
rect 403342 335384 403348 335396
rect 403400 335384 403406 335436
rect 421282 335384 421288 335436
rect 421340 335424 421346 335436
rect 446398 335424 446404 335436
rect 421340 335396 446404 335424
rect 421340 335384 421346 335396
rect 446398 335384 446404 335396
rect 446456 335384 446462 335436
rect 494514 335384 494520 335436
rect 494572 335424 494578 335436
rect 511350 335424 511356 335436
rect 494572 335396 511356 335424
rect 494572 335384 494578 335396
rect 511350 335384 511356 335396
rect 511408 335384 511414 335436
rect 522298 335384 522304 335436
rect 522356 335424 522362 335436
rect 538398 335424 538404 335436
rect 522356 335396 538404 335424
rect 522356 335384 522362 335396
rect 538398 335384 538404 335396
rect 538456 335384 538462 335436
rect 43346 335316 43352 335368
rect 43404 335356 43410 335368
rect 62758 335356 62764 335368
rect 43404 335328 62764 335356
rect 43404 335316 43410 335328
rect 62758 335316 62764 335328
rect 62816 335316 62822 335368
rect 144178 335316 144184 335368
rect 144236 335356 144242 335368
rect 160278 335356 160284 335368
rect 144236 335328 160284 335356
rect 144236 335316 144242 335328
rect 160278 335316 160284 335328
rect 160336 335316 160342 335368
rect 171778 335316 171784 335368
rect 171836 335356 171842 335368
rect 197446 335356 197452 335368
rect 171836 335328 197452 335356
rect 171836 335316 171842 335328
rect 197446 335316 197452 335328
rect 197504 335316 197510 335368
rect 199378 335316 199384 335368
rect 199436 335356 199442 335368
rect 223942 335356 223948 335368
rect 199436 335328 223948 335356
rect 199436 335316 199442 335328
rect 223942 335316 223948 335328
rect 224000 335316 224006 335368
rect 225598 335316 225604 335368
rect 225656 335356 225662 335368
rect 251266 335356 251272 335368
rect 225656 335328 251272 335356
rect 225656 335316 225662 335328
rect 251266 335316 251272 335328
rect 251324 335316 251330 335368
rect 253198 335316 253204 335368
rect 253256 335356 253262 335368
rect 278038 335356 278044 335368
rect 253256 335328 278044 335356
rect 253256 335316 253262 335328
rect 278038 335316 278044 335328
rect 278096 335316 278102 335368
rect 279418 335316 279424 335368
rect 279476 335356 279482 335368
rect 305454 335356 305460 335368
rect 279476 335328 305460 335356
rect 279476 335316 279482 335328
rect 305454 335316 305460 335328
rect 305512 335316 305518 335368
rect 307018 335316 307024 335368
rect 307076 335356 307082 335368
rect 331950 335356 331956 335368
rect 307076 335328 331956 335356
rect 307076 335316 307082 335328
rect 331950 335316 331956 335328
rect 332008 335316 332014 335368
rect 333238 335316 333244 335368
rect 333296 335356 333302 335368
rect 359458 335356 359464 335368
rect 333296 335328 359464 335356
rect 333296 335316 333302 335328
rect 359458 335316 359464 335328
rect 359516 335316 359522 335368
rect 359550 335316 359556 335368
rect 359608 335356 359614 335368
rect 386046 335356 386052 335368
rect 359608 335328 386052 335356
rect 359608 335316 359614 335328
rect 386046 335316 386052 335328
rect 386104 335316 386110 335368
rect 387058 335316 387064 335368
rect 387116 335356 387122 335368
rect 412910 335356 412916 335368
rect 387116 335328 412916 335356
rect 387116 335316 387122 335328
rect 412910 335316 412916 335328
rect 412968 335316 412974 335368
rect 414658 335316 414664 335368
rect 414716 335356 414722 335368
rect 440234 335356 440240 335368
rect 414716 335328 440240 335356
rect 414716 335316 414722 335328
rect 440234 335316 440240 335328
rect 440292 335316 440298 335368
rect 442258 335316 442264 335368
rect 442316 335356 442322 335368
rect 467006 335356 467012 335368
rect 442316 335328 467012 335356
rect 442316 335316 442322 335328
rect 467006 335316 467012 335328
rect 467064 335316 467070 335368
rect 468570 335316 468576 335368
rect 468628 335356 468634 335368
rect 494054 335356 494060 335368
rect 468628 335328 494060 335356
rect 468628 335316 468634 335328
rect 494054 335316 494060 335328
rect 494112 335316 494118 335368
rect 496078 335316 496084 335368
rect 496136 335356 496142 335368
rect 520918 335356 520924 335368
rect 496136 335328 520924 335356
rect 496136 335316 496142 335328
rect 520918 335316 520924 335328
rect 520976 335316 520982 335368
rect 522390 335316 522396 335368
rect 522448 335356 522454 335368
rect 547966 335356 547972 335368
rect 522448 335328 547972 335356
rect 522448 335316 522454 335328
rect 547966 335316 547972 335328
rect 548024 335316 548030 335368
rect 37918 333208 37924 333260
rect 37976 333248 37982 333260
rect 526438 333248 526444 333260
rect 37976 333220 526444 333248
rect 37976 333208 37982 333220
rect 526438 333208 526444 333220
rect 526496 333208 526502 333260
rect 35618 332528 35624 332580
rect 35676 332568 35682 332580
rect 36630 332568 36636 332580
rect 35676 332540 36636 332568
rect 35676 332528 35682 332540
rect 36630 332528 36636 332540
rect 36688 332528 36694 332580
rect 285766 332256 285772 332308
rect 285824 332296 285830 332308
rect 286134 332296 286140 332308
rect 285824 332268 286140 332296
rect 285824 332256 285830 332268
rect 286134 332256 286140 332268
rect 286192 332256 286198 332308
rect 339586 332256 339592 332308
rect 339644 332296 339650 332308
rect 340138 332296 340144 332308
rect 339644 332268 340144 332296
rect 339644 332256 339650 332268
rect 340138 332256 340144 332268
rect 340196 332256 340202 332308
rect 359550 330624 359556 330676
rect 359608 330624 359614 330676
rect 359568 330472 359596 330624
rect 359550 330420 359556 330472
rect 359608 330420 359614 330472
rect 445662 314644 445668 314696
rect 445720 314684 445726 314696
rect 445720 314656 454034 314684
rect 445720 314644 445726 314656
rect 13722 314576 13728 314628
rect 13780 314616 13786 314628
rect 64874 314616 64880 314628
rect 13780 314588 64880 314616
rect 13780 314576 13786 314588
rect 64874 314576 64880 314588
rect 64932 314576 64938 314628
rect 89714 314576 89720 314628
rect 89772 314616 89778 314628
rect 90450 314616 90456 314628
rect 89772 314588 90456 314616
rect 89772 314576 89778 314588
rect 90450 314576 90456 314588
rect 90508 314576 90514 314628
rect 95142 314576 95148 314628
rect 95200 314616 95206 314628
rect 146294 314616 146300 314628
rect 95200 314588 146300 314616
rect 95200 314576 95206 314588
rect 146294 314576 146300 314588
rect 146352 314576 146358 314628
rect 148962 314576 148968 314628
rect 149020 314616 149026 314628
rect 200114 314616 200120 314628
rect 149020 314588 200120 314616
rect 149020 314576 149026 314588
rect 200114 314576 200120 314588
rect 200172 314576 200178 314628
rect 202782 314576 202788 314628
rect 202840 314616 202846 314628
rect 253934 314616 253940 314628
rect 202840 314588 253940 314616
rect 202840 314576 202846 314588
rect 253934 314576 253940 314588
rect 253992 314576 253998 314628
rect 256602 314576 256608 314628
rect 256660 314616 256666 314628
rect 307754 314616 307760 314628
rect 256660 314588 307760 314616
rect 256660 314576 256666 314588
rect 307754 314576 307760 314588
rect 307812 314576 307818 314628
rect 338022 314576 338028 314628
rect 338080 314616 338086 314628
rect 389174 314616 389180 314628
rect 338080 314588 389180 314616
rect 338080 314576 338086 314588
rect 389174 314576 389180 314588
rect 389232 314576 389238 314628
rect 391842 314576 391848 314628
rect 391900 314616 391906 314628
rect 442994 314616 443000 314628
rect 391900 314588 443000 314616
rect 391900 314576 391906 314588
rect 442994 314576 443000 314588
rect 443052 314576 443058 314628
rect 446398 314576 446404 314628
rect 446456 314616 446462 314628
rect 447686 314616 447692 314628
rect 446456 314588 447692 314616
rect 446456 314576 446462 314588
rect 447686 314576 447692 314588
rect 447744 314576 447750 314628
rect 454006 314616 454034 314656
rect 496814 314616 496820 314628
rect 454006 314588 496820 314616
rect 496814 314576 496820 314588
rect 496872 314576 496878 314628
rect 500862 314576 500868 314628
rect 500920 314616 500926 314628
rect 550634 314616 550640 314628
rect 500920 314588 550640 314616
rect 500920 314576 500926 314588
rect 550634 314576 550640 314588
rect 550692 314576 550698 314628
rect 41322 314508 41328 314560
rect 41380 314548 41386 314560
rect 91094 314548 91100 314560
rect 41380 314520 91100 314548
rect 41380 314508 41386 314520
rect 91094 314508 91100 314520
rect 91152 314508 91158 314560
rect 122742 314508 122748 314560
rect 122800 314548 122806 314560
rect 172514 314548 172520 314560
rect 122800 314520 172520 314548
rect 122800 314508 122806 314520
rect 172514 314508 172520 314520
rect 172572 314508 172578 314560
rect 176562 314508 176568 314560
rect 176620 314548 176626 314560
rect 226334 314548 226340 314560
rect 176620 314520 226340 314548
rect 176620 314508 176626 314520
rect 226334 314508 226340 314520
rect 226392 314508 226398 314560
rect 230382 314508 230388 314560
rect 230440 314548 230446 314560
rect 280154 314548 280160 314560
rect 230440 314520 280160 314548
rect 230440 314508 230446 314520
rect 280154 314508 280160 314520
rect 280212 314508 280218 314560
rect 284202 314508 284208 314560
rect 284260 314548 284266 314560
rect 335354 314548 335360 314560
rect 284260 314520 335360 314548
rect 284260 314508 284266 314520
rect 335354 314508 335360 314520
rect 335412 314508 335418 314560
rect 365622 314508 365628 314560
rect 365680 314548 365686 314560
rect 415394 314548 415400 314560
rect 365680 314520 415400 314548
rect 365680 314508 365686 314520
rect 415394 314508 415400 314520
rect 415452 314508 415458 314560
rect 419442 314508 419448 314560
rect 419500 314548 419506 314560
rect 469214 314548 469220 314560
rect 419500 314520 444374 314548
rect 419500 314508 419506 314520
rect 68922 314440 68928 314492
rect 68980 314480 68986 314492
rect 118694 314480 118700 314492
rect 68980 314452 118700 314480
rect 68980 314440 68986 314452
rect 118694 314440 118700 314452
rect 118752 314440 118758 314492
rect 278682 314440 278688 314492
rect 278740 314480 278746 314492
rect 279510 314480 279516 314492
rect 278740 314452 279516 314480
rect 278740 314440 278746 314452
rect 279510 314440 279516 314452
rect 279568 314440 279574 314492
rect 311802 314440 311808 314492
rect 311860 314480 311866 314492
rect 361574 314480 361580 314492
rect 311860 314452 361580 314480
rect 311860 314440 311866 314452
rect 361574 314440 361580 314452
rect 361632 314440 361638 314492
rect 444346 314412 444374 314520
rect 454006 314520 469220 314548
rect 454006 314412 454034 314520
rect 469214 314508 469220 314520
rect 469272 314508 469278 314560
rect 473262 314508 473268 314560
rect 473320 314548 473326 314560
rect 523034 314548 523040 314560
rect 473320 314520 523040 314548
rect 473320 314508 473326 314520
rect 523034 314508 523040 314520
rect 523092 314508 523098 314560
rect 444346 314384 454034 314412
rect 170214 313624 170220 313676
rect 170272 313664 170278 313676
rect 170490 313664 170496 313676
rect 170272 313636 170496 313664
rect 170272 313624 170278 313636
rect 170490 313624 170496 313636
rect 170548 313624 170554 313676
rect 62758 311788 62764 311840
rect 62816 311828 62822 311840
rect 69750 311828 69756 311840
rect 62816 311800 69756 311828
rect 62816 311788 62822 311800
rect 69750 311788 69756 311800
rect 69808 311788 69814 311840
rect 96706 311788 96712 311840
rect 96764 311828 96770 311840
rect 96764 311800 103514 311828
rect 96764 311788 96770 311800
rect 15194 311720 15200 311772
rect 15252 311760 15258 311772
rect 42794 311760 42800 311772
rect 15252 311732 42800 311760
rect 15252 311720 15258 311732
rect 42794 311720 42800 311732
rect 42852 311720 42858 311772
rect 53098 311720 53104 311772
rect 53156 311760 53162 311772
rect 64138 311760 64144 311772
rect 53156 311732 64144 311760
rect 53156 311720 53162 311732
rect 64138 311720 64144 311732
rect 64196 311720 64202 311772
rect 69106 311720 69112 311772
rect 69164 311760 69170 311772
rect 96798 311760 96804 311772
rect 69164 311732 96804 311760
rect 69164 311720 69170 311732
rect 96798 311720 96804 311732
rect 96856 311720 96862 311772
rect 103486 311760 103514 311800
rect 200758 311788 200764 311840
rect 200816 311828 200822 311840
rect 204622 311828 204628 311840
rect 200816 311800 204628 311828
rect 200816 311788 200822 311800
rect 204622 311788 204628 311800
rect 204680 311788 204686 311840
rect 251818 311788 251824 311840
rect 251876 311828 251882 311840
rect 258718 311828 258724 311840
rect 251876 311800 258724 311828
rect 251876 311788 251882 311800
rect 258718 311788 258724 311800
rect 258776 311788 258782 311840
rect 332502 311788 332508 311840
rect 332560 311828 332566 311840
rect 335998 311828 336004 311840
rect 332560 311800 336004 311828
rect 332560 311788 332566 311800
rect 335998 311788 336004 311800
rect 336056 311788 336062 311840
rect 494698 311788 494704 311840
rect 494756 311828 494762 311840
rect 501598 311828 501604 311840
rect 494756 311800 501604 311828
rect 494756 311788 494762 311800
rect 501598 311788 501604 311800
rect 501656 311788 501662 311840
rect 123662 311760 123668 311772
rect 103486 311732 123668 311760
rect 123662 311720 123668 311732
rect 123720 311720 123726 311772
rect 149698 311720 149704 311772
rect 149756 311760 149762 311772
rect 548058 311760 548064 311772
rect 149756 311732 548064 311760
rect 149756 311720 149762 311732
rect 548058 311720 548064 311732
rect 548116 311720 548122 311772
rect 25958 311652 25964 311704
rect 26016 311692 26022 311704
rect 36814 311692 36820 311704
rect 26016 311664 36820 311692
rect 26016 311652 26022 311664
rect 36814 311652 36820 311664
rect 36872 311652 36878 311704
rect 79962 311652 79968 311704
rect 80020 311692 80026 311704
rect 90358 311692 90364 311704
rect 80020 311664 90364 311692
rect 80020 311652 80026 311664
rect 90358 311652 90364 311664
rect 90416 311652 90422 311704
rect 106550 311652 106556 311704
rect 106608 311692 106614 311704
rect 116578 311692 116584 311704
rect 106608 311664 116584 311692
rect 106608 311652 106614 311664
rect 116578 311652 116584 311664
rect 116636 311652 116642 311704
rect 133782 311652 133788 311704
rect 133840 311692 133846 311704
rect 144270 311692 144276 311704
rect 133840 311664 144276 311692
rect 133840 311652 133846 311664
rect 144270 311652 144276 311664
rect 144328 311652 144334 311704
rect 150526 311652 150532 311704
rect 150584 311692 150590 311704
rect 178126 311692 178132 311704
rect 150584 311664 178132 311692
rect 150584 311652 150590 311664
rect 178126 311652 178132 311664
rect 178184 311652 178190 311704
rect 187970 311652 187976 311704
rect 188028 311692 188034 311704
rect 199378 311692 199384 311704
rect 188028 311664 199384 311692
rect 188028 311652 188034 311664
rect 199378 311652 199384 311664
rect 199436 311652 199442 311704
rect 204346 311652 204352 311704
rect 204404 311692 204410 311704
rect 231854 311692 231860 311704
rect 204404 311664 231860 311692
rect 204404 311652 204410 311664
rect 231854 311652 231860 311664
rect 231912 311652 231918 311704
rect 242066 311652 242072 311704
rect 242124 311692 242130 311704
rect 253198 311692 253204 311704
rect 242124 311664 253204 311692
rect 242124 311652 242130 311664
rect 253198 311652 253204 311664
rect 253256 311652 253262 311704
rect 258166 311652 258172 311704
rect 258224 311692 258230 311704
rect 286134 311692 286140 311704
rect 258224 311664 286140 311692
rect 258224 311652 258230 311664
rect 286134 311652 286140 311664
rect 286192 311652 286198 311704
rect 312630 311692 312636 311704
rect 287026 311664 312636 311692
rect 122926 311584 122932 311636
rect 122984 311624 122990 311636
rect 150710 311624 150716 311636
rect 122984 311596 150716 311624
rect 122984 311584 122990 311596
rect 150710 311584 150716 311596
rect 150768 311584 150774 311636
rect 160554 311584 160560 311636
rect 160612 311624 160618 311636
rect 171778 311624 171784 311636
rect 160612 311596 171784 311624
rect 160612 311584 160618 311596
rect 171778 311584 171784 311596
rect 171836 311584 171842 311636
rect 215018 311584 215024 311636
rect 215076 311624 215082 311636
rect 225598 311624 225604 311636
rect 215076 311596 225604 311624
rect 215076 311584 215082 311596
rect 225598 311584 225604 311596
rect 225656 311584 225662 311636
rect 268930 311584 268936 311636
rect 268988 311624 268994 311636
rect 279418 311624 279424 311636
rect 268988 311596 279424 311624
rect 268988 311584 268994 311596
rect 279418 311584 279424 311596
rect 279476 311584 279482 311636
rect 285766 311584 285772 311636
rect 285824 311624 285830 311636
rect 287026 311624 287054 311664
rect 312630 311652 312636 311664
rect 312688 311652 312694 311704
rect 340138 311692 340144 311704
rect 316006 311664 340144 311692
rect 285824 311596 287054 311624
rect 285824 311584 285830 311596
rect 295978 311584 295984 311636
rect 296036 311624 296042 311636
rect 307018 311624 307024 311636
rect 296036 311596 307024 311624
rect 296036 311584 296042 311596
rect 307018 311584 307024 311596
rect 307076 311584 307082 311636
rect 311986 311584 311992 311636
rect 312044 311624 312050 311636
rect 316006 311624 316034 311664
rect 340138 311652 340144 311664
rect 340196 311652 340202 311704
rect 366726 311692 366732 311704
rect 344986 311664 366732 311692
rect 312044 311596 316034 311624
rect 312044 311584 312050 311596
rect 322842 311584 322848 311636
rect 322900 311624 322906 311636
rect 333238 311624 333244 311636
rect 322900 311596 333244 311624
rect 322900 311584 322906 311596
rect 333238 311584 333244 311596
rect 333296 311584 333302 311636
rect 339586 311584 339592 311636
rect 339644 311624 339650 311636
rect 344986 311624 345014 311664
rect 366726 311652 366732 311664
rect 366784 311652 366790 311704
rect 393590 311692 393596 311704
rect 373966 311664 393596 311692
rect 339644 311596 345014 311624
rect 339644 311584 339650 311596
rect 350074 311584 350080 311636
rect 350132 311624 350138 311636
rect 359550 311624 359556 311636
rect 350132 311596 359556 311624
rect 350132 311584 350138 311596
rect 359550 311584 359556 311596
rect 359608 311584 359614 311636
rect 365806 311584 365812 311636
rect 365864 311624 365870 311636
rect 373966 311624 373994 311664
rect 393590 311652 393596 311664
rect 393648 311652 393654 311704
rect 420914 311692 420920 311704
rect 402946 311664 420920 311692
rect 365864 311596 373994 311624
rect 365864 311584 365870 311596
rect 376570 311584 376576 311636
rect 376628 311624 376634 311636
rect 387058 311624 387064 311636
rect 376628 311596 387064 311624
rect 376628 311584 376634 311596
rect 387058 311584 387064 311596
rect 387116 311584 387122 311636
rect 393406 311584 393412 311636
rect 393464 311624 393470 311636
rect 402946 311624 402974 311664
rect 420914 311652 420920 311664
rect 420972 311652 420978 311704
rect 431034 311652 431040 311704
rect 431092 311692 431098 311704
rect 442258 311692 442264 311704
rect 431092 311664 442264 311692
rect 431092 311652 431098 311664
rect 442258 311652 442264 311664
rect 442316 311652 442322 311704
rect 447226 311652 447232 311704
rect 447284 311692 447290 311704
rect 474734 311692 474740 311704
rect 447284 311664 474740 311692
rect 447284 311652 447290 311664
rect 474734 311652 474740 311664
rect 474792 311652 474798 311704
rect 484946 311652 484952 311704
rect 485004 311692 485010 311704
rect 496078 311692 496084 311704
rect 485004 311664 496084 311692
rect 485004 311652 485010 311664
rect 496078 311652 496084 311664
rect 496136 311652 496142 311704
rect 501046 311652 501052 311704
rect 501104 311692 501110 311704
rect 528738 311692 528744 311704
rect 501104 311664 528744 311692
rect 501104 311652 501110 311664
rect 528738 311652 528744 311664
rect 528796 311652 528802 311704
rect 393464 311596 402974 311624
rect 393464 311584 393470 311596
rect 403986 311584 403992 311636
rect 404044 311624 404050 311636
rect 414658 311624 414664 311636
rect 404044 311596 414664 311624
rect 404044 311584 404050 311596
rect 414658 311584 414664 311596
rect 414716 311584 414722 311636
rect 458082 311584 458088 311636
rect 458140 311624 458146 311636
rect 468570 311624 468576 311636
rect 458140 311596 468576 311624
rect 458140 311584 458146 311596
rect 468570 311584 468576 311596
rect 468628 311584 468634 311636
rect 511902 311584 511908 311636
rect 511960 311624 511966 311636
rect 522390 311624 522396 311636
rect 511960 311596 522396 311624
rect 511960 311584 511966 311596
rect 522390 311584 522396 311596
rect 522448 311584 522454 311636
rect 36722 311516 36728 311568
rect 36780 311556 36786 311568
rect 538398 311556 538404 311568
rect 36780 311528 538404 311556
rect 36780 311516 36786 311528
rect 538398 311516 538404 311528
rect 538456 311516 538462 311568
rect 16298 308388 16304 308440
rect 16356 308428 16362 308440
rect 529014 308428 529020 308440
rect 16356 308400 529020 308428
rect 16356 308388 16362 308400
rect 529014 308388 529020 308400
rect 529072 308388 529078 308440
rect 25682 308048 25688 308100
rect 25740 308088 25746 308100
rect 149698 308088 149704 308100
rect 25740 308060 149704 308088
rect 25740 308048 25746 308060
rect 149698 308048 149704 308060
rect 149756 308048 149762 308100
rect 36814 307980 36820 308032
rect 36872 308020 36878 308032
rect 52638 308020 52644 308032
rect 36872 307992 52644 308020
rect 36872 307980 36878 307992
rect 52638 307980 52644 307992
rect 52696 307980 52702 308032
rect 232038 307980 232044 308032
rect 232096 308020 232102 308032
rect 251818 308020 251824 308032
rect 232096 307992 251824 308020
rect 232096 307980 232102 307992
rect 251818 307980 251824 307992
rect 251876 307980 251882 308032
rect 475010 307980 475016 308032
rect 475068 308020 475074 308032
rect 494698 308020 494704 308032
rect 475068 307992 494704 308020
rect 475068 307980 475074 307992
rect 494698 307980 494704 307992
rect 494756 307980 494762 308032
rect 62482 307912 62488 307964
rect 62540 307952 62546 307964
rect 79686 307952 79692 307964
rect 62540 307924 79692 307952
rect 62540 307912 62546 307924
rect 79686 307912 79692 307924
rect 79744 307912 79750 307964
rect 90358 307912 90364 307964
rect 90416 307952 90422 307964
rect 106642 307952 106648 307964
rect 90416 307924 106648 307952
rect 90416 307912 90422 307924
rect 106642 307912 106648 307924
rect 106700 307912 106706 307964
rect 116486 307912 116492 307964
rect 116544 307952 116550 307964
rect 133690 307952 133696 307964
rect 116544 307924 133696 307952
rect 116544 307912 116550 307924
rect 133690 307912 133696 307924
rect 133748 307912 133754 307964
rect 144178 307912 144184 307964
rect 144236 307952 144242 307964
rect 160646 307952 160652 307964
rect 144236 307924 160652 307952
rect 144236 307912 144242 307924
rect 160646 307912 160652 307924
rect 160704 307912 160710 307964
rect 170490 307912 170496 307964
rect 170548 307952 170554 307964
rect 187694 307952 187700 307964
rect 170548 307924 187700 307952
rect 170548 307912 170554 307924
rect 187694 307912 187700 307924
rect 187752 307912 187758 307964
rect 197446 307912 197452 307964
rect 197504 307952 197510 307964
rect 214650 307952 214656 307964
rect 197504 307924 214656 307952
rect 197504 307912 197510 307924
rect 214650 307912 214656 307924
rect 214708 307912 214714 307964
rect 224494 307912 224500 307964
rect 224552 307952 224558 307964
rect 241698 307952 241704 307964
rect 224552 307924 241704 307952
rect 224552 307912 224558 307924
rect 241698 307912 241704 307924
rect 241756 307912 241762 307964
rect 413462 307912 413468 307964
rect 413520 307952 413526 307964
rect 430666 307952 430672 307964
rect 413520 307924 430672 307952
rect 413520 307912 413526 307924
rect 430666 307912 430672 307924
rect 430724 307912 430730 307964
rect 440510 307912 440516 307964
rect 440568 307952 440574 307964
rect 457622 307952 457628 307964
rect 440568 307924 457628 307952
rect 440568 307912 440574 307924
rect 457622 307912 457628 307924
rect 457680 307912 457686 307964
rect 468570 307912 468576 307964
rect 468628 307952 468634 307964
rect 484670 307952 484676 307964
rect 468628 307924 484676 307952
rect 468628 307912 468634 307924
rect 484670 307912 484676 307924
rect 484728 307912 484734 307964
rect 36722 307844 36728 307896
rect 36780 307884 36786 307896
rect 62298 307884 62304 307896
rect 36780 307856 62304 307884
rect 36780 307844 36786 307856
rect 62298 307844 62304 307856
rect 62356 307844 62362 307896
rect 64138 307844 64144 307896
rect 64196 307884 64202 307896
rect 89346 307884 89352 307896
rect 64196 307856 89352 307884
rect 64196 307844 64202 307856
rect 89346 307844 89352 307856
rect 89404 307844 89410 307896
rect 90450 307844 90456 307896
rect 90508 307884 90514 307896
rect 116302 307884 116308 307896
rect 90508 307856 116308 307884
rect 90508 307844 90514 307856
rect 116302 307844 116308 307856
rect 116360 307844 116366 307896
rect 116578 307844 116584 307896
rect 116636 307884 116642 307896
rect 143350 307884 143356 307896
rect 116636 307856 143356 307884
rect 116636 307844 116642 307856
rect 143350 307844 143356 307856
rect 143408 307844 143414 307896
rect 144270 307844 144276 307896
rect 144328 307884 144334 307896
rect 170306 307884 170312 307896
rect 144328 307856 170312 307884
rect 144328 307844 144334 307856
rect 170306 307844 170312 307856
rect 170364 307844 170370 307896
rect 178034 307844 178040 307896
rect 178092 307884 178098 307896
rect 200758 307884 200764 307896
rect 178092 307856 200764 307884
rect 178092 307844 178098 307856
rect 200758 307844 200764 307856
rect 200816 307844 200822 307896
rect 251450 307844 251456 307896
rect 251508 307884 251514 307896
rect 268654 307884 268660 307896
rect 251508 307856 268660 307884
rect 251508 307844 251514 307856
rect 268654 307844 268660 307856
rect 268712 307844 268718 307896
rect 279510 307844 279516 307896
rect 279568 307884 279574 307896
rect 295702 307884 295708 307896
rect 279568 307856 295708 307884
rect 279568 307844 279574 307856
rect 295702 307844 295708 307856
rect 295760 307844 295766 307896
rect 305454 307844 305460 307896
rect 305512 307884 305518 307896
rect 322658 307884 322664 307896
rect 305512 307856 322664 307884
rect 305512 307844 305518 307856
rect 322658 307844 322664 307856
rect 322716 307844 322722 307896
rect 334618 307844 334624 307896
rect 334676 307884 334682 307896
rect 349706 307884 349712 307896
rect 334676 307856 349712 307884
rect 334676 307844 334682 307856
rect 349706 307844 349712 307856
rect 349764 307844 349770 307896
rect 359458 307844 359464 307896
rect 359516 307884 359522 307896
rect 376662 307884 376668 307896
rect 359516 307856 376668 307884
rect 359516 307844 359522 307856
rect 376662 307844 376668 307856
rect 376720 307844 376726 307896
rect 386506 307844 386512 307896
rect 386564 307884 386570 307896
rect 403618 307884 403624 307896
rect 386564 307856 403624 307884
rect 386564 307844 386570 307856
rect 403618 307844 403624 307856
rect 403676 307844 403682 307896
rect 421006 307844 421012 307896
rect 421064 307884 421070 307896
rect 443638 307884 443644 307896
rect 421064 307856 443644 307884
rect 421064 307844 421070 307856
rect 443638 307844 443644 307856
rect 443696 307844 443702 307896
rect 494514 307844 494520 307896
rect 494572 307884 494578 307896
rect 511626 307884 511632 307896
rect 494572 307856 511632 307884
rect 494572 307844 494578 307856
rect 511626 307844 511632 307856
rect 511684 307844 511690 307896
rect 522298 307844 522304 307896
rect 522356 307884 522362 307896
rect 538674 307884 538680 307896
rect 522356 307856 538680 307884
rect 522356 307844 522362 307856
rect 538674 307844 538680 307856
rect 538732 307844 538738 307896
rect 43070 307776 43076 307828
rect 43128 307816 43134 307828
rect 62758 307816 62764 307828
rect 43128 307788 62764 307816
rect 43128 307776 43134 307788
rect 62758 307776 62764 307788
rect 62816 307776 62822 307828
rect 171778 307776 171784 307828
rect 171836 307816 171842 307828
rect 197354 307816 197360 307828
rect 171836 307788 197360 307816
rect 171836 307776 171842 307788
rect 197354 307776 197360 307788
rect 197412 307776 197418 307828
rect 199378 307776 199384 307828
rect 199436 307816 199442 307828
rect 224310 307816 224316 307828
rect 199436 307788 224316 307816
rect 199436 307776 199442 307788
rect 224310 307776 224316 307788
rect 224368 307776 224374 307828
rect 225598 307776 225604 307828
rect 225656 307816 225662 307828
rect 251358 307816 251364 307828
rect 225656 307788 251364 307816
rect 225656 307776 225662 307788
rect 251358 307776 251364 307788
rect 251416 307776 251422 307828
rect 253198 307776 253204 307828
rect 253256 307816 253262 307828
rect 278314 307816 278320 307828
rect 253256 307788 278320 307816
rect 253256 307776 253262 307788
rect 278314 307776 278320 307788
rect 278372 307776 278378 307828
rect 279418 307776 279424 307828
rect 279476 307816 279482 307828
rect 305362 307816 305368 307828
rect 279476 307788 305368 307816
rect 279476 307776 279482 307788
rect 305362 307776 305368 307788
rect 305420 307776 305426 307828
rect 307018 307776 307024 307828
rect 307076 307816 307082 307828
rect 332318 307816 332324 307828
rect 307076 307788 332324 307816
rect 307076 307776 307082 307788
rect 332318 307776 332324 307788
rect 332376 307776 332382 307828
rect 333238 307776 333244 307828
rect 333296 307816 333302 307828
rect 359366 307816 359372 307828
rect 333296 307788 359372 307816
rect 333296 307776 333302 307788
rect 359366 307776 359372 307788
rect 359424 307776 359430 307828
rect 359550 307776 359556 307828
rect 359608 307816 359614 307828
rect 386322 307816 386328 307828
rect 359608 307788 386328 307816
rect 359608 307776 359614 307788
rect 386322 307776 386328 307788
rect 386380 307776 386386 307828
rect 387058 307776 387064 307828
rect 387116 307816 387122 307828
rect 413278 307816 413284 307828
rect 387116 307788 413284 307816
rect 387116 307776 387122 307788
rect 413278 307776 413284 307788
rect 413336 307776 413342 307828
rect 414658 307776 414664 307828
rect 414716 307816 414722 307828
rect 440326 307816 440332 307828
rect 414716 307788 440332 307816
rect 414716 307776 414722 307788
rect 440326 307776 440332 307788
rect 440384 307776 440390 307828
rect 442258 307776 442264 307828
rect 442316 307816 442322 307828
rect 467282 307816 467288 307828
rect 442316 307788 467288 307816
rect 442316 307776 442322 307788
rect 467282 307776 467288 307788
rect 467340 307776 467346 307828
rect 468478 307776 468484 307828
rect 468536 307816 468542 307828
rect 494330 307816 494336 307828
rect 468536 307788 494336 307816
rect 468536 307776 468542 307788
rect 494330 307776 494336 307788
rect 494388 307776 494394 307828
rect 496078 307776 496084 307828
rect 496136 307816 496142 307828
rect 521286 307816 521292 307828
rect 496136 307788 521292 307816
rect 496136 307776 496142 307788
rect 521286 307776 521292 307788
rect 521344 307776 521350 307828
rect 522390 307776 522396 307828
rect 522448 307816 522454 307828
rect 548334 307816 548340 307828
rect 522448 307788 548340 307816
rect 522448 307776 522454 307788
rect 548334 307776 548340 307788
rect 548392 307776 548398 307828
rect 37918 305600 37924 305652
rect 37976 305640 37982 305652
rect 526438 305640 526444 305652
rect 37976 305612 526444 305640
rect 37976 305600 37982 305612
rect 526438 305600 526444 305612
rect 526496 305600 526502 305652
rect 13722 286968 13728 287020
rect 13780 287008 13786 287020
rect 64874 287008 64880 287020
rect 13780 286980 64880 287008
rect 13780 286968 13786 286980
rect 64874 286968 64880 286980
rect 64932 286968 64938 287020
rect 95142 286968 95148 287020
rect 95200 287008 95206 287020
rect 146294 287008 146300 287020
rect 95200 286980 146300 287008
rect 95200 286968 95206 286980
rect 146294 286968 146300 286980
rect 146352 286968 146358 287020
rect 148962 286968 148968 287020
rect 149020 287008 149026 287020
rect 200114 287008 200120 287020
rect 149020 286980 200120 287008
rect 149020 286968 149026 286980
rect 200114 286968 200120 286980
rect 200172 286968 200178 287020
rect 202782 286968 202788 287020
rect 202840 287008 202846 287020
rect 253934 287008 253940 287020
rect 202840 286980 253940 287008
rect 202840 286968 202846 286980
rect 253934 286968 253940 286980
rect 253992 286968 253998 287020
rect 256602 286968 256608 287020
rect 256660 287008 256666 287020
rect 307754 287008 307760 287020
rect 256660 286980 307760 287008
rect 256660 286968 256666 286980
rect 307754 286968 307760 286980
rect 307812 286968 307818 287020
rect 338022 286968 338028 287020
rect 338080 287008 338086 287020
rect 389174 287008 389180 287020
rect 338080 286980 389180 287008
rect 338080 286968 338086 286980
rect 389174 286968 389180 286980
rect 389232 286968 389238 287020
rect 391842 286968 391848 287020
rect 391900 287008 391906 287020
rect 442994 287008 443000 287020
rect 391900 286980 443000 287008
rect 391900 286968 391906 286980
rect 442994 286968 443000 286980
rect 443052 286968 443058 287020
rect 445662 286968 445668 287020
rect 445720 287008 445726 287020
rect 496814 287008 496820 287020
rect 445720 286980 496820 287008
rect 445720 286968 445726 286980
rect 496814 286968 496820 286980
rect 496872 286968 496878 287020
rect 500862 286968 500868 287020
rect 500920 287008 500926 287020
rect 550634 287008 550640 287020
rect 500920 286980 550640 287008
rect 500920 286968 500926 286980
rect 550634 286968 550640 286980
rect 550692 286968 550698 287020
rect 35618 286900 35624 286952
rect 35676 286940 35682 286952
rect 36814 286940 36820 286952
rect 35676 286912 36820 286940
rect 35676 286900 35682 286912
rect 36814 286900 36820 286912
rect 36872 286900 36878 286952
rect 41322 286900 41328 286952
rect 41380 286940 41386 286952
rect 91094 286940 91100 286952
rect 41380 286912 91100 286940
rect 41380 286900 41386 286912
rect 91094 286900 91100 286912
rect 91152 286900 91158 286952
rect 122742 286900 122748 286952
rect 122800 286940 122806 286952
rect 172514 286940 172520 286952
rect 122800 286912 172520 286940
rect 122800 286900 122806 286912
rect 172514 286900 172520 286912
rect 172572 286900 172578 286952
rect 176562 286900 176568 286952
rect 176620 286940 176626 286952
rect 226334 286940 226340 286952
rect 176620 286912 226340 286940
rect 176620 286900 176626 286912
rect 226334 286900 226340 286912
rect 226392 286900 226398 286952
rect 230382 286900 230388 286952
rect 230440 286940 230446 286952
rect 280154 286940 280160 286952
rect 230440 286912 280160 286940
rect 230440 286900 230446 286912
rect 280154 286900 280160 286912
rect 280212 286900 280218 286952
rect 284202 286900 284208 286952
rect 284260 286940 284266 286952
rect 335354 286940 335360 286952
rect 284260 286912 335360 286940
rect 284260 286900 284266 286912
rect 335354 286900 335360 286912
rect 335412 286900 335418 286952
rect 365622 286900 365628 286952
rect 365680 286940 365686 286952
rect 415394 286940 415400 286952
rect 365680 286912 415400 286940
rect 365680 286900 365686 286912
rect 415394 286900 415400 286912
rect 415452 286900 415458 286952
rect 419442 286900 419448 286952
rect 419500 286940 419506 286952
rect 469214 286940 469220 286952
rect 419500 286912 469220 286940
rect 419500 286900 419506 286912
rect 469214 286900 469220 286912
rect 469272 286900 469278 286952
rect 473262 286900 473268 286952
rect 473320 286940 473326 286952
rect 523034 286940 523040 286952
rect 473320 286912 523040 286940
rect 473320 286900 473326 286912
rect 523034 286900 523040 286912
rect 523092 286900 523098 286952
rect 68922 286832 68928 286884
rect 68980 286872 68986 286884
rect 118694 286872 118700 286884
rect 68980 286844 118700 286872
rect 68980 286832 68986 286844
rect 118694 286832 118700 286844
rect 118752 286832 118758 286884
rect 311802 286832 311808 286884
rect 311860 286872 311866 286884
rect 361574 286872 361580 286884
rect 311860 286844 361580 286872
rect 311860 286832 311866 286844
rect 361574 286832 361580 286844
rect 361632 286832 361638 286884
rect 200758 286764 200764 286816
rect 200816 286804 200822 286816
rect 204622 286804 204628 286816
rect 200816 286776 204628 286804
rect 200816 286764 200822 286776
rect 204622 286764 204628 286776
rect 204680 286764 204686 286816
rect 278682 286764 278688 286816
rect 278740 286804 278746 286816
rect 279510 286804 279516 286816
rect 278740 286776 279516 286804
rect 278740 286764 278746 286776
rect 279510 286764 279516 286776
rect 279568 286764 279574 286816
rect 332502 286764 332508 286816
rect 332560 286804 332566 286816
rect 334618 286804 334624 286816
rect 332560 286776 334624 286804
rect 332560 286764 332566 286776
rect 334618 286764 334624 286776
rect 334676 286764 334682 286816
rect 467650 286764 467656 286816
rect 467708 286804 467714 286816
rect 468570 286804 468576 286816
rect 467708 286776 468576 286804
rect 467708 286764 467714 286776
rect 468570 286764 468576 286776
rect 468628 286764 468634 286816
rect 62758 284248 62764 284300
rect 62816 284288 62822 284300
rect 70026 284288 70032 284300
rect 62816 284260 70032 284288
rect 62816 284248 62822 284260
rect 70026 284248 70032 284260
rect 70084 284248 70090 284300
rect 96706 284248 96712 284300
rect 96764 284288 96770 284300
rect 96764 284260 103514 284288
rect 96764 284248 96770 284260
rect 15194 284180 15200 284232
rect 15252 284220 15258 284232
rect 42978 284220 42984 284232
rect 15252 284192 42984 284220
rect 15252 284180 15258 284192
rect 42978 284180 42984 284192
rect 43036 284180 43042 284232
rect 52730 284180 52736 284232
rect 52788 284220 52794 284232
rect 64138 284220 64144 284232
rect 52788 284192 64144 284220
rect 52788 284180 52794 284192
rect 64138 284180 64144 284192
rect 64196 284180 64202 284232
rect 69106 284180 69112 284232
rect 69164 284220 69170 284232
rect 96982 284220 96988 284232
rect 69164 284192 96988 284220
rect 69164 284180 69170 284192
rect 96982 284180 96988 284192
rect 97040 284180 97046 284232
rect 103486 284220 103514 284260
rect 146938 284248 146944 284300
rect 146996 284288 147002 284300
rect 146996 284260 151814 284288
rect 146996 284248 147002 284260
rect 124030 284220 124036 284232
rect 103486 284192 124036 284220
rect 124030 284180 124036 284192
rect 124088 284180 124094 284232
rect 133690 284180 133696 284232
rect 133748 284220 133754 284232
rect 144270 284220 144276 284232
rect 133748 284192 144276 284220
rect 133748 284180 133754 284192
rect 144270 284180 144276 284192
rect 144328 284180 144334 284232
rect 150526 284180 150532 284232
rect 150584 284220 150590 284232
rect 151786 284220 151814 284260
rect 251818 284248 251824 284300
rect 251876 284288 251882 284300
rect 258994 284288 259000 284300
rect 251876 284260 259000 284288
rect 251876 284248 251882 284260
rect 258994 284248 259000 284260
rect 259052 284248 259058 284300
rect 443638 284248 443644 284300
rect 443696 284288 443702 284300
rect 447962 284288 447968 284300
rect 443696 284260 447968 284288
rect 443696 284248 443702 284260
rect 447962 284248 447968 284260
rect 448020 284248 448026 284300
rect 494698 284248 494704 284300
rect 494756 284288 494762 284300
rect 501966 284288 501972 284300
rect 494756 284260 501972 284288
rect 494756 284248 494762 284260
rect 501966 284248 501972 284260
rect 502024 284248 502030 284300
rect 548334 284220 548340 284232
rect 150584 284192 151124 284220
rect 151786 284192 548340 284220
rect 150584 284180 150590 284192
rect 25682 284112 25688 284164
rect 25740 284152 25746 284164
rect 36722 284152 36728 284164
rect 25740 284124 36728 284152
rect 25740 284112 25746 284124
rect 36722 284112 36728 284124
rect 36780 284112 36786 284164
rect 79686 284112 79692 284164
rect 79744 284152 79750 284164
rect 90450 284152 90456 284164
rect 79744 284124 90456 284152
rect 79744 284112 79750 284124
rect 90450 284112 90456 284124
rect 90508 284112 90514 284164
rect 106642 284112 106648 284164
rect 106700 284152 106706 284164
rect 116578 284152 116584 284164
rect 106700 284124 116584 284152
rect 106700 284112 106706 284124
rect 116578 284112 116584 284124
rect 116636 284112 116642 284164
rect 122926 284112 122932 284164
rect 122984 284152 122990 284164
rect 150986 284152 150992 284164
rect 122984 284124 150992 284152
rect 122984 284112 122990 284124
rect 150986 284112 150992 284124
rect 151044 284112 151050 284164
rect 151096 284152 151124 284192
rect 548334 284180 548340 284192
rect 548392 284180 548398 284232
rect 178034 284152 178040 284164
rect 151096 284124 178040 284152
rect 178034 284112 178040 284124
rect 178092 284112 178098 284164
rect 187694 284112 187700 284164
rect 187752 284152 187758 284164
rect 199378 284152 199384 284164
rect 187752 284124 199384 284152
rect 187752 284112 187758 284124
rect 199378 284112 199384 284124
rect 199436 284112 199442 284164
rect 204346 284112 204352 284164
rect 204404 284152 204410 284164
rect 232038 284152 232044 284164
rect 204404 284124 232044 284152
rect 204404 284112 204410 284124
rect 232038 284112 232044 284124
rect 232096 284112 232102 284164
rect 241698 284112 241704 284164
rect 241756 284152 241762 284164
rect 253198 284152 253204 284164
rect 241756 284124 253204 284152
rect 241756 284112 241762 284124
rect 253198 284112 253204 284124
rect 253256 284112 253262 284164
rect 258166 284112 258172 284164
rect 258224 284152 258230 284164
rect 286042 284152 286048 284164
rect 258224 284124 286048 284152
rect 258224 284112 258230 284124
rect 286042 284112 286048 284124
rect 286100 284112 286106 284164
rect 312998 284152 313004 284164
rect 287026 284124 313004 284152
rect 160646 284044 160652 284096
rect 160704 284084 160710 284096
rect 171778 284084 171784 284096
rect 160704 284056 171784 284084
rect 160704 284044 160710 284056
rect 171778 284044 171784 284056
rect 171836 284044 171842 284096
rect 214650 284044 214656 284096
rect 214708 284084 214714 284096
rect 225598 284084 225604 284096
rect 214708 284056 225604 284084
rect 214708 284044 214714 284056
rect 225598 284044 225604 284056
rect 225656 284044 225662 284096
rect 268654 284044 268660 284096
rect 268712 284084 268718 284096
rect 279418 284084 279424 284096
rect 268712 284056 279424 284084
rect 268712 284044 268718 284056
rect 279418 284044 279424 284056
rect 279476 284044 279482 284096
rect 285766 284044 285772 284096
rect 285824 284084 285830 284096
rect 287026 284084 287054 284124
rect 312998 284112 313004 284124
rect 313056 284112 313062 284164
rect 340046 284152 340052 284164
rect 316006 284124 340052 284152
rect 285824 284056 287054 284084
rect 285824 284044 285830 284056
rect 295702 284044 295708 284096
rect 295760 284084 295766 284096
rect 307018 284084 307024 284096
rect 295760 284056 307024 284084
rect 295760 284044 295766 284056
rect 307018 284044 307024 284056
rect 307076 284044 307082 284096
rect 311986 284044 311992 284096
rect 312044 284084 312050 284096
rect 316006 284084 316034 284124
rect 340046 284112 340052 284124
rect 340104 284112 340110 284164
rect 367002 284152 367008 284164
rect 344986 284124 367008 284152
rect 312044 284056 316034 284084
rect 312044 284044 312050 284056
rect 322658 284044 322664 284096
rect 322716 284084 322722 284096
rect 333238 284084 333244 284096
rect 322716 284056 333244 284084
rect 322716 284044 322722 284056
rect 333238 284044 333244 284056
rect 333296 284044 333302 284096
rect 339586 284044 339592 284096
rect 339644 284084 339650 284096
rect 344986 284084 345014 284124
rect 367002 284112 367008 284124
rect 367060 284112 367066 284164
rect 393958 284152 393964 284164
rect 373966 284124 393964 284152
rect 339644 284056 345014 284084
rect 339644 284044 339650 284056
rect 349706 284044 349712 284096
rect 349764 284084 349770 284096
rect 359550 284084 359556 284096
rect 349764 284056 359556 284084
rect 349764 284044 349770 284056
rect 359550 284044 359556 284056
rect 359608 284044 359614 284096
rect 365806 284044 365812 284096
rect 365864 284084 365870 284096
rect 373966 284084 373994 284124
rect 393958 284112 393964 284124
rect 394016 284112 394022 284164
rect 421006 284152 421012 284164
rect 402946 284124 421012 284152
rect 365864 284056 373994 284084
rect 365864 284044 365870 284056
rect 376662 284044 376668 284096
rect 376720 284084 376726 284096
rect 387058 284084 387064 284096
rect 376720 284056 387064 284084
rect 376720 284044 376726 284056
rect 387058 284044 387064 284056
rect 387116 284044 387122 284096
rect 393406 284044 393412 284096
rect 393464 284084 393470 284096
rect 402946 284084 402974 284124
rect 421006 284112 421012 284124
rect 421064 284112 421070 284164
rect 430666 284112 430672 284164
rect 430724 284152 430730 284164
rect 442258 284152 442264 284164
rect 430724 284124 442264 284152
rect 430724 284112 430730 284124
rect 442258 284112 442264 284124
rect 442316 284112 442322 284164
rect 447226 284112 447232 284164
rect 447284 284152 447290 284164
rect 475010 284152 475016 284164
rect 447284 284124 475016 284152
rect 447284 284112 447290 284124
rect 475010 284112 475016 284124
rect 475068 284112 475074 284164
rect 484670 284112 484676 284164
rect 484728 284152 484734 284164
rect 496078 284152 496084 284164
rect 484728 284124 496084 284152
rect 484728 284112 484734 284124
rect 496078 284112 496084 284124
rect 496136 284112 496142 284164
rect 501046 284112 501052 284164
rect 501104 284152 501110 284164
rect 529014 284152 529020 284164
rect 501104 284124 529020 284152
rect 501104 284112 501110 284124
rect 529014 284112 529020 284124
rect 529072 284112 529078 284164
rect 393464 284056 402974 284084
rect 393464 284044 393470 284056
rect 403710 284044 403716 284096
rect 403768 284084 403774 284096
rect 414658 284084 414664 284096
rect 403768 284056 414664 284084
rect 403768 284044 403774 284056
rect 414658 284044 414664 284056
rect 414716 284044 414722 284096
rect 457714 284044 457720 284096
rect 457772 284084 457778 284096
rect 468478 284084 468484 284096
rect 457772 284056 468484 284084
rect 457772 284044 457778 284056
rect 468478 284044 468484 284056
rect 468536 284044 468542 284096
rect 511718 284044 511724 284096
rect 511776 284084 511782 284096
rect 522390 284084 522396 284096
rect 511776 284056 522396 284084
rect 511776 284044 511782 284056
rect 522390 284044 522396 284056
rect 522448 284044 522454 284096
rect 36630 283976 36636 284028
rect 36688 284016 36694 284028
rect 538674 284016 538680 284028
rect 36688 283988 538680 284016
rect 36688 283976 36694 283988
rect 538674 283976 538680 283988
rect 538732 283976 538738 284028
rect 16022 280780 16028 280832
rect 16080 280820 16086 280832
rect 528738 280820 528744 280832
rect 16080 280792 528744 280820
rect 16080 280780 16086 280792
rect 528738 280780 528744 280792
rect 528796 280780 528802 280832
rect 25958 280440 25964 280492
rect 26016 280480 26022 280492
rect 146938 280480 146944 280492
rect 26016 280452 146944 280480
rect 26016 280440 26022 280452
rect 146938 280440 146944 280452
rect 146996 280440 147002 280492
rect 36814 280372 36820 280424
rect 36872 280412 36878 280424
rect 52454 280412 52460 280424
rect 36872 280384 52460 280412
rect 36872 280372 36878 280384
rect 52454 280372 52460 280384
rect 52512 280372 52518 280424
rect 232314 280372 232320 280424
rect 232372 280412 232378 280424
rect 251818 280412 251824 280424
rect 232372 280384 251824 280412
rect 232372 280372 232378 280384
rect 251818 280372 251824 280384
rect 251876 280372 251882 280424
rect 475378 280372 475384 280424
rect 475436 280412 475442 280424
rect 494698 280412 494704 280424
rect 475436 280384 494704 280412
rect 475436 280372 475442 280384
rect 494698 280372 494704 280384
rect 494756 280372 494762 280424
rect 62482 280304 62488 280356
rect 62540 280344 62546 280356
rect 79318 280344 79324 280356
rect 62540 280316 79324 280344
rect 62540 280304 62546 280316
rect 79318 280304 79324 280316
rect 79376 280304 79382 280356
rect 90358 280304 90364 280356
rect 90416 280344 90422 280356
rect 106366 280344 106372 280356
rect 90416 280316 106372 280344
rect 90416 280304 90422 280316
rect 106366 280304 106372 280316
rect 106424 280304 106430 280356
rect 116486 280304 116492 280356
rect 116544 280344 116550 280356
rect 133414 280344 133420 280356
rect 116544 280316 133420 280344
rect 116544 280304 116550 280316
rect 133414 280304 133420 280316
rect 133472 280304 133478 280356
rect 170490 280304 170496 280356
rect 170548 280344 170554 280356
rect 187786 280344 187792 280356
rect 170548 280316 187792 280344
rect 170548 280304 170554 280316
rect 187786 280304 187792 280316
rect 187844 280304 187850 280356
rect 197538 280304 197544 280356
rect 197596 280344 197602 280356
rect 214374 280344 214380 280356
rect 197596 280316 214380 280344
rect 197596 280304 197602 280316
rect 214374 280304 214380 280316
rect 214432 280304 214438 280356
rect 224494 280304 224500 280356
rect 224552 280344 224558 280356
rect 241514 280344 241520 280356
rect 224552 280316 241520 280344
rect 224552 280304 224558 280316
rect 241514 280304 241520 280316
rect 241572 280304 241578 280356
rect 413462 280304 413468 280356
rect 413520 280344 413526 280356
rect 430574 280344 430580 280356
rect 413520 280316 430580 280344
rect 413520 280304 413526 280316
rect 430574 280304 430580 280316
rect 430632 280304 430638 280356
rect 440510 280304 440516 280356
rect 440568 280344 440574 280356
rect 457254 280344 457260 280356
rect 440568 280316 457260 280344
rect 440568 280304 440574 280316
rect 457254 280304 457260 280316
rect 457312 280304 457318 280356
rect 468570 280304 468576 280356
rect 468628 280344 468634 280356
rect 484394 280344 484400 280356
rect 468628 280316 484400 280344
rect 468628 280304 468634 280316
rect 484394 280304 484400 280316
rect 484452 280304 484458 280356
rect 36722 280236 36728 280288
rect 36780 280276 36786 280288
rect 62114 280276 62120 280288
rect 36780 280248 62120 280276
rect 36780 280236 36786 280248
rect 62114 280236 62120 280248
rect 62172 280236 62178 280288
rect 64138 280236 64144 280288
rect 64196 280276 64202 280288
rect 89070 280276 89076 280288
rect 64196 280248 89076 280276
rect 64196 280236 64202 280248
rect 89070 280236 89076 280248
rect 89128 280236 89134 280288
rect 90450 280236 90456 280288
rect 90508 280276 90514 280288
rect 115934 280276 115940 280288
rect 90508 280248 115940 280276
rect 90508 280236 90514 280248
rect 115934 280236 115940 280248
rect 115992 280236 115998 280288
rect 116578 280236 116584 280288
rect 116636 280276 116642 280288
rect 142982 280276 142988 280288
rect 116636 280248 142988 280276
rect 116636 280236 116642 280248
rect 142982 280236 142988 280248
rect 143040 280236 143046 280288
rect 144270 280236 144276 280288
rect 144328 280276 144334 280288
rect 170030 280276 170036 280288
rect 144328 280248 170036 280276
rect 144328 280236 144334 280248
rect 170030 280236 170036 280248
rect 170088 280236 170094 280288
rect 178402 280236 178408 280288
rect 178460 280276 178466 280288
rect 200758 280276 200764 280288
rect 178460 280248 200764 280276
rect 178460 280236 178466 280248
rect 200758 280236 200764 280248
rect 200816 280236 200822 280288
rect 251450 280236 251456 280288
rect 251508 280276 251514 280288
rect 268286 280276 268292 280288
rect 251508 280248 268292 280276
rect 251508 280236 251514 280248
rect 268286 280236 268292 280248
rect 268344 280236 268350 280288
rect 279510 280236 279516 280288
rect 279568 280276 279574 280288
rect 295794 280276 295800 280288
rect 279568 280248 295800 280276
rect 279568 280236 279574 280248
rect 295794 280236 295800 280248
rect 295852 280236 295858 280288
rect 305546 280236 305552 280288
rect 305604 280276 305610 280288
rect 322382 280276 322388 280288
rect 305604 280248 322388 280276
rect 305604 280236 305610 280248
rect 322382 280236 322388 280248
rect 322440 280236 322446 280288
rect 335998 280236 336004 280288
rect 336056 280276 336062 280288
rect 349798 280276 349804 280288
rect 336056 280248 349804 280276
rect 336056 280236 336062 280248
rect 349798 280236 349804 280248
rect 349856 280236 349862 280288
rect 359642 280236 359648 280288
rect 359700 280276 359706 280288
rect 376294 280276 376300 280288
rect 359700 280248 376300 280276
rect 359700 280236 359706 280248
rect 376294 280236 376300 280248
rect 376352 280236 376358 280288
rect 386506 280236 386512 280288
rect 386564 280276 386570 280288
rect 403342 280276 403348 280288
rect 386564 280248 403348 280276
rect 386564 280236 386570 280248
rect 403342 280236 403348 280248
rect 403400 280236 403406 280288
rect 421282 280236 421288 280288
rect 421340 280276 421346 280288
rect 446398 280276 446404 280288
rect 421340 280248 446404 280276
rect 421340 280236 421346 280248
rect 446398 280236 446404 280248
rect 446456 280236 446462 280288
rect 494514 280236 494520 280288
rect 494572 280276 494578 280288
rect 511350 280276 511356 280288
rect 494572 280248 511356 280276
rect 494572 280236 494578 280248
rect 511350 280236 511356 280248
rect 511408 280236 511414 280288
rect 522298 280236 522304 280288
rect 522356 280276 522362 280288
rect 538398 280276 538404 280288
rect 522356 280248 538404 280276
rect 522356 280236 522362 280248
rect 538398 280236 538404 280248
rect 538456 280236 538462 280288
rect 43346 280168 43352 280220
rect 43404 280208 43410 280220
rect 62758 280208 62764 280220
rect 43404 280180 62764 280208
rect 43404 280168 43410 280180
rect 62758 280168 62764 280180
rect 62816 280168 62822 280220
rect 144178 280168 144184 280220
rect 144236 280208 144242 280220
rect 160278 280208 160284 280220
rect 144236 280180 160284 280208
rect 144236 280168 144242 280180
rect 160278 280168 160284 280180
rect 160336 280168 160342 280220
rect 171778 280168 171784 280220
rect 171836 280208 171842 280220
rect 197446 280208 197452 280220
rect 171836 280180 197452 280208
rect 171836 280168 171842 280180
rect 197446 280168 197452 280180
rect 197504 280168 197510 280220
rect 199378 280168 199384 280220
rect 199436 280208 199442 280220
rect 223942 280208 223948 280220
rect 199436 280180 223948 280208
rect 199436 280168 199442 280180
rect 223942 280168 223948 280180
rect 224000 280168 224006 280220
rect 225598 280168 225604 280220
rect 225656 280208 225662 280220
rect 251174 280208 251180 280220
rect 225656 280180 251180 280208
rect 225656 280168 225662 280180
rect 251174 280168 251180 280180
rect 251232 280168 251238 280220
rect 253198 280168 253204 280220
rect 253256 280208 253262 280220
rect 278038 280208 278044 280220
rect 253256 280180 278044 280208
rect 253256 280168 253262 280180
rect 278038 280168 278044 280180
rect 278096 280168 278102 280220
rect 279418 280168 279424 280220
rect 279476 280208 279482 280220
rect 305454 280208 305460 280220
rect 279476 280180 305460 280208
rect 279476 280168 279482 280180
rect 305454 280168 305460 280180
rect 305512 280168 305518 280220
rect 307018 280168 307024 280220
rect 307076 280208 307082 280220
rect 331950 280208 331956 280220
rect 307076 280180 331956 280208
rect 307076 280168 307082 280180
rect 331950 280168 331956 280180
rect 332008 280168 332014 280220
rect 333238 280168 333244 280220
rect 333296 280208 333302 280220
rect 359458 280208 359464 280220
rect 333296 280180 359464 280208
rect 333296 280168 333302 280180
rect 359458 280168 359464 280180
rect 359516 280168 359522 280220
rect 359734 280168 359740 280220
rect 359792 280208 359798 280220
rect 386046 280208 386052 280220
rect 359792 280180 386052 280208
rect 359792 280168 359798 280180
rect 386046 280168 386052 280180
rect 386104 280168 386110 280220
rect 387058 280168 387064 280220
rect 387116 280208 387122 280220
rect 412910 280208 412916 280220
rect 387116 280180 412916 280208
rect 387116 280168 387122 280180
rect 412910 280168 412916 280180
rect 412968 280168 412974 280220
rect 414658 280168 414664 280220
rect 414716 280208 414722 280220
rect 440234 280208 440240 280220
rect 414716 280180 440240 280208
rect 414716 280168 414722 280180
rect 440234 280168 440240 280180
rect 440292 280168 440298 280220
rect 442258 280168 442264 280220
rect 442316 280208 442322 280220
rect 467006 280208 467012 280220
rect 442316 280180 467012 280208
rect 442316 280168 442322 280180
rect 467006 280168 467012 280180
rect 467064 280168 467070 280220
rect 468478 280168 468484 280220
rect 468536 280208 468542 280220
rect 494054 280208 494060 280220
rect 468536 280180 494060 280208
rect 468536 280168 468542 280180
rect 494054 280168 494060 280180
rect 494112 280168 494118 280220
rect 496078 280168 496084 280220
rect 496136 280208 496142 280220
rect 520918 280208 520924 280220
rect 496136 280180 520924 280208
rect 496136 280168 496142 280180
rect 520918 280168 520924 280180
rect 520976 280168 520982 280220
rect 522390 280168 522396 280220
rect 522448 280208 522454 280220
rect 548058 280208 548064 280220
rect 522448 280180 548064 280208
rect 522448 280168 522454 280180
rect 548058 280168 548064 280180
rect 548116 280168 548122 280220
rect 37918 279420 37924 279472
rect 37976 279460 37982 279472
rect 526438 279460 526444 279472
rect 37976 279432 526444 279460
rect 37976 279420 37982 279432
rect 526438 279420 526444 279432
rect 526496 279420 526502 279472
rect 285766 278264 285772 278316
rect 285824 278304 285830 278316
rect 286134 278304 286140 278316
rect 285824 278276 286140 278304
rect 285824 278264 285830 278276
rect 286134 278264 286140 278276
rect 286192 278264 286198 278316
rect 339586 278264 339592 278316
rect 339644 278304 339650 278316
rect 340138 278304 340144 278316
rect 339644 278276 340144 278304
rect 339644 278264 339650 278276
rect 340138 278264 340144 278276
rect 340196 278264 340202 278316
rect 68922 277516 68928 277568
rect 68980 277556 68986 277568
rect 118694 277556 118700 277568
rect 68980 277528 118700 277556
rect 68980 277516 68986 277528
rect 118694 277516 118700 277528
rect 118752 277516 118758 277568
rect 311802 277516 311808 277568
rect 311860 277556 311866 277568
rect 361574 277556 361580 277568
rect 311860 277528 361580 277556
rect 311860 277516 311866 277528
rect 361574 277516 361580 277528
rect 361632 277516 361638 277568
rect 35618 277448 35624 277500
rect 35676 277488 35682 277500
rect 36630 277488 36636 277500
rect 35676 277460 36636 277488
rect 35676 277448 35682 277460
rect 36630 277448 36636 277460
rect 36688 277448 36694 277500
rect 41322 277448 41328 277500
rect 41380 277488 41386 277500
rect 91094 277488 91100 277500
rect 41380 277460 91100 277488
rect 41380 277448 41386 277460
rect 91094 277448 91100 277460
rect 91152 277448 91158 277500
rect 122742 277448 122748 277500
rect 122800 277488 122806 277500
rect 172514 277488 172520 277500
rect 122800 277460 172520 277488
rect 122800 277448 122806 277460
rect 172514 277448 172520 277460
rect 172572 277448 172578 277500
rect 176562 277448 176568 277500
rect 176620 277488 176626 277500
rect 226334 277488 226340 277500
rect 176620 277460 226340 277488
rect 176620 277448 176626 277460
rect 226334 277448 226340 277460
rect 226392 277448 226398 277500
rect 230382 277448 230388 277500
rect 230440 277488 230446 277500
rect 280154 277488 280160 277500
rect 230440 277460 280160 277488
rect 230440 277448 230446 277460
rect 280154 277448 280160 277460
rect 280212 277448 280218 277500
rect 284202 277448 284208 277500
rect 284260 277488 284266 277500
rect 335354 277488 335360 277500
rect 284260 277460 335360 277488
rect 284260 277448 284266 277460
rect 335354 277448 335360 277460
rect 335412 277448 335418 277500
rect 365622 277448 365628 277500
rect 365680 277488 365686 277500
rect 415394 277488 415400 277500
rect 365680 277460 415400 277488
rect 365680 277448 365686 277460
rect 415394 277448 415400 277460
rect 415452 277448 415458 277500
rect 419442 277448 419448 277500
rect 419500 277488 419506 277500
rect 469214 277488 469220 277500
rect 419500 277460 469220 277488
rect 419500 277448 419506 277460
rect 469214 277448 469220 277460
rect 469272 277448 469278 277500
rect 473262 277448 473268 277500
rect 473320 277488 473326 277500
rect 523034 277488 523040 277500
rect 473320 277460 523040 277488
rect 473320 277448 473326 277460
rect 523034 277448 523040 277460
rect 523092 277448 523098 277500
rect 13722 277380 13728 277432
rect 13780 277420 13786 277432
rect 64874 277420 64880 277432
rect 13780 277392 64880 277420
rect 13780 277380 13786 277392
rect 64874 277380 64880 277392
rect 64932 277380 64938 277432
rect 95142 277380 95148 277432
rect 95200 277420 95206 277432
rect 146294 277420 146300 277432
rect 95200 277392 146300 277420
rect 95200 277380 95206 277392
rect 146294 277380 146300 277392
rect 146352 277380 146358 277432
rect 148962 277380 148968 277432
rect 149020 277420 149026 277432
rect 200114 277420 200120 277432
rect 149020 277392 200120 277420
rect 149020 277380 149026 277392
rect 200114 277380 200120 277392
rect 200172 277380 200178 277432
rect 202782 277380 202788 277432
rect 202840 277420 202846 277432
rect 253934 277420 253940 277432
rect 202840 277392 253940 277420
rect 202840 277380 202846 277392
rect 253934 277380 253940 277392
rect 253992 277380 253998 277432
rect 256602 277380 256608 277432
rect 256660 277420 256666 277432
rect 307754 277420 307760 277432
rect 256660 277392 307760 277420
rect 256660 277380 256666 277392
rect 307754 277380 307760 277392
rect 307812 277380 307818 277432
rect 338022 277380 338028 277432
rect 338080 277420 338086 277432
rect 389174 277420 389180 277432
rect 338080 277392 389180 277420
rect 338080 277380 338086 277392
rect 389174 277380 389180 277392
rect 389232 277380 389238 277432
rect 391842 277380 391848 277432
rect 391900 277420 391906 277432
rect 442994 277420 443000 277432
rect 391900 277392 443000 277420
rect 391900 277380 391906 277392
rect 442994 277380 443000 277392
rect 443052 277380 443058 277432
rect 445662 277380 445668 277432
rect 445720 277420 445726 277432
rect 496814 277420 496820 277432
rect 445720 277392 496820 277420
rect 445720 277380 445726 277392
rect 496814 277380 496820 277392
rect 496872 277380 496878 277432
rect 500862 277380 500868 277432
rect 500920 277420 500926 277432
rect 550634 277420 550640 277432
rect 500920 277392 550640 277420
rect 500920 277380 500926 277392
rect 550634 277380 550640 277392
rect 550692 277380 550698 277432
rect 170214 259632 170220 259684
rect 170272 259672 170278 259684
rect 170490 259672 170496 259684
rect 170272 259644 170496 259672
rect 170272 259632 170278 259644
rect 170490 259632 170496 259644
rect 170548 259632 170554 259684
rect 446398 259428 446404 259480
rect 446456 259468 446462 259480
rect 447686 259468 447692 259480
rect 446456 259440 447692 259468
rect 446456 259428 446462 259440
rect 447686 259428 447692 259440
rect 447744 259428 447750 259480
rect 35618 259360 35624 259412
rect 35676 259400 35682 259412
rect 36814 259400 36820 259412
rect 35676 259372 36820 259400
rect 35676 259360 35682 259372
rect 36814 259360 36820 259372
rect 36872 259360 36878 259412
rect 278682 259360 278688 259412
rect 278740 259400 278746 259412
rect 279510 259400 279516 259412
rect 278740 259372 279516 259400
rect 278740 259360 278746 259372
rect 279510 259360 279516 259372
rect 279568 259360 279574 259412
rect 332594 259360 332600 259412
rect 332652 259400 332658 259412
rect 335998 259400 336004 259412
rect 332652 259372 336004 259400
rect 332652 259360 332658 259372
rect 335998 259360 336004 259372
rect 336056 259360 336062 259412
rect 467650 259360 467656 259412
rect 467708 259400 467714 259412
rect 468570 259400 468576 259412
rect 467708 259372 468576 259400
rect 467708 259360 467714 259372
rect 468570 259360 468576 259372
rect 468628 259360 468634 259412
rect 26050 256640 26056 256692
rect 26108 256680 26114 256692
rect 36722 256680 36728 256692
rect 26108 256652 36728 256680
rect 26108 256640 26114 256652
rect 36722 256640 36728 256652
rect 36780 256640 36786 256692
rect 62758 256640 62764 256692
rect 62816 256680 62822 256692
rect 69750 256680 69756 256692
rect 62816 256652 69756 256680
rect 62816 256640 62822 256652
rect 69750 256640 69756 256652
rect 69808 256640 69814 256692
rect 96614 256640 96620 256692
rect 96672 256680 96678 256692
rect 96672 256652 103514 256680
rect 96672 256640 96678 256652
rect 15194 256572 15200 256624
rect 15252 256612 15258 256624
rect 42794 256612 42800 256624
rect 15252 256584 42800 256612
rect 15252 256572 15258 256584
rect 42794 256572 42800 256584
rect 42852 256572 42858 256624
rect 53098 256572 53104 256624
rect 53156 256612 53162 256624
rect 64138 256612 64144 256624
rect 53156 256584 64144 256612
rect 53156 256572 53162 256584
rect 64138 256572 64144 256584
rect 64196 256572 64202 256624
rect 69106 256572 69112 256624
rect 69164 256612 69170 256624
rect 96706 256612 96712 256624
rect 69164 256584 96712 256612
rect 69164 256572 69170 256584
rect 96706 256572 96712 256584
rect 96764 256572 96770 256624
rect 103486 256612 103514 256652
rect 200758 256640 200764 256692
rect 200816 256680 200822 256692
rect 204622 256680 204628 256692
rect 200816 256652 204628 256680
rect 200816 256640 200822 256652
rect 204622 256640 204628 256652
rect 204680 256640 204686 256692
rect 251818 256640 251824 256692
rect 251876 256680 251882 256692
rect 258718 256680 258724 256692
rect 251876 256652 258724 256680
rect 251876 256640 251882 256652
rect 258718 256640 258724 256652
rect 258776 256640 258782 256692
rect 494698 256640 494704 256692
rect 494756 256680 494762 256692
rect 501598 256680 501604 256692
rect 494756 256652 501604 256680
rect 494756 256640 494762 256652
rect 501598 256640 501604 256652
rect 501656 256640 501662 256692
rect 123662 256612 123668 256624
rect 103486 256584 123668 256612
rect 123662 256572 123668 256584
rect 123720 256572 123726 256624
rect 149698 256572 149704 256624
rect 149756 256612 149762 256624
rect 547966 256612 547972 256624
rect 149756 256584 547972 256612
rect 149756 256572 149762 256584
rect 547966 256572 547972 256584
rect 548024 256572 548030 256624
rect 79962 256504 79968 256556
rect 80020 256544 80026 256556
rect 90450 256544 90456 256556
rect 80020 256516 90456 256544
rect 80020 256504 80026 256516
rect 90450 256504 90456 256516
rect 90508 256504 90514 256556
rect 106550 256504 106556 256556
rect 106608 256544 106614 256556
rect 116578 256544 116584 256556
rect 106608 256516 116584 256544
rect 106608 256504 106614 256516
rect 116578 256504 116584 256516
rect 116636 256504 116642 256556
rect 133782 256504 133788 256556
rect 133840 256544 133846 256556
rect 144270 256544 144276 256556
rect 133840 256516 144276 256544
rect 133840 256504 133846 256516
rect 144270 256504 144276 256516
rect 144328 256504 144334 256556
rect 150526 256504 150532 256556
rect 150584 256544 150590 256556
rect 178126 256544 178132 256556
rect 150584 256516 178132 256544
rect 150584 256504 150590 256516
rect 178126 256504 178132 256516
rect 178184 256504 178190 256556
rect 187970 256504 187976 256556
rect 188028 256544 188034 256556
rect 199378 256544 199384 256556
rect 188028 256516 199384 256544
rect 188028 256504 188034 256516
rect 199378 256504 199384 256516
rect 199436 256504 199442 256556
rect 204346 256504 204352 256556
rect 204404 256544 204410 256556
rect 231946 256544 231952 256556
rect 204404 256516 231952 256544
rect 204404 256504 204410 256516
rect 231946 256504 231952 256516
rect 232004 256504 232010 256556
rect 242066 256504 242072 256556
rect 242124 256544 242130 256556
rect 253198 256544 253204 256556
rect 242124 256516 253204 256544
rect 242124 256504 242130 256516
rect 253198 256504 253204 256516
rect 253256 256504 253262 256556
rect 258166 256504 258172 256556
rect 258224 256544 258230 256556
rect 258224 256516 281764 256544
rect 258224 256504 258230 256516
rect 122926 256436 122932 256488
rect 122984 256476 122990 256488
rect 150710 256476 150716 256488
rect 122984 256448 150716 256476
rect 122984 256436 122990 256448
rect 150710 256436 150716 256448
rect 150768 256436 150774 256488
rect 160554 256436 160560 256488
rect 160612 256476 160618 256488
rect 171778 256476 171784 256488
rect 160612 256448 171784 256476
rect 160612 256436 160618 256448
rect 171778 256436 171784 256448
rect 171836 256436 171842 256488
rect 215018 256436 215024 256488
rect 215076 256476 215082 256488
rect 225598 256476 225604 256488
rect 215076 256448 225604 256476
rect 215076 256436 215082 256448
rect 225598 256436 225604 256448
rect 225656 256436 225662 256488
rect 268930 256436 268936 256488
rect 268988 256476 268994 256488
rect 279418 256476 279424 256488
rect 268988 256448 279424 256476
rect 268988 256436 268994 256448
rect 279418 256436 279424 256448
rect 279476 256436 279482 256488
rect 281736 256476 281764 256516
rect 285766 256504 285772 256556
rect 285824 256544 285830 256556
rect 312630 256544 312636 256556
rect 285824 256516 312636 256544
rect 285824 256504 285830 256516
rect 312630 256504 312636 256516
rect 312688 256504 312694 256556
rect 340138 256544 340144 256556
rect 316006 256516 340144 256544
rect 286134 256476 286140 256488
rect 281736 256448 286140 256476
rect 286134 256436 286140 256448
rect 286192 256436 286198 256488
rect 295978 256436 295984 256488
rect 296036 256476 296042 256488
rect 307018 256476 307024 256488
rect 296036 256448 307024 256476
rect 296036 256436 296042 256448
rect 307018 256436 307024 256448
rect 307076 256436 307082 256488
rect 311986 256436 311992 256488
rect 312044 256476 312050 256488
rect 316006 256476 316034 256516
rect 340138 256504 340144 256516
rect 340196 256504 340202 256556
rect 344986 256516 364334 256544
rect 312044 256448 316034 256476
rect 312044 256436 312050 256448
rect 322842 256436 322848 256488
rect 322900 256476 322906 256488
rect 333238 256476 333244 256488
rect 322900 256448 333244 256476
rect 322900 256436 322906 256448
rect 333238 256436 333244 256448
rect 333296 256436 333302 256488
rect 339586 256436 339592 256488
rect 339644 256476 339650 256488
rect 344986 256476 345014 256516
rect 339644 256448 345014 256476
rect 339644 256436 339650 256448
rect 350074 256436 350080 256488
rect 350132 256476 350138 256488
rect 359550 256476 359556 256488
rect 350132 256448 359556 256476
rect 350132 256436 350138 256448
rect 359550 256436 359556 256448
rect 359608 256436 359614 256488
rect 364306 256476 364334 256516
rect 365806 256504 365812 256556
rect 365864 256544 365870 256556
rect 393590 256544 393596 256556
rect 365864 256516 393596 256544
rect 365864 256504 365870 256516
rect 393590 256504 393596 256516
rect 393648 256504 393654 256556
rect 420914 256544 420920 256556
rect 402946 256516 420920 256544
rect 366726 256476 366732 256488
rect 364306 256448 366732 256476
rect 366726 256436 366732 256448
rect 366784 256436 366790 256488
rect 376570 256436 376576 256488
rect 376628 256476 376634 256488
rect 387058 256476 387064 256488
rect 376628 256448 387064 256476
rect 376628 256436 376634 256448
rect 387058 256436 387064 256448
rect 387116 256436 387122 256488
rect 393406 256436 393412 256488
rect 393464 256476 393470 256488
rect 402946 256476 402974 256516
rect 420914 256504 420920 256516
rect 420972 256504 420978 256556
rect 431034 256504 431040 256556
rect 431092 256544 431098 256556
rect 442258 256544 442264 256556
rect 431092 256516 442264 256544
rect 431092 256504 431098 256516
rect 442258 256504 442264 256516
rect 442316 256504 442322 256556
rect 447226 256504 447232 256556
rect 447284 256544 447290 256556
rect 474734 256544 474740 256556
rect 447284 256516 474740 256544
rect 447284 256504 447290 256516
rect 474734 256504 474740 256516
rect 474792 256504 474798 256556
rect 484946 256504 484952 256556
rect 485004 256544 485010 256556
rect 496078 256544 496084 256556
rect 485004 256516 496084 256544
rect 485004 256504 485010 256516
rect 496078 256504 496084 256516
rect 496136 256504 496142 256556
rect 501046 256504 501052 256556
rect 501104 256544 501110 256556
rect 528646 256544 528652 256556
rect 501104 256516 528652 256544
rect 501104 256504 501110 256516
rect 528646 256504 528652 256516
rect 528704 256504 528710 256556
rect 393464 256448 402974 256476
rect 393464 256436 393470 256448
rect 403986 256436 403992 256488
rect 404044 256476 404050 256488
rect 414658 256476 414664 256488
rect 404044 256448 414664 256476
rect 404044 256436 404050 256448
rect 414658 256436 414664 256448
rect 414716 256436 414722 256488
rect 458082 256436 458088 256488
rect 458140 256476 458146 256488
rect 468478 256476 468484 256488
rect 458140 256448 468484 256476
rect 458140 256436 458146 256448
rect 468478 256436 468484 256448
rect 468536 256436 468542 256488
rect 511810 256436 511816 256488
rect 511868 256476 511874 256488
rect 522390 256476 522396 256488
rect 511868 256448 522396 256476
rect 511868 256436 511874 256448
rect 522390 256436 522396 256448
rect 522448 256436 522454 256488
rect 36538 256368 36544 256420
rect 36596 256408 36602 256420
rect 538398 256408 538404 256420
rect 36596 256380 538404 256408
rect 36596 256368 36602 256380
rect 538398 256368 538404 256380
rect 538456 256368 538462 256420
rect 16298 254532 16304 254584
rect 16356 254572 16362 254584
rect 529014 254572 529020 254584
rect 16356 254544 529020 254572
rect 16356 254532 16362 254544
rect 529014 254532 529020 254544
rect 529072 254532 529078 254584
rect 25682 254192 25688 254244
rect 25740 254232 25746 254244
rect 148318 254232 148324 254244
rect 25740 254204 148324 254232
rect 25740 254192 25746 254204
rect 148318 254192 148324 254204
rect 148376 254192 148382 254244
rect 36814 254124 36820 254176
rect 36872 254164 36878 254176
rect 52638 254164 52644 254176
rect 36872 254136 52644 254164
rect 36872 254124 36878 254136
rect 52638 254124 52644 254136
rect 52696 254124 52702 254176
rect 232038 254124 232044 254176
rect 232096 254164 232102 254176
rect 251818 254164 251824 254176
rect 232096 254136 251824 254164
rect 232096 254124 232102 254136
rect 251818 254124 251824 254136
rect 251876 254124 251882 254176
rect 475010 254124 475016 254176
rect 475068 254164 475074 254176
rect 494698 254164 494704 254176
rect 475068 254136 494704 254164
rect 475068 254124 475074 254136
rect 494698 254124 494704 254136
rect 494756 254124 494762 254176
rect 62482 254056 62488 254108
rect 62540 254096 62546 254108
rect 79686 254096 79692 254108
rect 62540 254068 79692 254096
rect 62540 254056 62546 254068
rect 79686 254056 79692 254068
rect 79744 254056 79750 254108
rect 90358 254056 90364 254108
rect 90416 254096 90422 254108
rect 106642 254096 106648 254108
rect 90416 254068 106648 254096
rect 90416 254056 90422 254068
rect 106642 254056 106648 254068
rect 106700 254056 106706 254108
rect 116486 254056 116492 254108
rect 116544 254096 116550 254108
rect 133690 254096 133696 254108
rect 116544 254068 133696 254096
rect 116544 254056 116550 254068
rect 133690 254056 133696 254068
rect 133748 254056 133754 254108
rect 170490 254056 170496 254108
rect 170548 254096 170554 254108
rect 187694 254096 187700 254108
rect 170548 254068 187700 254096
rect 170548 254056 170554 254068
rect 187694 254056 187700 254068
rect 187752 254056 187758 254108
rect 197446 254056 197452 254108
rect 197504 254096 197510 254108
rect 214650 254096 214656 254108
rect 197504 254068 214656 254096
rect 197504 254056 197510 254068
rect 214650 254056 214656 254068
rect 214708 254056 214714 254108
rect 224494 254056 224500 254108
rect 224552 254096 224558 254108
rect 241698 254096 241704 254108
rect 224552 254068 241704 254096
rect 224552 254056 224558 254068
rect 241698 254056 241704 254068
rect 241756 254056 241762 254108
rect 413462 254056 413468 254108
rect 413520 254096 413526 254108
rect 430666 254096 430672 254108
rect 413520 254068 430672 254096
rect 413520 254056 413526 254068
rect 430666 254056 430672 254068
rect 430724 254056 430730 254108
rect 440510 254056 440516 254108
rect 440568 254096 440574 254108
rect 457622 254096 457628 254108
rect 440568 254068 457628 254096
rect 440568 254056 440574 254068
rect 457622 254056 457628 254068
rect 457680 254056 457686 254108
rect 468570 254056 468576 254108
rect 468628 254096 468634 254108
rect 484670 254096 484676 254108
rect 468628 254068 484676 254096
rect 468628 254056 468634 254068
rect 484670 254056 484676 254068
rect 484728 254056 484734 254108
rect 36722 253988 36728 254040
rect 36780 254028 36786 254040
rect 62298 254028 62304 254040
rect 36780 254000 62304 254028
rect 36780 253988 36786 254000
rect 62298 253988 62304 254000
rect 62356 253988 62362 254040
rect 64138 253988 64144 254040
rect 64196 254028 64202 254040
rect 89346 254028 89352 254040
rect 64196 254000 89352 254028
rect 64196 253988 64202 254000
rect 89346 253988 89352 254000
rect 89404 253988 89410 254040
rect 90450 253988 90456 254040
rect 90508 254028 90514 254040
rect 116302 254028 116308 254040
rect 90508 254000 116308 254028
rect 90508 253988 90514 254000
rect 116302 253988 116308 254000
rect 116360 253988 116366 254040
rect 116578 253988 116584 254040
rect 116636 254028 116642 254040
rect 143350 254028 143356 254040
rect 116636 254000 143356 254028
rect 116636 253988 116642 254000
rect 143350 253988 143356 254000
rect 143408 253988 143414 254040
rect 144270 253988 144276 254040
rect 144328 254028 144334 254040
rect 170306 254028 170312 254040
rect 144328 254000 170312 254028
rect 144328 253988 144334 254000
rect 170306 253988 170312 254000
rect 170364 253988 170370 254040
rect 178034 253988 178040 254040
rect 178092 254028 178098 254040
rect 200758 254028 200764 254040
rect 178092 254000 200764 254028
rect 178092 253988 178098 254000
rect 200758 253988 200764 254000
rect 200816 253988 200822 254040
rect 251450 253988 251456 254040
rect 251508 254028 251514 254040
rect 268654 254028 268660 254040
rect 251508 254000 268660 254028
rect 251508 253988 251514 254000
rect 268654 253988 268660 254000
rect 268712 253988 268718 254040
rect 279418 253988 279424 254040
rect 279476 254028 279482 254040
rect 295702 254028 295708 254040
rect 279476 254000 295708 254028
rect 279476 253988 279482 254000
rect 295702 253988 295708 254000
rect 295760 253988 295766 254040
rect 305454 253988 305460 254040
rect 305512 254028 305518 254040
rect 322658 254028 322664 254040
rect 305512 254000 322664 254028
rect 305512 253988 305518 254000
rect 322658 253988 322664 254000
rect 322716 253988 322722 254040
rect 334618 253988 334624 254040
rect 334676 254028 334682 254040
rect 349706 254028 349712 254040
rect 334676 254000 349712 254028
rect 334676 253988 334682 254000
rect 349706 253988 349712 254000
rect 349764 253988 349770 254040
rect 359458 253988 359464 254040
rect 359516 254028 359522 254040
rect 376662 254028 376668 254040
rect 359516 254000 376668 254028
rect 359516 253988 359522 254000
rect 376662 253988 376668 254000
rect 376720 253988 376726 254040
rect 386506 253988 386512 254040
rect 386564 254028 386570 254040
rect 403618 254028 403624 254040
rect 386564 254000 403624 254028
rect 386564 253988 386570 254000
rect 403618 253988 403624 254000
rect 403676 253988 403682 254040
rect 421006 253988 421012 254040
rect 421064 254028 421070 254040
rect 443638 254028 443644 254040
rect 421064 254000 443644 254028
rect 421064 253988 421070 254000
rect 443638 253988 443644 254000
rect 443696 253988 443702 254040
rect 494514 253988 494520 254040
rect 494572 254028 494578 254040
rect 511626 254028 511632 254040
rect 494572 254000 511632 254028
rect 494572 253988 494578 254000
rect 511626 253988 511632 254000
rect 511684 253988 511690 254040
rect 522390 253988 522396 254040
rect 522448 254028 522454 254040
rect 538674 254028 538680 254040
rect 522448 254000 538680 254028
rect 522448 253988 522454 254000
rect 538674 253988 538680 254000
rect 538732 253988 538738 254040
rect 43070 253920 43076 253972
rect 43128 253960 43134 253972
rect 62758 253960 62764 253972
rect 43128 253932 62764 253960
rect 43128 253920 43134 253932
rect 62758 253920 62764 253932
rect 62816 253920 62822 253972
rect 144178 253920 144184 253972
rect 144236 253960 144242 253972
rect 160646 253960 160652 253972
rect 144236 253932 160652 253960
rect 144236 253920 144242 253932
rect 160646 253920 160652 253932
rect 160704 253920 160710 253972
rect 171778 253920 171784 253972
rect 171836 253960 171842 253972
rect 197354 253960 197360 253972
rect 171836 253932 197360 253960
rect 171836 253920 171842 253932
rect 197354 253920 197360 253932
rect 197412 253920 197418 253972
rect 199378 253920 199384 253972
rect 199436 253960 199442 253972
rect 224310 253960 224316 253972
rect 199436 253932 224316 253960
rect 199436 253920 199442 253932
rect 224310 253920 224316 253932
rect 224368 253920 224374 253972
rect 225598 253920 225604 253972
rect 225656 253960 225662 253972
rect 251358 253960 251364 253972
rect 225656 253932 251364 253960
rect 225656 253920 225662 253932
rect 251358 253920 251364 253932
rect 251416 253920 251422 253972
rect 253198 253920 253204 253972
rect 253256 253960 253262 253972
rect 278314 253960 278320 253972
rect 253256 253932 278320 253960
rect 253256 253920 253262 253932
rect 278314 253920 278320 253932
rect 278372 253920 278378 253972
rect 279510 253920 279516 253972
rect 279568 253960 279574 253972
rect 305362 253960 305368 253972
rect 279568 253932 305368 253960
rect 279568 253920 279574 253932
rect 305362 253920 305368 253932
rect 305420 253920 305426 253972
rect 307018 253920 307024 253972
rect 307076 253960 307082 253972
rect 332318 253960 332324 253972
rect 307076 253932 332324 253960
rect 307076 253920 307082 253932
rect 332318 253920 332324 253932
rect 332376 253920 332382 253972
rect 333238 253920 333244 253972
rect 333296 253960 333302 253972
rect 359366 253960 359372 253972
rect 333296 253932 359372 253960
rect 333296 253920 333302 253932
rect 359366 253920 359372 253932
rect 359424 253920 359430 253972
rect 359550 253920 359556 253972
rect 359608 253960 359614 253972
rect 386322 253960 386328 253972
rect 359608 253932 386328 253960
rect 359608 253920 359614 253932
rect 386322 253920 386328 253932
rect 386380 253920 386386 253972
rect 387058 253920 387064 253972
rect 387116 253960 387122 253972
rect 413278 253960 413284 253972
rect 387116 253932 413284 253960
rect 387116 253920 387122 253932
rect 413278 253920 413284 253932
rect 413336 253920 413342 253972
rect 414658 253920 414664 253972
rect 414716 253960 414722 253972
rect 440326 253960 440332 253972
rect 414716 253932 440332 253960
rect 414716 253920 414722 253932
rect 440326 253920 440332 253932
rect 440384 253920 440390 253972
rect 442258 253920 442264 253972
rect 442316 253960 442322 253972
rect 467282 253960 467288 253972
rect 442316 253932 467288 253960
rect 442316 253920 442322 253932
rect 467282 253920 467288 253932
rect 467340 253920 467346 253972
rect 468478 253920 468484 253972
rect 468536 253960 468542 253972
rect 494330 253960 494336 253972
rect 468536 253932 494336 253960
rect 468536 253920 468542 253932
rect 494330 253920 494336 253932
rect 494388 253920 494394 253972
rect 496078 253920 496084 253972
rect 496136 253960 496142 253972
rect 521286 253960 521292 253972
rect 496136 253932 521292 253960
rect 496136 253920 496142 253932
rect 521286 253920 521292 253932
rect 521344 253920 521350 253972
rect 522298 253920 522304 253972
rect 522356 253960 522362 253972
rect 548334 253960 548340 253972
rect 522356 253932 548340 253960
rect 522356 253920 522362 253932
rect 548334 253920 548340 253932
rect 548392 253920 548398 253972
rect 37918 251812 37924 251864
rect 37976 251852 37982 251864
rect 526438 251852 526444 251864
rect 37976 251824 526444 251852
rect 37976 251812 37982 251824
rect 526438 251812 526444 251824
rect 526496 251812 526502 251864
rect 68922 251268 68928 251320
rect 68980 251308 68986 251320
rect 118694 251308 118700 251320
rect 68980 251280 118700 251308
rect 68980 251268 68986 251280
rect 118694 251268 118700 251280
rect 118752 251268 118758 251320
rect 122742 251268 122748 251320
rect 122800 251308 122806 251320
rect 172514 251308 172520 251320
rect 122800 251280 172520 251308
rect 122800 251268 122806 251280
rect 172514 251268 172520 251280
rect 172572 251268 172578 251320
rect 230382 251268 230388 251320
rect 230440 251308 230446 251320
rect 280154 251308 280160 251320
rect 230440 251280 280160 251308
rect 230440 251268 230446 251280
rect 280154 251268 280160 251280
rect 280212 251268 280218 251320
rect 311802 251268 311808 251320
rect 311860 251308 311866 251320
rect 361574 251308 361580 251320
rect 311860 251280 361580 251308
rect 311860 251268 311866 251280
rect 361574 251268 361580 251280
rect 361632 251268 361638 251320
rect 500862 251268 500868 251320
rect 500920 251308 500926 251320
rect 550634 251308 550640 251320
rect 500920 251280 550640 251308
rect 500920 251268 500926 251280
rect 550634 251268 550640 251280
rect 550692 251268 550698 251320
rect 41322 251200 41328 251252
rect 41380 251240 41386 251252
rect 91094 251240 91100 251252
rect 41380 251212 91100 251240
rect 41380 251200 41386 251212
rect 91094 251200 91100 251212
rect 91152 251200 91158 251252
rect 148962 251200 148968 251252
rect 149020 251240 149026 251252
rect 200114 251240 200120 251252
rect 149020 251212 200120 251240
rect 149020 251200 149026 251212
rect 200114 251200 200120 251212
rect 200172 251200 200178 251252
rect 202782 251200 202788 251252
rect 202840 251240 202846 251252
rect 253934 251240 253940 251252
rect 202840 251212 253940 251240
rect 202840 251200 202846 251212
rect 253934 251200 253940 251212
rect 253992 251200 253998 251252
rect 284202 251200 284208 251252
rect 284260 251240 284266 251252
rect 335354 251240 335360 251252
rect 284260 251212 335360 251240
rect 284260 251200 284266 251212
rect 335354 251200 335360 251212
rect 335412 251200 335418 251252
rect 365622 251200 365628 251252
rect 365680 251240 365686 251252
rect 415394 251240 415400 251252
rect 365680 251212 415400 251240
rect 365680 251200 365686 251212
rect 415394 251200 415400 251212
rect 415452 251200 415458 251252
rect 419442 251200 419448 251252
rect 419500 251240 419506 251252
rect 469214 251240 469220 251252
rect 419500 251212 469220 251240
rect 419500 251200 419506 251212
rect 469214 251200 469220 251212
rect 469272 251200 469278 251252
rect 473262 251200 473268 251252
rect 473320 251240 473326 251252
rect 523034 251240 523040 251252
rect 473320 251212 523040 251240
rect 473320 251200 473326 251212
rect 523034 251200 523040 251212
rect 523092 251200 523098 251252
rect 521746 235356 521752 235408
rect 521804 235396 521810 235408
rect 522390 235396 522396 235408
rect 521804 235368 522396 235396
rect 521804 235356 521810 235368
rect 522390 235356 522396 235368
rect 522448 235356 522454 235408
rect 13722 233180 13728 233232
rect 13780 233220 13786 233232
rect 64874 233220 64880 233232
rect 13780 233192 64880 233220
rect 13780 233180 13786 233192
rect 64874 233180 64880 233192
rect 64932 233180 64938 233232
rect 95142 233180 95148 233232
rect 95200 233220 95206 233232
rect 146294 233220 146300 233232
rect 95200 233192 146300 233220
rect 95200 233180 95206 233192
rect 146294 233180 146300 233192
rect 146352 233180 146358 233232
rect 176562 233180 176568 233232
rect 176620 233220 176626 233232
rect 226334 233220 226340 233232
rect 176620 233192 226340 233220
rect 176620 233180 176626 233192
rect 226334 233180 226340 233192
rect 226392 233180 226398 233232
rect 256602 233180 256608 233232
rect 256660 233220 256666 233232
rect 307754 233220 307760 233232
rect 256660 233192 307760 233220
rect 256660 233180 256666 233192
rect 307754 233180 307760 233192
rect 307812 233180 307818 233232
rect 332502 233180 332508 233232
rect 332560 233220 332566 233232
rect 334618 233220 334624 233232
rect 332560 233192 334624 233220
rect 332560 233180 332566 233192
rect 334618 233180 334624 233192
rect 334676 233180 334682 233232
rect 338022 233180 338028 233232
rect 338080 233220 338086 233232
rect 389174 233220 389180 233232
rect 338080 233192 389180 233220
rect 338080 233180 338086 233192
rect 389174 233180 389180 233192
rect 389232 233180 389238 233232
rect 391842 233180 391848 233232
rect 391900 233220 391906 233232
rect 442994 233220 443000 233232
rect 391900 233192 443000 233220
rect 391900 233180 391906 233192
rect 442994 233180 443000 233192
rect 443052 233180 443058 233232
rect 445662 233180 445668 233232
rect 445720 233220 445726 233232
rect 496814 233220 496820 233232
rect 445720 233192 496820 233220
rect 445720 233180 445726 233192
rect 496814 233180 496820 233192
rect 496872 233180 496878 233232
rect 467650 233112 467656 233164
rect 467708 233152 467714 233164
rect 468570 233152 468576 233164
rect 467708 233124 468576 233152
rect 467708 233112 467714 233124
rect 468570 233112 468576 233124
rect 468628 233112 468634 233164
rect 35618 232704 35624 232756
rect 35676 232744 35682 232756
rect 36814 232744 36820 232756
rect 35676 232716 36820 232744
rect 35676 232704 35682 232716
rect 36814 232704 36820 232716
rect 36872 232704 36878 232756
rect 257982 231820 257988 231872
rect 258040 231860 258046 231872
rect 258718 231860 258724 231872
rect 258040 231832 258724 231860
rect 258040 231820 258046 231832
rect 258718 231820 258724 231832
rect 258776 231820 258782 231872
rect 494698 231820 494704 231872
rect 494756 231860 494762 231872
rect 501598 231860 501604 231872
rect 494756 231832 501604 231860
rect 494756 231820 494762 231832
rect 501598 231820 501604 231832
rect 501656 231820 501662 231872
rect 26050 230392 26056 230444
rect 26108 230432 26114 230444
rect 36722 230432 36728 230444
rect 26108 230404 36728 230432
rect 26108 230392 26114 230404
rect 36722 230392 36728 230404
rect 36780 230392 36786 230444
rect 62758 230392 62764 230444
rect 62816 230432 62822 230444
rect 69750 230432 69756 230444
rect 62816 230404 69756 230432
rect 62816 230392 62822 230404
rect 69750 230392 69756 230404
rect 69808 230392 69814 230444
rect 96706 230392 96712 230444
rect 96764 230432 96770 230444
rect 96764 230404 103514 230432
rect 96764 230392 96770 230404
rect 15194 230324 15200 230376
rect 15252 230364 15258 230376
rect 42794 230364 42800 230376
rect 15252 230336 42800 230364
rect 15252 230324 15258 230336
rect 42794 230324 42800 230336
rect 42852 230324 42858 230376
rect 53098 230324 53104 230376
rect 53156 230364 53162 230376
rect 64138 230364 64144 230376
rect 53156 230336 64144 230364
rect 53156 230324 53162 230336
rect 64138 230324 64144 230336
rect 64196 230324 64202 230376
rect 69106 230324 69112 230376
rect 69164 230364 69170 230376
rect 96798 230364 96804 230376
rect 69164 230336 96804 230364
rect 69164 230324 69170 230336
rect 96798 230324 96804 230336
rect 96856 230324 96862 230376
rect 103486 230364 103514 230404
rect 146938 230392 146944 230444
rect 146996 230432 147002 230444
rect 146996 230404 151814 230432
rect 146996 230392 147002 230404
rect 123662 230364 123668 230376
rect 103486 230336 123668 230364
rect 123662 230324 123668 230336
rect 123720 230324 123726 230376
rect 133782 230324 133788 230376
rect 133840 230364 133846 230376
rect 144270 230364 144276 230376
rect 133840 230336 144276 230364
rect 133840 230324 133846 230336
rect 144270 230324 144276 230336
rect 144328 230324 144334 230376
rect 150710 230364 150716 230376
rect 146588 230336 150716 230364
rect 79962 230256 79968 230308
rect 80020 230296 80026 230308
rect 90450 230296 90456 230308
rect 80020 230268 90456 230296
rect 80020 230256 80026 230268
rect 90450 230256 90456 230268
rect 90508 230256 90514 230308
rect 106550 230256 106556 230308
rect 106608 230296 106614 230308
rect 116578 230296 116584 230308
rect 106608 230268 116584 230296
rect 106608 230256 106614 230268
rect 116578 230256 116584 230268
rect 116636 230256 116642 230308
rect 122926 230256 122932 230308
rect 122984 230296 122990 230308
rect 146588 230296 146616 230336
rect 150710 230324 150716 230336
rect 150768 230324 150774 230376
rect 151786 230364 151814 230404
rect 200758 230392 200764 230444
rect 200816 230432 200822 230444
rect 204622 230432 204628 230444
rect 200816 230404 204628 230432
rect 200816 230392 200822 230404
rect 204622 230392 204628 230404
rect 204680 230392 204686 230444
rect 251818 230392 251824 230444
rect 251876 230432 251882 230444
rect 257982 230432 257988 230444
rect 251876 230404 257988 230432
rect 251876 230392 251882 230404
rect 257982 230392 257988 230404
rect 258040 230392 258046 230444
rect 443638 230392 443644 230444
rect 443696 230432 443702 230444
rect 447686 230432 447692 230444
rect 443696 230404 447692 230432
rect 443696 230392 443702 230404
rect 447686 230392 447692 230404
rect 447744 230392 447750 230444
rect 547966 230364 547972 230376
rect 151786 230336 547972 230364
rect 547966 230324 547972 230336
rect 548024 230324 548030 230376
rect 122984 230268 146616 230296
rect 122984 230256 122990 230268
rect 150526 230256 150532 230308
rect 150584 230296 150590 230308
rect 178126 230296 178132 230308
rect 150584 230268 178132 230296
rect 150584 230256 150590 230268
rect 178126 230256 178132 230268
rect 178184 230256 178190 230308
rect 187970 230256 187976 230308
rect 188028 230296 188034 230308
rect 199378 230296 199384 230308
rect 188028 230268 199384 230296
rect 188028 230256 188034 230268
rect 199378 230256 199384 230268
rect 199436 230256 199442 230308
rect 204346 230256 204352 230308
rect 204404 230296 204410 230308
rect 231854 230296 231860 230308
rect 204404 230268 231860 230296
rect 204404 230256 204410 230268
rect 231854 230256 231860 230268
rect 231912 230256 231918 230308
rect 242066 230256 242072 230308
rect 242124 230296 242130 230308
rect 253198 230296 253204 230308
rect 242124 230268 253204 230296
rect 242124 230256 242130 230268
rect 253198 230256 253204 230268
rect 253256 230256 253262 230308
rect 258166 230256 258172 230308
rect 258224 230296 258230 230308
rect 286134 230296 286140 230308
rect 258224 230268 286140 230296
rect 258224 230256 258230 230268
rect 286134 230256 286140 230268
rect 286192 230256 286198 230308
rect 312630 230296 312636 230308
rect 287026 230268 312636 230296
rect 160554 230188 160560 230240
rect 160612 230228 160618 230240
rect 171778 230228 171784 230240
rect 160612 230200 171784 230228
rect 160612 230188 160618 230200
rect 171778 230188 171784 230200
rect 171836 230188 171842 230240
rect 215018 230188 215024 230240
rect 215076 230228 215082 230240
rect 225598 230228 225604 230240
rect 215076 230200 225604 230228
rect 215076 230188 215082 230200
rect 225598 230188 225604 230200
rect 225656 230188 225662 230240
rect 268930 230188 268936 230240
rect 268988 230228 268994 230240
rect 279510 230228 279516 230240
rect 268988 230200 279516 230228
rect 268988 230188 268994 230200
rect 279510 230188 279516 230200
rect 279568 230188 279574 230240
rect 285766 230188 285772 230240
rect 285824 230228 285830 230240
rect 287026 230228 287054 230268
rect 312630 230256 312636 230268
rect 312688 230256 312694 230308
rect 340138 230296 340144 230308
rect 316006 230268 340144 230296
rect 285824 230200 287054 230228
rect 285824 230188 285830 230200
rect 295978 230188 295984 230240
rect 296036 230228 296042 230240
rect 307018 230228 307024 230240
rect 296036 230200 307024 230228
rect 296036 230188 296042 230200
rect 307018 230188 307024 230200
rect 307076 230188 307082 230240
rect 311986 230188 311992 230240
rect 312044 230228 312050 230240
rect 316006 230228 316034 230268
rect 340138 230256 340144 230268
rect 340196 230256 340202 230308
rect 366726 230296 366732 230308
rect 344986 230268 366732 230296
rect 312044 230200 316034 230228
rect 312044 230188 312050 230200
rect 322842 230188 322848 230240
rect 322900 230228 322906 230240
rect 333238 230228 333244 230240
rect 322900 230200 333244 230228
rect 322900 230188 322906 230200
rect 333238 230188 333244 230200
rect 333296 230188 333302 230240
rect 339586 230188 339592 230240
rect 339644 230228 339650 230240
rect 344986 230228 345014 230268
rect 366726 230256 366732 230268
rect 366784 230256 366790 230308
rect 393590 230296 393596 230308
rect 373966 230268 393596 230296
rect 339644 230200 345014 230228
rect 339644 230188 339650 230200
rect 350074 230188 350080 230240
rect 350132 230228 350138 230240
rect 359550 230228 359556 230240
rect 350132 230200 359556 230228
rect 350132 230188 350138 230200
rect 359550 230188 359556 230200
rect 359608 230188 359614 230240
rect 365806 230188 365812 230240
rect 365864 230228 365870 230240
rect 373966 230228 373994 230268
rect 393590 230256 393596 230268
rect 393648 230256 393654 230308
rect 420914 230296 420920 230308
rect 402946 230268 420920 230296
rect 365864 230200 373994 230228
rect 365864 230188 365870 230200
rect 376570 230188 376576 230240
rect 376628 230228 376634 230240
rect 387058 230228 387064 230240
rect 376628 230200 387064 230228
rect 376628 230188 376634 230200
rect 387058 230188 387064 230200
rect 387116 230188 387122 230240
rect 393406 230188 393412 230240
rect 393464 230228 393470 230240
rect 402946 230228 402974 230268
rect 420914 230256 420920 230268
rect 420972 230256 420978 230308
rect 431034 230256 431040 230308
rect 431092 230296 431098 230308
rect 442258 230296 442264 230308
rect 431092 230268 442264 230296
rect 431092 230256 431098 230268
rect 442258 230256 442264 230268
rect 442316 230256 442322 230308
rect 447226 230256 447232 230308
rect 447284 230296 447290 230308
rect 474734 230296 474740 230308
rect 447284 230268 474740 230296
rect 447284 230256 447290 230268
rect 474734 230256 474740 230268
rect 474792 230256 474798 230308
rect 484946 230256 484952 230308
rect 485004 230296 485010 230308
rect 496078 230296 496084 230308
rect 485004 230268 496084 230296
rect 485004 230256 485010 230268
rect 496078 230256 496084 230268
rect 496136 230256 496142 230308
rect 501046 230256 501052 230308
rect 501104 230296 501110 230308
rect 528646 230296 528652 230308
rect 501104 230268 528652 230296
rect 501104 230256 501110 230268
rect 528646 230256 528652 230268
rect 528704 230256 528710 230308
rect 393464 230200 402974 230228
rect 393464 230188 393470 230200
rect 403986 230188 403992 230240
rect 404044 230228 404050 230240
rect 414658 230228 414664 230240
rect 404044 230200 414664 230228
rect 404044 230188 404050 230200
rect 414658 230188 414664 230200
rect 414716 230188 414722 230240
rect 458082 230188 458088 230240
rect 458140 230228 458146 230240
rect 468478 230228 468484 230240
rect 458140 230200 468484 230228
rect 458140 230188 458146 230200
rect 468478 230188 468484 230200
rect 468536 230188 468542 230240
rect 511902 230188 511908 230240
rect 511960 230228 511966 230240
rect 522298 230228 522304 230240
rect 511960 230200 522304 230228
rect 511960 230188 511966 230200
rect 522298 230188 522304 230200
rect 522356 230188 522362 230240
rect 36630 230120 36636 230172
rect 36688 230160 36694 230172
rect 538398 230160 538404 230172
rect 36688 230132 538404 230160
rect 36688 230120 36694 230132
rect 538398 230120 538404 230132
rect 538456 230120 538462 230172
rect 15286 226992 15292 227044
rect 15344 227032 15350 227044
rect 528738 227032 528744 227044
rect 15344 227004 528744 227032
rect 15344 226992 15350 227004
rect 528738 226992 528744 227004
rect 528796 226992 528802 227044
rect 25958 226584 25964 226636
rect 26016 226624 26022 226636
rect 146938 226624 146944 226636
rect 26016 226596 146944 226624
rect 26016 226584 26022 226596
rect 146938 226584 146944 226596
rect 146996 226584 147002 226636
rect 36814 226516 36820 226568
rect 36872 226556 36878 226568
rect 52454 226556 52460 226568
rect 36872 226528 52460 226556
rect 36872 226516 36878 226528
rect 52454 226516 52460 226528
rect 52512 226516 52518 226568
rect 62482 226516 62488 226568
rect 62540 226556 62546 226568
rect 79318 226556 79324 226568
rect 62540 226528 79324 226556
rect 62540 226516 62546 226528
rect 79318 226516 79324 226528
rect 79376 226516 79382 226568
rect 259362 226516 259368 226568
rect 259420 226556 259426 226568
rect 279602 226556 279608 226568
rect 259420 226528 279608 226556
rect 259420 226516 259426 226528
rect 279602 226516 279608 226528
rect 279660 226516 279666 226568
rect 448330 226516 448336 226568
rect 448388 226556 448394 226568
rect 468662 226556 468668 226568
rect 448388 226528 468668 226556
rect 448388 226516 448394 226528
rect 468662 226516 468668 226528
rect 468720 226516 468726 226568
rect 43346 226448 43352 226500
rect 43404 226488 43410 226500
rect 62758 226488 62764 226500
rect 43404 226460 62764 226488
rect 43404 226448 43410 226460
rect 62758 226448 62764 226460
rect 62816 226448 62822 226500
rect 90358 226448 90364 226500
rect 90416 226488 90422 226500
rect 106366 226488 106372 226500
rect 90416 226460 106372 226488
rect 90416 226448 90422 226460
rect 106366 226448 106372 226460
rect 106424 226448 106430 226500
rect 116486 226448 116492 226500
rect 116544 226488 116550 226500
rect 133414 226488 133420 226500
rect 116544 226460 133420 226488
rect 116544 226448 116550 226460
rect 133414 226448 133420 226460
rect 133472 226448 133478 226500
rect 170490 226448 170496 226500
rect 170548 226488 170554 226500
rect 187786 226488 187792 226500
rect 170548 226460 187792 226488
rect 170548 226448 170554 226460
rect 187786 226448 187792 226460
rect 187844 226448 187850 226500
rect 197538 226448 197544 226500
rect 197596 226488 197602 226500
rect 214374 226488 214380 226500
rect 197596 226460 214380 226488
rect 197596 226448 197602 226460
rect 214374 226448 214380 226460
rect 214432 226448 214438 226500
rect 224494 226448 224500 226500
rect 224552 226488 224558 226500
rect 241514 226488 241520 226500
rect 224552 226460 241520 226488
rect 224552 226448 224558 226460
rect 241514 226448 241520 226460
rect 241572 226448 241578 226500
rect 251450 226448 251456 226500
rect 251508 226488 251514 226500
rect 268286 226488 268292 226500
rect 251508 226460 268292 226488
rect 251508 226448 251514 226460
rect 268286 226448 268292 226460
rect 268344 226448 268350 226500
rect 413462 226448 413468 226500
rect 413520 226488 413526 226500
rect 430574 226488 430580 226500
rect 413520 226460 430580 226488
rect 413520 226448 413526 226460
rect 430574 226448 430580 226460
rect 430632 226448 430638 226500
rect 440510 226448 440516 226500
rect 440568 226488 440574 226500
rect 457254 226488 457260 226500
rect 440568 226460 457260 226488
rect 440568 226448 440574 226460
rect 457254 226448 457260 226460
rect 457312 226448 457318 226500
rect 36722 226380 36728 226432
rect 36780 226420 36786 226432
rect 62114 226420 62120 226432
rect 36780 226392 62120 226420
rect 36780 226380 36786 226392
rect 62114 226380 62120 226392
rect 62172 226380 62178 226432
rect 64138 226380 64144 226432
rect 64196 226420 64202 226432
rect 89070 226420 89076 226432
rect 64196 226392 89076 226420
rect 64196 226380 64202 226392
rect 89070 226380 89076 226392
rect 89128 226380 89134 226432
rect 90450 226380 90456 226432
rect 90508 226420 90514 226432
rect 115934 226420 115940 226432
rect 90508 226392 115940 226420
rect 90508 226380 90514 226392
rect 115934 226380 115940 226392
rect 115992 226380 115998 226432
rect 116578 226380 116584 226432
rect 116636 226420 116642 226432
rect 142982 226420 142988 226432
rect 116636 226392 142988 226420
rect 116636 226380 116642 226392
rect 142982 226380 142988 226392
rect 143040 226380 143046 226432
rect 144270 226380 144276 226432
rect 144328 226420 144334 226432
rect 170030 226420 170036 226432
rect 144328 226392 170036 226420
rect 144328 226380 144334 226392
rect 170030 226380 170036 226392
rect 170088 226380 170094 226432
rect 178402 226380 178408 226432
rect 178460 226420 178466 226432
rect 200758 226420 200764 226432
rect 178460 226392 200764 226420
rect 178460 226380 178466 226392
rect 200758 226380 200764 226392
rect 200816 226380 200822 226432
rect 232314 226380 232320 226432
rect 232372 226420 232378 226432
rect 251818 226420 251824 226432
rect 232372 226392 251824 226420
rect 232372 226380 232378 226392
rect 251818 226380 251824 226392
rect 251876 226380 251882 226432
rect 279418 226380 279424 226432
rect 279476 226420 279482 226432
rect 295794 226420 295800 226432
rect 279476 226392 295800 226420
rect 279476 226380 279482 226392
rect 295794 226380 295800 226392
rect 295852 226380 295858 226432
rect 305638 226380 305644 226432
rect 305696 226420 305702 226432
rect 322382 226420 322388 226432
rect 305696 226392 322388 226420
rect 305696 226380 305702 226392
rect 322382 226380 322388 226392
rect 322440 226380 322446 226432
rect 335998 226380 336004 226432
rect 336056 226420 336062 226432
rect 349798 226420 349804 226432
rect 336056 226392 349804 226420
rect 336056 226380 336062 226392
rect 349798 226380 349804 226392
rect 349856 226380 349862 226432
rect 359550 226380 359556 226432
rect 359608 226420 359614 226432
rect 376294 226420 376300 226432
rect 359608 226392 376300 226420
rect 359608 226380 359614 226392
rect 376294 226380 376300 226392
rect 376352 226380 376358 226432
rect 386506 226380 386512 226432
rect 386564 226420 386570 226432
rect 403342 226420 403348 226432
rect 386564 226392 403348 226420
rect 386564 226380 386570 226392
rect 403342 226380 403348 226392
rect 403400 226380 403406 226432
rect 421282 226380 421288 226432
rect 421340 226420 421346 226432
rect 445018 226420 445024 226432
rect 421340 226392 445024 226420
rect 421340 226380 421346 226392
rect 445018 226380 445024 226392
rect 445076 226380 445082 226432
rect 468570 226380 468576 226432
rect 468628 226420 468634 226432
rect 484394 226420 484400 226432
rect 468628 226392 484400 226420
rect 468628 226380 468634 226392
rect 484394 226380 484400 226392
rect 484452 226380 484458 226432
rect 494514 226380 494520 226432
rect 494572 226420 494578 226432
rect 511350 226420 511356 226432
rect 494572 226392 511356 226420
rect 494572 226380 494578 226392
rect 511350 226380 511356 226392
rect 511408 226380 511414 226432
rect 522390 226380 522396 226432
rect 522448 226420 522454 226432
rect 538398 226420 538404 226432
rect 522448 226392 538404 226420
rect 522448 226380 522454 226392
rect 538398 226380 538404 226392
rect 538456 226380 538462 226432
rect 70302 226312 70308 226364
rect 70360 226352 70366 226364
rect 90542 226352 90548 226364
rect 70360 226324 90548 226352
rect 70360 226312 70366 226324
rect 90542 226312 90548 226324
rect 90600 226312 90606 226364
rect 144178 226312 144184 226364
rect 144236 226352 144242 226364
rect 160278 226352 160284 226364
rect 144236 226324 160284 226352
rect 144236 226312 144242 226324
rect 160278 226312 160284 226324
rect 160336 226312 160342 226364
rect 171778 226312 171784 226364
rect 171836 226352 171842 226364
rect 197446 226352 197452 226364
rect 171836 226324 197452 226352
rect 171836 226312 171842 226324
rect 197446 226312 197452 226324
rect 197504 226312 197510 226364
rect 199378 226312 199384 226364
rect 199436 226352 199442 226364
rect 223942 226352 223948 226364
rect 199436 226324 223948 226352
rect 199436 226312 199442 226324
rect 223942 226312 223948 226324
rect 224000 226312 224006 226364
rect 225598 226312 225604 226364
rect 225656 226352 225662 226364
rect 251174 226352 251180 226364
rect 225656 226324 251180 226352
rect 225656 226312 225662 226324
rect 251174 226312 251180 226324
rect 251232 226312 251238 226364
rect 253198 226312 253204 226364
rect 253256 226352 253262 226364
rect 278038 226352 278044 226364
rect 253256 226324 278044 226352
rect 253256 226312 253262 226324
rect 278038 226312 278044 226324
rect 278096 226312 278102 226364
rect 279510 226312 279516 226364
rect 279568 226352 279574 226364
rect 305546 226352 305552 226364
rect 279568 226324 305552 226352
rect 279568 226312 279574 226324
rect 305546 226312 305552 226324
rect 305604 226312 305610 226364
rect 307018 226312 307024 226364
rect 307076 226352 307082 226364
rect 331950 226352 331956 226364
rect 307076 226324 331956 226352
rect 307076 226312 307082 226324
rect 331950 226312 331956 226324
rect 332008 226312 332014 226364
rect 333238 226312 333244 226364
rect 333296 226352 333302 226364
rect 359458 226352 359464 226364
rect 333296 226324 359464 226352
rect 333296 226312 333302 226324
rect 359458 226312 359464 226324
rect 359516 226312 359522 226364
rect 359734 226312 359740 226364
rect 359792 226352 359798 226364
rect 386046 226352 386052 226364
rect 359792 226324 386052 226352
rect 359792 226312 359798 226324
rect 386046 226312 386052 226324
rect 386104 226312 386110 226364
rect 387058 226312 387064 226364
rect 387116 226352 387122 226364
rect 412910 226352 412916 226364
rect 387116 226324 412916 226352
rect 387116 226312 387122 226324
rect 412910 226312 412916 226324
rect 412968 226312 412974 226364
rect 414658 226312 414664 226364
rect 414716 226352 414722 226364
rect 440234 226352 440240 226364
rect 414716 226324 440240 226352
rect 414716 226312 414722 226324
rect 440234 226312 440240 226324
rect 440292 226312 440298 226364
rect 442258 226312 442264 226364
rect 442316 226352 442322 226364
rect 467006 226352 467012 226364
rect 442316 226324 467012 226352
rect 442316 226312 442322 226324
rect 467006 226312 467012 226324
rect 467064 226312 467070 226364
rect 468478 226312 468484 226364
rect 468536 226352 468542 226364
rect 494054 226352 494060 226364
rect 468536 226324 494060 226352
rect 468536 226312 468542 226324
rect 494054 226312 494060 226324
rect 494112 226312 494118 226364
rect 496078 226312 496084 226364
rect 496136 226352 496142 226364
rect 520918 226352 520924 226364
rect 496136 226324 520924 226352
rect 496136 226312 496142 226324
rect 520918 226312 520924 226324
rect 520976 226312 520982 226364
rect 522298 226312 522304 226364
rect 522356 226352 522362 226364
rect 548058 226352 548064 226364
rect 522356 226324 548064 226352
rect 522356 226312 522362 226324
rect 548058 226312 548064 226324
rect 548116 226312 548122 226364
rect 37918 225564 37924 225616
rect 37976 225604 37982 225616
rect 526438 225604 526444 225616
rect 37976 225576 526444 225604
rect 37976 225564 37982 225576
rect 526438 225564 526444 225576
rect 526496 225564 526502 225616
rect 285766 224272 285772 224324
rect 285824 224312 285830 224324
rect 286134 224312 286140 224324
rect 285824 224284 286140 224312
rect 285824 224272 285830 224284
rect 286134 224272 286140 224284
rect 286192 224272 286198 224324
rect 339586 224272 339592 224324
rect 339644 224312 339650 224324
rect 340138 224312 340144 224324
rect 339644 224284 340144 224312
rect 339644 224272 339650 224284
rect 340138 224272 340144 224284
rect 340196 224272 340202 224324
rect 35618 223592 35624 223644
rect 35676 223632 35682 223644
rect 36630 223632 36636 223644
rect 35676 223604 36636 223632
rect 35676 223592 35682 223604
rect 36630 223592 36636 223604
rect 36688 223592 36694 223644
rect 90542 206252 90548 206304
rect 90600 206292 90606 206304
rect 96798 206292 96804 206304
rect 90600 206264 96804 206292
rect 90600 206252 90606 206264
rect 96798 206252 96804 206264
rect 96856 206252 96862 206304
rect 468662 206252 468668 206304
rect 468720 206292 468726 206304
rect 474734 206292 474740 206304
rect 468720 206264 474740 206292
rect 468720 206252 468726 206264
rect 474734 206252 474740 206264
rect 474792 206252 474798 206304
rect 474826 205708 474832 205760
rect 474884 205708 474890 205760
rect 279602 205640 279608 205692
rect 279660 205680 279666 205692
rect 286134 205680 286140 205692
rect 279660 205652 286140 205680
rect 279660 205640 279666 205652
rect 286134 205640 286140 205652
rect 286192 205640 286198 205692
rect 445018 205640 445024 205692
rect 445076 205680 445082 205692
rect 447686 205680 447692 205692
rect 445076 205652 447692 205680
rect 445076 205640 445082 205652
rect 447686 205640 447692 205652
rect 447744 205640 447750 205692
rect 474844 205680 474872 205708
rect 475194 205680 475200 205692
rect 474844 205652 475200 205680
rect 475194 205640 475200 205652
rect 475252 205640 475258 205692
rect 521746 205640 521752 205692
rect 521804 205680 521810 205692
rect 522390 205680 522396 205692
rect 521804 205652 522396 205680
rect 521804 205640 521810 205652
rect 522390 205640 522396 205652
rect 522448 205640 522454 205692
rect 13722 205572 13728 205624
rect 13780 205612 13786 205624
rect 64874 205612 64880 205624
rect 13780 205584 64880 205612
rect 13780 205572 13786 205584
rect 64874 205572 64880 205584
rect 64932 205572 64938 205624
rect 95142 205572 95148 205624
rect 95200 205612 95206 205624
rect 146294 205612 146300 205624
rect 95200 205584 146300 205612
rect 95200 205572 95206 205584
rect 146294 205572 146300 205584
rect 146352 205572 146358 205624
rect 148962 205572 148968 205624
rect 149020 205612 149026 205624
rect 200114 205612 200120 205624
rect 149020 205584 200120 205612
rect 149020 205572 149026 205584
rect 200114 205572 200120 205584
rect 200172 205572 200178 205624
rect 202782 205572 202788 205624
rect 202840 205612 202846 205624
rect 253934 205612 253940 205624
rect 202840 205584 253940 205612
rect 202840 205572 202846 205584
rect 253934 205572 253940 205584
rect 253992 205572 253998 205624
rect 256602 205572 256608 205624
rect 256660 205612 256666 205624
rect 307754 205612 307760 205624
rect 256660 205584 307760 205612
rect 256660 205572 256666 205584
rect 307754 205572 307760 205584
rect 307812 205572 307818 205624
rect 338022 205572 338028 205624
rect 338080 205612 338086 205624
rect 389174 205612 389180 205624
rect 338080 205584 389180 205612
rect 338080 205572 338086 205584
rect 389174 205572 389180 205584
rect 389232 205572 389238 205624
rect 391842 205572 391848 205624
rect 391900 205612 391906 205624
rect 442994 205612 443000 205624
rect 391900 205584 443000 205612
rect 391900 205572 391906 205584
rect 442994 205572 443000 205584
rect 443052 205572 443058 205624
rect 445662 205572 445668 205624
rect 445720 205612 445726 205624
rect 496814 205612 496820 205624
rect 445720 205584 496820 205612
rect 445720 205572 445726 205584
rect 496814 205572 496820 205584
rect 496872 205572 496878 205624
rect 500862 205572 500868 205624
rect 500920 205612 500926 205624
rect 550634 205612 550640 205624
rect 500920 205584 550640 205612
rect 500920 205572 500926 205584
rect 550634 205572 550640 205584
rect 550692 205572 550698 205624
rect 35618 205504 35624 205556
rect 35676 205544 35682 205556
rect 36814 205544 36820 205556
rect 35676 205516 36820 205544
rect 35676 205504 35682 205516
rect 36814 205504 36820 205516
rect 36872 205504 36878 205556
rect 41322 205504 41328 205556
rect 41380 205544 41386 205556
rect 91094 205544 91100 205556
rect 41380 205516 91100 205544
rect 41380 205504 41386 205516
rect 91094 205504 91100 205516
rect 91152 205504 91158 205556
rect 122742 205504 122748 205556
rect 122800 205544 122806 205556
rect 172514 205544 172520 205556
rect 122800 205516 172520 205544
rect 122800 205504 122806 205516
rect 172514 205504 172520 205516
rect 172572 205504 172578 205556
rect 176562 205504 176568 205556
rect 176620 205544 176626 205556
rect 226334 205544 226340 205556
rect 176620 205516 226340 205544
rect 176620 205504 176626 205516
rect 226334 205504 226340 205516
rect 226392 205504 226398 205556
rect 230382 205504 230388 205556
rect 230440 205544 230446 205556
rect 280154 205544 280160 205556
rect 230440 205516 280160 205544
rect 230440 205504 230446 205516
rect 280154 205504 280160 205516
rect 280212 205504 280218 205556
rect 284202 205504 284208 205556
rect 284260 205544 284266 205556
rect 335354 205544 335360 205556
rect 284260 205516 335360 205544
rect 284260 205504 284266 205516
rect 335354 205504 335360 205516
rect 335412 205504 335418 205556
rect 365622 205504 365628 205556
rect 365680 205544 365686 205556
rect 415394 205544 415400 205556
rect 365680 205516 415400 205544
rect 365680 205504 365686 205516
rect 415394 205504 415400 205516
rect 415452 205504 415458 205556
rect 419442 205504 419448 205556
rect 419500 205544 419506 205556
rect 469214 205544 469220 205556
rect 419500 205516 469220 205544
rect 419500 205504 419506 205516
rect 469214 205504 469220 205516
rect 469272 205504 469278 205556
rect 473262 205504 473268 205556
rect 473320 205544 473326 205556
rect 523034 205544 523040 205556
rect 473320 205516 523040 205544
rect 473320 205504 473326 205516
rect 523034 205504 523040 205516
rect 523092 205504 523098 205556
rect 68922 205436 68928 205488
rect 68980 205476 68986 205488
rect 118694 205476 118700 205488
rect 68980 205448 118700 205476
rect 68980 205436 68986 205448
rect 118694 205436 118700 205448
rect 118752 205436 118758 205488
rect 200758 205436 200764 205488
rect 200816 205476 200822 205488
rect 204622 205476 204628 205488
rect 200816 205448 204628 205476
rect 200816 205436 200822 205448
rect 204622 205436 204628 205448
rect 204680 205436 204686 205488
rect 311802 205436 311808 205488
rect 311860 205476 311866 205488
rect 361574 205476 361580 205488
rect 311860 205448 361580 205476
rect 311860 205436 311866 205448
rect 361574 205436 361580 205448
rect 361632 205436 361638 205488
rect 467650 205436 467656 205488
rect 467708 205476 467714 205488
rect 468570 205476 468576 205488
rect 467708 205448 468576 205476
rect 467708 205436 467714 205448
rect 468570 205436 468576 205448
rect 468628 205436 468634 205488
rect 53098 202784 53104 202836
rect 53156 202824 53162 202836
rect 64138 202824 64144 202836
rect 53156 202796 64144 202824
rect 53156 202784 53162 202796
rect 64138 202784 64144 202796
rect 64196 202784 64202 202836
rect 251818 202784 251824 202836
rect 251876 202824 251882 202836
rect 258994 202824 259000 202836
rect 251876 202796 259000 202824
rect 251876 202784 251882 202796
rect 258994 202784 259000 202796
rect 259052 202784 259058 202836
rect 332318 202784 332324 202836
rect 332376 202824 332382 202836
rect 335998 202824 336004 202836
rect 332376 202796 336004 202824
rect 332376 202784 332382 202796
rect 335998 202784 336004 202796
rect 336056 202784 336062 202836
rect 15194 202716 15200 202768
rect 15252 202756 15258 202768
rect 42978 202756 42984 202768
rect 15252 202728 42984 202756
rect 15252 202716 15258 202728
rect 42978 202716 42984 202728
rect 43036 202716 43042 202768
rect 62758 202716 62764 202768
rect 62816 202756 62822 202768
rect 70026 202756 70032 202768
rect 62816 202728 70032 202756
rect 62816 202716 62822 202728
rect 70026 202716 70032 202728
rect 70084 202716 70090 202768
rect 79686 202716 79692 202768
rect 79744 202756 79750 202768
rect 90450 202756 90456 202768
rect 79744 202728 90456 202756
rect 79744 202716 79750 202728
rect 90450 202716 90456 202728
rect 90508 202716 90514 202768
rect 96706 202716 96712 202768
rect 96764 202756 96770 202768
rect 124030 202756 124036 202768
rect 96764 202728 124036 202756
rect 96764 202716 96770 202728
rect 124030 202716 124036 202728
rect 124088 202716 124094 202768
rect 148318 202716 148324 202768
rect 148376 202756 148382 202768
rect 548334 202756 548340 202768
rect 148376 202728 548340 202756
rect 148376 202716 148382 202728
rect 548334 202716 548340 202728
rect 548392 202716 548398 202768
rect 25682 202648 25688 202700
rect 25740 202688 25746 202700
rect 36722 202688 36728 202700
rect 25740 202660 36728 202688
rect 25740 202648 25746 202660
rect 36722 202648 36728 202660
rect 36780 202648 36786 202700
rect 106642 202648 106648 202700
rect 106700 202688 106706 202700
rect 116578 202688 116584 202700
rect 106700 202660 116584 202688
rect 106700 202648 106706 202660
rect 116578 202648 116584 202660
rect 116636 202648 116642 202700
rect 133690 202648 133696 202700
rect 133748 202688 133754 202700
rect 144270 202688 144276 202700
rect 133748 202660 144276 202688
rect 133748 202648 133754 202660
rect 144270 202648 144276 202660
rect 144328 202648 144334 202700
rect 150526 202648 150532 202700
rect 150584 202688 150590 202700
rect 178034 202688 178040 202700
rect 150584 202660 178040 202688
rect 150584 202648 150590 202660
rect 178034 202648 178040 202660
rect 178092 202648 178098 202700
rect 187694 202648 187700 202700
rect 187752 202688 187758 202700
rect 199378 202688 199384 202700
rect 187752 202660 199384 202688
rect 187752 202648 187758 202660
rect 199378 202648 199384 202660
rect 199436 202648 199442 202700
rect 204346 202648 204352 202700
rect 204404 202688 204410 202700
rect 232038 202688 232044 202700
rect 204404 202660 232044 202688
rect 204404 202648 204410 202660
rect 232038 202648 232044 202660
rect 232096 202648 232102 202700
rect 241698 202648 241704 202700
rect 241756 202688 241762 202700
rect 253198 202688 253204 202700
rect 241756 202660 253204 202688
rect 241756 202648 241762 202660
rect 253198 202648 253204 202660
rect 253256 202648 253262 202700
rect 268654 202648 268660 202700
rect 268712 202688 268718 202700
rect 279510 202688 279516 202700
rect 268712 202660 279516 202688
rect 268712 202648 268718 202660
rect 279510 202648 279516 202660
rect 279568 202648 279574 202700
rect 285766 202648 285772 202700
rect 285824 202688 285830 202700
rect 312998 202688 313004 202700
rect 285824 202660 313004 202688
rect 285824 202648 285830 202660
rect 312998 202648 313004 202660
rect 313056 202648 313062 202700
rect 340046 202688 340052 202700
rect 316006 202660 340052 202688
rect 122926 202580 122932 202632
rect 122984 202620 122990 202632
rect 150986 202620 150992 202632
rect 122984 202592 150992 202620
rect 122984 202580 122990 202592
rect 150986 202580 150992 202592
rect 151044 202580 151050 202632
rect 160646 202580 160652 202632
rect 160704 202620 160710 202632
rect 171778 202620 171784 202632
rect 160704 202592 171784 202620
rect 160704 202580 160710 202592
rect 171778 202580 171784 202592
rect 171836 202580 171842 202632
rect 214650 202580 214656 202632
rect 214708 202620 214714 202632
rect 225598 202620 225604 202632
rect 214708 202592 225604 202620
rect 214708 202580 214714 202592
rect 225598 202580 225604 202592
rect 225656 202580 225662 202632
rect 295702 202580 295708 202632
rect 295760 202620 295766 202632
rect 307018 202620 307024 202632
rect 295760 202592 307024 202620
rect 295760 202580 295766 202592
rect 307018 202580 307024 202592
rect 307076 202580 307082 202632
rect 311986 202580 311992 202632
rect 312044 202620 312050 202632
rect 316006 202620 316034 202660
rect 340046 202648 340052 202660
rect 340104 202648 340110 202700
rect 367002 202688 367008 202700
rect 344986 202660 367008 202688
rect 312044 202592 316034 202620
rect 312044 202580 312050 202592
rect 322658 202580 322664 202632
rect 322716 202620 322722 202632
rect 333238 202620 333244 202632
rect 322716 202592 333244 202620
rect 322716 202580 322722 202592
rect 333238 202580 333244 202592
rect 333296 202580 333302 202632
rect 339586 202580 339592 202632
rect 339644 202620 339650 202632
rect 344986 202620 345014 202660
rect 367002 202648 367008 202660
rect 367060 202648 367066 202700
rect 393590 202688 393596 202700
rect 373966 202660 393596 202688
rect 339644 202592 345014 202620
rect 339644 202580 339650 202592
rect 349706 202580 349712 202632
rect 349764 202620 349770 202632
rect 359550 202620 359556 202632
rect 349764 202592 359556 202620
rect 349764 202580 349770 202592
rect 359550 202580 359556 202592
rect 359608 202580 359614 202632
rect 365806 202580 365812 202632
rect 365864 202620 365870 202632
rect 373966 202620 373994 202660
rect 393590 202648 393596 202660
rect 393648 202648 393654 202700
rect 421006 202688 421012 202700
rect 402946 202660 421012 202688
rect 365864 202592 373994 202620
rect 365864 202580 365870 202592
rect 376662 202580 376668 202632
rect 376720 202620 376726 202632
rect 387058 202620 387064 202632
rect 376720 202592 387064 202620
rect 376720 202580 376726 202592
rect 387058 202580 387064 202592
rect 387116 202580 387122 202632
rect 393406 202580 393412 202632
rect 393464 202620 393470 202632
rect 402946 202620 402974 202660
rect 421006 202648 421012 202660
rect 421064 202648 421070 202700
rect 430666 202648 430672 202700
rect 430724 202688 430730 202700
rect 442258 202688 442264 202700
rect 430724 202660 442264 202688
rect 430724 202648 430730 202660
rect 442258 202648 442264 202660
rect 442316 202648 442322 202700
rect 457714 202648 457720 202700
rect 457772 202688 457778 202700
rect 468478 202688 468484 202700
rect 457772 202660 468484 202688
rect 457772 202648 457778 202660
rect 468478 202648 468484 202660
rect 468536 202648 468542 202700
rect 475194 202648 475200 202700
rect 475252 202688 475258 202700
rect 501966 202688 501972 202700
rect 475252 202660 501972 202688
rect 475252 202648 475258 202660
rect 501966 202648 501972 202660
rect 502024 202648 502030 202700
rect 529014 202688 529020 202700
rect 509206 202660 529020 202688
rect 393464 202592 402974 202620
rect 393464 202580 393470 202592
rect 403710 202580 403716 202632
rect 403768 202620 403774 202632
rect 414658 202620 414664 202632
rect 403768 202592 414664 202620
rect 403768 202580 403774 202592
rect 414658 202580 414664 202592
rect 414716 202580 414722 202632
rect 484670 202580 484676 202632
rect 484728 202620 484734 202632
rect 496078 202620 496084 202632
rect 484728 202592 496084 202620
rect 484728 202580 484734 202592
rect 496078 202580 496084 202592
rect 496136 202580 496142 202632
rect 501046 202580 501052 202632
rect 501104 202620 501110 202632
rect 509206 202620 509234 202660
rect 529014 202648 529020 202660
rect 529072 202648 529078 202700
rect 501104 202592 509234 202620
rect 501104 202580 501110 202592
rect 511718 202580 511724 202632
rect 511776 202620 511782 202632
rect 522298 202620 522304 202632
rect 511776 202592 522304 202620
rect 511776 202580 511782 202592
rect 522298 202580 522304 202592
rect 522356 202580 522362 202632
rect 36538 202512 36544 202564
rect 36596 202552 36602 202564
rect 538674 202552 538680 202564
rect 36596 202524 538680 202552
rect 36596 202512 36602 202524
rect 538674 202512 538680 202524
rect 538732 202512 538738 202564
rect 16022 200744 16028 200796
rect 16080 200784 16086 200796
rect 529014 200784 529020 200796
rect 16080 200756 529020 200784
rect 16080 200744 16086 200756
rect 529014 200744 529020 200756
rect 529072 200744 529078 200796
rect 25682 200404 25688 200456
rect 25740 200444 25746 200456
rect 149698 200444 149704 200456
rect 25740 200416 149704 200444
rect 25740 200404 25746 200416
rect 149698 200404 149704 200416
rect 149756 200404 149762 200456
rect 36722 200336 36728 200388
rect 36780 200376 36786 200388
rect 52638 200376 52644 200388
rect 36780 200348 52644 200376
rect 36780 200336 36786 200348
rect 52638 200336 52644 200348
rect 52696 200336 52702 200388
rect 232038 200336 232044 200388
rect 232096 200376 232102 200388
rect 251818 200376 251824 200388
rect 232096 200348 251824 200376
rect 232096 200336 232102 200348
rect 251818 200336 251824 200348
rect 251876 200336 251882 200388
rect 43070 200268 43076 200320
rect 43128 200308 43134 200320
rect 62758 200308 62764 200320
rect 43128 200280 62764 200308
rect 43128 200268 43134 200280
rect 62758 200268 62764 200280
rect 62816 200268 62822 200320
rect 90358 200268 90364 200320
rect 90416 200308 90422 200320
rect 106642 200308 106648 200320
rect 90416 200280 106648 200308
rect 90416 200268 90422 200280
rect 106642 200268 106648 200280
rect 106700 200268 106706 200320
rect 116486 200268 116492 200320
rect 116544 200308 116550 200320
rect 133690 200308 133696 200320
rect 116544 200280 133696 200308
rect 116544 200268 116550 200280
rect 133690 200268 133696 200280
rect 133748 200268 133754 200320
rect 144178 200268 144184 200320
rect 144236 200308 144242 200320
rect 160646 200308 160652 200320
rect 144236 200280 160652 200308
rect 144236 200268 144242 200280
rect 160646 200268 160652 200280
rect 160704 200268 160710 200320
rect 170490 200268 170496 200320
rect 170548 200308 170554 200320
rect 187694 200308 187700 200320
rect 170548 200280 187700 200308
rect 170548 200268 170554 200280
rect 187694 200268 187700 200280
rect 187752 200268 187758 200320
rect 197446 200268 197452 200320
rect 197504 200308 197510 200320
rect 214650 200308 214656 200320
rect 197504 200280 214656 200308
rect 197504 200268 197510 200280
rect 214650 200268 214656 200280
rect 214708 200268 214714 200320
rect 224494 200268 224500 200320
rect 224552 200308 224558 200320
rect 241698 200308 241704 200320
rect 224552 200280 241704 200308
rect 224552 200268 224558 200280
rect 241698 200268 241704 200280
rect 241756 200268 241762 200320
rect 413462 200268 413468 200320
rect 413520 200308 413526 200320
rect 430666 200308 430672 200320
rect 413520 200280 430672 200308
rect 413520 200268 413526 200280
rect 430666 200268 430672 200280
rect 430724 200268 430730 200320
rect 440510 200268 440516 200320
rect 440568 200308 440574 200320
rect 457622 200308 457628 200320
rect 440568 200280 457628 200308
rect 440568 200268 440574 200280
rect 457622 200268 457628 200280
rect 457680 200268 457686 200320
rect 468570 200268 468576 200320
rect 468628 200308 468634 200320
rect 484670 200308 484676 200320
rect 468628 200280 484676 200308
rect 468628 200268 468634 200280
rect 484670 200268 484676 200280
rect 484728 200268 484734 200320
rect 494514 200268 494520 200320
rect 494572 200308 494578 200320
rect 511626 200308 511632 200320
rect 494572 200280 511632 200308
rect 494572 200268 494578 200280
rect 511626 200268 511632 200280
rect 511684 200268 511690 200320
rect 36814 200200 36820 200252
rect 36872 200240 36878 200252
rect 62298 200240 62304 200252
rect 36872 200212 62304 200240
rect 36872 200200 36878 200212
rect 62298 200200 62304 200212
rect 62356 200200 62362 200252
rect 64138 200200 64144 200252
rect 64196 200240 64202 200252
rect 89346 200240 89352 200252
rect 64196 200212 89352 200240
rect 64196 200200 64202 200212
rect 89346 200200 89352 200212
rect 89404 200200 89410 200252
rect 90450 200200 90456 200252
rect 90508 200240 90514 200252
rect 116302 200240 116308 200252
rect 90508 200212 116308 200240
rect 90508 200200 90514 200212
rect 116302 200200 116308 200212
rect 116360 200200 116366 200252
rect 116578 200200 116584 200252
rect 116636 200240 116642 200252
rect 143350 200240 143356 200252
rect 116636 200212 143356 200240
rect 116636 200200 116642 200212
rect 143350 200200 143356 200212
rect 143408 200200 143414 200252
rect 144270 200200 144276 200252
rect 144328 200240 144334 200252
rect 170306 200240 170312 200252
rect 144328 200212 170312 200240
rect 144328 200200 144334 200212
rect 170306 200200 170312 200212
rect 170364 200200 170370 200252
rect 178034 200200 178040 200252
rect 178092 200240 178098 200252
rect 200758 200240 200764 200252
rect 178092 200212 200764 200240
rect 178092 200200 178098 200212
rect 200758 200200 200764 200212
rect 200816 200200 200822 200252
rect 251450 200200 251456 200252
rect 251508 200240 251514 200252
rect 268654 200240 268660 200252
rect 251508 200212 268660 200240
rect 251508 200200 251514 200212
rect 268654 200200 268660 200212
rect 268712 200200 268718 200252
rect 279418 200200 279424 200252
rect 279476 200240 279482 200252
rect 295702 200240 295708 200252
rect 279476 200212 295708 200240
rect 279476 200200 279482 200212
rect 295702 200200 295708 200212
rect 295760 200200 295766 200252
rect 305454 200200 305460 200252
rect 305512 200240 305518 200252
rect 322658 200240 322664 200252
rect 305512 200212 322664 200240
rect 305512 200200 305518 200212
rect 322658 200200 322664 200212
rect 322716 200200 322722 200252
rect 335998 200200 336004 200252
rect 336056 200240 336062 200252
rect 349706 200240 349712 200252
rect 336056 200212 349712 200240
rect 336056 200200 336062 200212
rect 349706 200200 349712 200212
rect 349764 200200 349770 200252
rect 359458 200200 359464 200252
rect 359516 200240 359522 200252
rect 376662 200240 376668 200252
rect 359516 200212 376668 200240
rect 359516 200200 359522 200212
rect 376662 200200 376668 200212
rect 376720 200200 376726 200252
rect 386506 200200 386512 200252
rect 386564 200240 386570 200252
rect 403618 200240 403624 200252
rect 386564 200212 403624 200240
rect 386564 200200 386570 200212
rect 403618 200200 403624 200212
rect 403676 200200 403682 200252
rect 421006 200200 421012 200252
rect 421064 200240 421070 200252
rect 446398 200240 446404 200252
rect 421064 200212 446404 200240
rect 421064 200200 421070 200212
rect 446398 200200 446404 200212
rect 446456 200200 446462 200252
rect 475010 200200 475016 200252
rect 475068 200240 475074 200252
rect 494698 200240 494704 200252
rect 475068 200212 494704 200240
rect 475068 200200 475074 200212
rect 494698 200200 494704 200212
rect 494756 200200 494762 200252
rect 522390 200200 522396 200252
rect 522448 200240 522454 200252
rect 538674 200240 538680 200252
rect 522448 200212 538680 200240
rect 522448 200200 522454 200212
rect 538674 200200 538680 200212
rect 538732 200200 538738 200252
rect 62482 200132 62488 200184
rect 62540 200172 62546 200184
rect 79686 200172 79692 200184
rect 62540 200144 79692 200172
rect 62540 200132 62546 200144
rect 79686 200132 79692 200144
rect 79744 200132 79750 200184
rect 171778 200132 171784 200184
rect 171836 200172 171842 200184
rect 197354 200172 197360 200184
rect 171836 200144 197360 200172
rect 171836 200132 171842 200144
rect 197354 200132 197360 200144
rect 197412 200132 197418 200184
rect 199378 200132 199384 200184
rect 199436 200172 199442 200184
rect 224310 200172 224316 200184
rect 199436 200144 224316 200172
rect 199436 200132 199442 200144
rect 224310 200132 224316 200144
rect 224368 200132 224374 200184
rect 225598 200132 225604 200184
rect 225656 200172 225662 200184
rect 251358 200172 251364 200184
rect 225656 200144 251364 200172
rect 225656 200132 225662 200144
rect 251358 200132 251364 200144
rect 251416 200132 251422 200184
rect 253198 200132 253204 200184
rect 253256 200172 253262 200184
rect 278314 200172 278320 200184
rect 253256 200144 278320 200172
rect 253256 200132 253262 200144
rect 278314 200132 278320 200144
rect 278372 200132 278378 200184
rect 279510 200132 279516 200184
rect 279568 200172 279574 200184
rect 305362 200172 305368 200184
rect 279568 200144 305368 200172
rect 279568 200132 279574 200144
rect 305362 200132 305368 200144
rect 305420 200132 305426 200184
rect 307018 200132 307024 200184
rect 307076 200172 307082 200184
rect 332318 200172 332324 200184
rect 307076 200144 332324 200172
rect 307076 200132 307082 200144
rect 332318 200132 332324 200144
rect 332376 200132 332382 200184
rect 333238 200132 333244 200184
rect 333296 200172 333302 200184
rect 359366 200172 359372 200184
rect 333296 200144 359372 200172
rect 333296 200132 333302 200144
rect 359366 200132 359372 200144
rect 359424 200132 359430 200184
rect 359550 200132 359556 200184
rect 359608 200172 359614 200184
rect 386322 200172 386328 200184
rect 359608 200144 386328 200172
rect 359608 200132 359614 200144
rect 386322 200132 386328 200144
rect 386380 200132 386386 200184
rect 387058 200132 387064 200184
rect 387116 200172 387122 200184
rect 413278 200172 413284 200184
rect 387116 200144 413284 200172
rect 387116 200132 387122 200144
rect 413278 200132 413284 200144
rect 413336 200132 413342 200184
rect 414658 200132 414664 200184
rect 414716 200172 414722 200184
rect 440326 200172 440332 200184
rect 414716 200144 440332 200172
rect 414716 200132 414722 200144
rect 440326 200132 440332 200144
rect 440384 200132 440390 200184
rect 442258 200132 442264 200184
rect 442316 200172 442322 200184
rect 467282 200172 467288 200184
rect 442316 200144 467288 200172
rect 442316 200132 442322 200144
rect 467282 200132 467288 200144
rect 467340 200132 467346 200184
rect 468478 200132 468484 200184
rect 468536 200172 468542 200184
rect 494330 200172 494336 200184
rect 468536 200144 494336 200172
rect 468536 200132 468542 200144
rect 494330 200132 494336 200144
rect 494388 200132 494394 200184
rect 496078 200132 496084 200184
rect 496136 200172 496142 200184
rect 521286 200172 521292 200184
rect 496136 200144 521292 200172
rect 496136 200132 496142 200144
rect 521286 200132 521292 200144
rect 521344 200132 521350 200184
rect 522298 200132 522304 200184
rect 522356 200172 522362 200184
rect 548334 200172 548340 200184
rect 522356 200144 548340 200172
rect 522356 200132 522362 200144
rect 548334 200132 548340 200144
rect 548392 200132 548398 200184
rect 37918 197956 37924 198008
rect 37976 197996 37982 198008
rect 526438 197996 526444 198008
rect 37976 197968 526444 197996
rect 37976 197956 37982 197968
rect 526438 197956 526444 197968
rect 526496 197956 526502 198008
rect 445662 179392 445668 179444
rect 445720 179432 445726 179444
rect 445720 179404 454034 179432
rect 445720 179392 445726 179404
rect 13722 179324 13728 179376
rect 13780 179364 13786 179376
rect 64874 179364 64880 179376
rect 13780 179336 64880 179364
rect 13780 179324 13786 179336
rect 64874 179324 64880 179336
rect 64932 179324 64938 179376
rect 95142 179324 95148 179376
rect 95200 179364 95206 179376
rect 146294 179364 146300 179376
rect 95200 179336 146300 179364
rect 95200 179324 95206 179336
rect 146294 179324 146300 179336
rect 146352 179324 146358 179376
rect 148962 179324 148968 179376
rect 149020 179364 149026 179376
rect 200114 179364 200120 179376
rect 149020 179336 200120 179364
rect 149020 179324 149026 179336
rect 200114 179324 200120 179336
rect 200172 179324 200178 179376
rect 202782 179324 202788 179376
rect 202840 179364 202846 179376
rect 253934 179364 253940 179376
rect 202840 179336 253940 179364
rect 202840 179324 202846 179336
rect 253934 179324 253940 179336
rect 253992 179324 253998 179376
rect 256602 179324 256608 179376
rect 256660 179364 256666 179376
rect 307754 179364 307760 179376
rect 256660 179336 307760 179364
rect 256660 179324 256666 179336
rect 307754 179324 307760 179336
rect 307812 179324 307818 179376
rect 338022 179324 338028 179376
rect 338080 179364 338086 179376
rect 389174 179364 389180 179376
rect 338080 179336 389180 179364
rect 338080 179324 338086 179336
rect 389174 179324 389180 179336
rect 389232 179324 389238 179376
rect 391842 179324 391848 179376
rect 391900 179364 391906 179376
rect 442994 179364 443000 179376
rect 391900 179336 443000 179364
rect 391900 179324 391906 179336
rect 442994 179324 443000 179336
rect 443052 179324 443058 179376
rect 446398 179324 446404 179376
rect 446456 179364 446462 179376
rect 447686 179364 447692 179376
rect 446456 179336 447692 179364
rect 446456 179324 446462 179336
rect 447686 179324 447692 179336
rect 447744 179324 447750 179376
rect 454006 179364 454034 179404
rect 521746 179392 521752 179444
rect 521804 179432 521810 179444
rect 522390 179432 522396 179444
rect 521804 179404 522396 179432
rect 521804 179392 521810 179404
rect 522390 179392 522396 179404
rect 522448 179392 522454 179444
rect 496814 179364 496820 179376
rect 454006 179336 496820 179364
rect 496814 179324 496820 179336
rect 496872 179324 496878 179376
rect 500862 179324 500868 179376
rect 500920 179364 500926 179376
rect 550634 179364 550640 179376
rect 500920 179336 550640 179364
rect 500920 179324 500926 179336
rect 550634 179324 550640 179336
rect 550692 179324 550698 179376
rect 35618 179256 35624 179308
rect 35676 179296 35682 179308
rect 36722 179296 36728 179308
rect 35676 179268 36728 179296
rect 35676 179256 35682 179268
rect 36722 179256 36728 179268
rect 36780 179256 36786 179308
rect 41322 179256 41328 179308
rect 41380 179296 41386 179308
rect 91094 179296 91100 179308
rect 41380 179268 91100 179296
rect 41380 179256 41386 179268
rect 91094 179256 91100 179268
rect 91152 179256 91158 179308
rect 122742 179256 122748 179308
rect 122800 179296 122806 179308
rect 172514 179296 172520 179308
rect 122800 179268 172520 179296
rect 122800 179256 122806 179268
rect 172514 179256 172520 179268
rect 172572 179256 172578 179308
rect 176562 179256 176568 179308
rect 176620 179296 176626 179308
rect 226334 179296 226340 179308
rect 176620 179268 226340 179296
rect 176620 179256 176626 179268
rect 226334 179256 226340 179268
rect 226392 179256 226398 179308
rect 230382 179256 230388 179308
rect 230440 179296 230446 179308
rect 280154 179296 280160 179308
rect 230440 179268 280160 179296
rect 230440 179256 230446 179268
rect 280154 179256 280160 179268
rect 280212 179256 280218 179308
rect 284202 179256 284208 179308
rect 284260 179296 284266 179308
rect 335354 179296 335360 179308
rect 284260 179268 335360 179296
rect 284260 179256 284266 179268
rect 335354 179256 335360 179268
rect 335412 179256 335418 179308
rect 365622 179256 365628 179308
rect 365680 179296 365686 179308
rect 415394 179296 415400 179308
rect 365680 179268 415400 179296
rect 365680 179256 365686 179268
rect 415394 179256 415400 179268
rect 415452 179256 415458 179308
rect 419442 179256 419448 179308
rect 419500 179296 419506 179308
rect 469214 179296 469220 179308
rect 419500 179268 444374 179296
rect 419500 179256 419506 179268
rect 68922 179188 68928 179240
rect 68980 179228 68986 179240
rect 118694 179228 118700 179240
rect 68980 179200 118700 179228
rect 68980 179188 68986 179200
rect 118694 179188 118700 179200
rect 118752 179188 118758 179240
rect 311802 179188 311808 179240
rect 311860 179228 311866 179240
rect 361574 179228 361580 179240
rect 311860 179200 361580 179228
rect 311860 179188 311866 179200
rect 361574 179188 361580 179200
rect 361632 179188 361638 179240
rect 444346 179160 444374 179268
rect 456766 179268 469220 179296
rect 456766 179160 456794 179268
rect 469214 179256 469220 179268
rect 469272 179256 469278 179308
rect 473262 179256 473268 179308
rect 473320 179296 473326 179308
rect 523034 179296 523040 179308
rect 473320 179268 523040 179296
rect 473320 179256 473326 179268
rect 523034 179256 523040 179268
rect 523092 179256 523098 179308
rect 467650 179188 467656 179240
rect 467708 179228 467714 179240
rect 468570 179228 468576 179240
rect 467708 179200 468576 179228
rect 467708 179188 467714 179200
rect 468570 179188 468576 179200
rect 468628 179188 468634 179240
rect 444346 179132 456794 179160
rect 62758 176604 62764 176656
rect 62816 176644 62822 176656
rect 69750 176644 69756 176656
rect 62816 176616 69756 176644
rect 62816 176604 62822 176616
rect 69750 176604 69756 176616
rect 69808 176604 69814 176656
rect 96706 176604 96712 176656
rect 96764 176644 96770 176656
rect 96764 176616 103514 176644
rect 96764 176604 96770 176616
rect 15194 176536 15200 176588
rect 15252 176576 15258 176588
rect 42794 176576 42800 176588
rect 15252 176548 42800 176576
rect 15252 176536 15258 176548
rect 42794 176536 42800 176548
rect 42852 176536 42858 176588
rect 53098 176536 53104 176588
rect 53156 176576 53162 176588
rect 64138 176576 64144 176588
rect 53156 176548 64144 176576
rect 53156 176536 53162 176548
rect 64138 176536 64144 176548
rect 64196 176536 64202 176588
rect 69106 176536 69112 176588
rect 69164 176576 69170 176588
rect 96798 176576 96804 176588
rect 69164 176548 96804 176576
rect 69164 176536 69170 176548
rect 96798 176536 96804 176548
rect 96856 176536 96862 176588
rect 103486 176576 103514 176616
rect 146938 176604 146944 176656
rect 146996 176644 147002 176656
rect 146996 176616 151814 176644
rect 146996 176604 147002 176616
rect 123662 176576 123668 176588
rect 103486 176548 123668 176576
rect 123662 176536 123668 176548
rect 123720 176536 123726 176588
rect 133782 176536 133788 176588
rect 133840 176576 133846 176588
rect 144270 176576 144276 176588
rect 133840 176548 144276 176576
rect 133840 176536 133846 176548
rect 144270 176536 144276 176548
rect 144328 176536 144334 176588
rect 150526 176536 150532 176588
rect 150584 176576 150590 176588
rect 151786 176576 151814 176616
rect 200758 176604 200764 176656
rect 200816 176644 200822 176656
rect 204622 176644 204628 176656
rect 200816 176616 204628 176644
rect 200816 176604 200822 176616
rect 204622 176604 204628 176616
rect 204680 176604 204686 176656
rect 251818 176604 251824 176656
rect 251876 176644 251882 176656
rect 258718 176644 258724 176656
rect 251876 176616 258724 176644
rect 251876 176604 251882 176616
rect 258718 176604 258724 176616
rect 258776 176604 258782 176656
rect 332502 176604 332508 176656
rect 332560 176644 332566 176656
rect 335998 176644 336004 176656
rect 332560 176616 336004 176644
rect 332560 176604 332566 176616
rect 335998 176604 336004 176616
rect 336056 176604 336062 176656
rect 494698 176604 494704 176656
rect 494756 176644 494762 176656
rect 501598 176644 501604 176656
rect 494756 176616 501604 176644
rect 494756 176604 494762 176616
rect 501598 176604 501604 176616
rect 501656 176604 501662 176656
rect 547966 176576 547972 176588
rect 150584 176548 150940 176576
rect 151786 176548 547972 176576
rect 150584 176536 150590 176548
rect 26050 176468 26056 176520
rect 26108 176508 26114 176520
rect 36814 176508 36820 176520
rect 26108 176480 36820 176508
rect 26108 176468 26114 176480
rect 36814 176468 36820 176480
rect 36872 176468 36878 176520
rect 79962 176468 79968 176520
rect 80020 176508 80026 176520
rect 90450 176508 90456 176520
rect 80020 176480 90456 176508
rect 80020 176468 80026 176480
rect 90450 176468 90456 176480
rect 90508 176468 90514 176520
rect 106550 176468 106556 176520
rect 106608 176508 106614 176520
rect 116578 176508 116584 176520
rect 106608 176480 116584 176508
rect 106608 176468 106614 176480
rect 116578 176468 116584 176480
rect 116636 176468 116642 176520
rect 122926 176468 122932 176520
rect 122984 176508 122990 176520
rect 150710 176508 150716 176520
rect 122984 176480 150716 176508
rect 122984 176468 122990 176480
rect 150710 176468 150716 176480
rect 150768 176468 150774 176520
rect 150912 176508 150940 176548
rect 547966 176536 547972 176548
rect 548024 176536 548030 176588
rect 178126 176508 178132 176520
rect 150912 176480 178132 176508
rect 178126 176468 178132 176480
rect 178184 176468 178190 176520
rect 187970 176468 187976 176520
rect 188028 176508 188034 176520
rect 199378 176508 199384 176520
rect 188028 176480 199384 176508
rect 188028 176468 188034 176480
rect 199378 176468 199384 176480
rect 199436 176468 199442 176520
rect 204346 176468 204352 176520
rect 204404 176508 204410 176520
rect 231854 176508 231860 176520
rect 204404 176480 231860 176508
rect 204404 176468 204410 176480
rect 231854 176468 231860 176480
rect 231912 176468 231918 176520
rect 242066 176468 242072 176520
rect 242124 176508 242130 176520
rect 253198 176508 253204 176520
rect 242124 176480 253204 176508
rect 242124 176468 242130 176480
rect 253198 176468 253204 176480
rect 253256 176468 253262 176520
rect 258166 176468 258172 176520
rect 258224 176508 258230 176520
rect 286134 176508 286140 176520
rect 258224 176480 286140 176508
rect 258224 176468 258230 176480
rect 286134 176468 286140 176480
rect 286192 176468 286198 176520
rect 312630 176508 312636 176520
rect 287026 176480 312636 176508
rect 160554 176400 160560 176452
rect 160612 176440 160618 176452
rect 171778 176440 171784 176452
rect 160612 176412 171784 176440
rect 160612 176400 160618 176412
rect 171778 176400 171784 176412
rect 171836 176400 171842 176452
rect 215018 176400 215024 176452
rect 215076 176440 215082 176452
rect 225598 176440 225604 176452
rect 215076 176412 225604 176440
rect 215076 176400 215082 176412
rect 225598 176400 225604 176412
rect 225656 176400 225662 176452
rect 268930 176400 268936 176452
rect 268988 176440 268994 176452
rect 279510 176440 279516 176452
rect 268988 176412 279516 176440
rect 268988 176400 268994 176412
rect 279510 176400 279516 176412
rect 279568 176400 279574 176452
rect 285766 176400 285772 176452
rect 285824 176440 285830 176452
rect 287026 176440 287054 176480
rect 312630 176468 312636 176480
rect 312688 176468 312694 176520
rect 340138 176508 340144 176520
rect 316006 176480 340144 176508
rect 285824 176412 287054 176440
rect 285824 176400 285830 176412
rect 295978 176400 295984 176452
rect 296036 176440 296042 176452
rect 307018 176440 307024 176452
rect 296036 176412 307024 176440
rect 296036 176400 296042 176412
rect 307018 176400 307024 176412
rect 307076 176400 307082 176452
rect 311986 176400 311992 176452
rect 312044 176440 312050 176452
rect 316006 176440 316034 176480
rect 340138 176468 340144 176480
rect 340196 176468 340202 176520
rect 366726 176508 366732 176520
rect 344986 176480 366732 176508
rect 312044 176412 316034 176440
rect 312044 176400 312050 176412
rect 322842 176400 322848 176452
rect 322900 176440 322906 176452
rect 333238 176440 333244 176452
rect 322900 176412 333244 176440
rect 322900 176400 322906 176412
rect 333238 176400 333244 176412
rect 333296 176400 333302 176452
rect 339586 176400 339592 176452
rect 339644 176440 339650 176452
rect 344986 176440 345014 176480
rect 366726 176468 366732 176480
rect 366784 176468 366790 176520
rect 393590 176508 393596 176520
rect 373966 176480 393596 176508
rect 339644 176412 345014 176440
rect 339644 176400 339650 176412
rect 350074 176400 350080 176452
rect 350132 176440 350138 176452
rect 359550 176440 359556 176452
rect 350132 176412 359556 176440
rect 350132 176400 350138 176412
rect 359550 176400 359556 176412
rect 359608 176400 359614 176452
rect 365806 176400 365812 176452
rect 365864 176440 365870 176452
rect 373966 176440 373994 176480
rect 393590 176468 393596 176480
rect 393648 176468 393654 176520
rect 420914 176508 420920 176520
rect 402946 176480 420920 176508
rect 365864 176412 373994 176440
rect 365864 176400 365870 176412
rect 376570 176400 376576 176452
rect 376628 176440 376634 176452
rect 387058 176440 387064 176452
rect 376628 176412 387064 176440
rect 376628 176400 376634 176412
rect 387058 176400 387064 176412
rect 387116 176400 387122 176452
rect 393406 176400 393412 176452
rect 393464 176440 393470 176452
rect 402946 176440 402974 176480
rect 420914 176468 420920 176480
rect 420972 176468 420978 176520
rect 431034 176468 431040 176520
rect 431092 176508 431098 176520
rect 442258 176508 442264 176520
rect 431092 176480 442264 176508
rect 431092 176468 431098 176480
rect 442258 176468 442264 176480
rect 442316 176468 442322 176520
rect 447226 176468 447232 176520
rect 447284 176508 447290 176520
rect 474734 176508 474740 176520
rect 447284 176480 474740 176508
rect 447284 176468 447290 176480
rect 474734 176468 474740 176480
rect 474792 176468 474798 176520
rect 484946 176468 484952 176520
rect 485004 176508 485010 176520
rect 496078 176508 496084 176520
rect 485004 176480 496084 176508
rect 485004 176468 485010 176480
rect 496078 176468 496084 176480
rect 496136 176468 496142 176520
rect 501046 176468 501052 176520
rect 501104 176508 501110 176520
rect 528646 176508 528652 176520
rect 501104 176480 528652 176508
rect 501104 176468 501110 176480
rect 528646 176468 528652 176480
rect 528704 176468 528710 176520
rect 393464 176412 402974 176440
rect 393464 176400 393470 176412
rect 403986 176400 403992 176452
rect 404044 176440 404050 176452
rect 414658 176440 414664 176452
rect 404044 176412 414664 176440
rect 404044 176400 404050 176412
rect 414658 176400 414664 176412
rect 414716 176400 414722 176452
rect 458082 176400 458088 176452
rect 458140 176440 458146 176452
rect 468478 176440 468484 176452
rect 458140 176412 468484 176440
rect 458140 176400 458146 176412
rect 468478 176400 468484 176412
rect 468536 176400 468542 176452
rect 511902 176400 511908 176452
rect 511960 176440 511966 176452
rect 522298 176440 522304 176452
rect 511960 176412 522304 176440
rect 511960 176400 511966 176412
rect 522298 176400 522304 176412
rect 522356 176400 522362 176452
rect 36630 176332 36636 176384
rect 36688 176372 36694 176384
rect 538398 176372 538404 176384
rect 36688 176344 538404 176372
rect 36688 176332 36694 176344
rect 538398 176332 538404 176344
rect 538456 176332 538462 176384
rect 16298 173136 16304 173188
rect 16356 173176 16362 173188
rect 528646 173176 528652 173188
rect 16356 173148 528652 173176
rect 16356 173136 16362 173148
rect 528646 173136 528652 173148
rect 528704 173136 528710 173188
rect 26050 172796 26056 172848
rect 26108 172836 26114 172848
rect 146938 172836 146944 172848
rect 26108 172808 146944 172836
rect 26108 172796 26114 172808
rect 146938 172796 146944 172808
rect 146996 172796 147002 172848
rect 36722 172728 36728 172780
rect 36780 172768 36786 172780
rect 52454 172768 52460 172780
rect 36780 172740 52460 172768
rect 36780 172728 36786 172740
rect 52454 172728 52460 172740
rect 52512 172728 52518 172780
rect 232314 172728 232320 172780
rect 232372 172768 232378 172780
rect 251818 172768 251824 172780
rect 232372 172740 251824 172768
rect 232372 172728 232378 172740
rect 251818 172728 251824 172740
rect 251876 172728 251882 172780
rect 475378 172728 475384 172780
rect 475436 172768 475442 172780
rect 494698 172768 494704 172780
rect 475436 172740 494704 172768
rect 475436 172728 475442 172740
rect 494698 172728 494704 172740
rect 494756 172728 494762 172780
rect 62482 172660 62488 172712
rect 62540 172700 62546 172712
rect 79318 172700 79324 172712
rect 62540 172672 79324 172700
rect 62540 172660 62546 172672
rect 79318 172660 79324 172672
rect 79376 172660 79382 172712
rect 90450 172660 90456 172712
rect 90508 172700 90514 172712
rect 106458 172700 106464 172712
rect 90508 172672 106464 172700
rect 90508 172660 90514 172672
rect 106458 172660 106464 172672
rect 106516 172660 106522 172712
rect 116486 172660 116492 172712
rect 116544 172700 116550 172712
rect 133414 172700 133420 172712
rect 116544 172672 133420 172700
rect 116544 172660 116550 172672
rect 133414 172660 133420 172672
rect 133472 172660 133478 172712
rect 170490 172660 170496 172712
rect 170548 172700 170554 172712
rect 187786 172700 187792 172712
rect 170548 172672 187792 172700
rect 170548 172660 170554 172672
rect 187786 172660 187792 172672
rect 187844 172660 187850 172712
rect 197538 172660 197544 172712
rect 197596 172700 197602 172712
rect 214374 172700 214380 172712
rect 197596 172672 214380 172700
rect 197596 172660 197602 172672
rect 214374 172660 214380 172672
rect 214432 172660 214438 172712
rect 224494 172660 224500 172712
rect 224552 172700 224558 172712
rect 241606 172700 241612 172712
rect 224552 172672 241612 172700
rect 224552 172660 224558 172672
rect 241606 172660 241612 172672
rect 241664 172660 241670 172712
rect 413462 172660 413468 172712
rect 413520 172700 413526 172712
rect 430574 172700 430580 172712
rect 413520 172672 430580 172700
rect 413520 172660 413526 172672
rect 430574 172660 430580 172672
rect 430632 172660 430638 172712
rect 440510 172660 440516 172712
rect 440568 172700 440574 172712
rect 457254 172700 457260 172712
rect 440568 172672 457260 172700
rect 440568 172660 440574 172672
rect 457254 172660 457260 172672
rect 457312 172660 457318 172712
rect 468478 172660 468484 172712
rect 468536 172700 468542 172712
rect 484394 172700 484400 172712
rect 468536 172672 484400 172700
rect 468536 172660 468542 172672
rect 484394 172660 484400 172672
rect 484452 172660 484458 172712
rect 36814 172592 36820 172644
rect 36872 172632 36878 172644
rect 62114 172632 62120 172644
rect 36872 172604 62120 172632
rect 36872 172592 36878 172604
rect 62114 172592 62120 172604
rect 62172 172592 62178 172644
rect 64138 172592 64144 172644
rect 64196 172632 64202 172644
rect 89070 172632 89076 172644
rect 64196 172604 89076 172632
rect 64196 172592 64202 172604
rect 89070 172592 89076 172604
rect 89128 172592 89134 172644
rect 90358 172592 90364 172644
rect 90416 172632 90422 172644
rect 116118 172632 116124 172644
rect 90416 172604 116124 172632
rect 90416 172592 90422 172604
rect 116118 172592 116124 172604
rect 116176 172592 116182 172644
rect 116578 172592 116584 172644
rect 116636 172632 116642 172644
rect 142982 172632 142988 172644
rect 116636 172604 142988 172632
rect 116636 172592 116642 172604
rect 142982 172592 142988 172604
rect 143040 172592 143046 172644
rect 144178 172592 144184 172644
rect 144236 172632 144242 172644
rect 170030 172632 170036 172644
rect 144236 172604 170036 172632
rect 144236 172592 144242 172604
rect 170030 172592 170036 172604
rect 170088 172592 170094 172644
rect 178402 172592 178408 172644
rect 178460 172632 178466 172644
rect 200758 172632 200764 172644
rect 178460 172604 200764 172632
rect 178460 172592 178466 172604
rect 200758 172592 200764 172604
rect 200816 172592 200822 172644
rect 251450 172592 251456 172644
rect 251508 172632 251514 172644
rect 268286 172632 268292 172644
rect 251508 172604 268292 172632
rect 251508 172592 251514 172604
rect 268286 172592 268292 172604
rect 268344 172592 268350 172644
rect 279418 172592 279424 172644
rect 279476 172632 279482 172644
rect 295794 172632 295800 172644
rect 279476 172604 295800 172632
rect 279476 172592 279482 172604
rect 295794 172592 295800 172604
rect 295852 172592 295858 172644
rect 305546 172592 305552 172644
rect 305604 172632 305610 172644
rect 322382 172632 322388 172644
rect 305604 172604 322388 172632
rect 305604 172592 305610 172604
rect 322382 172592 322388 172604
rect 322440 172592 322446 172644
rect 334618 172592 334624 172644
rect 334676 172632 334682 172644
rect 349798 172632 349804 172644
rect 334676 172604 349804 172632
rect 334676 172592 334682 172604
rect 349798 172592 349804 172604
rect 349856 172592 349862 172644
rect 359642 172592 359648 172644
rect 359700 172632 359706 172644
rect 376294 172632 376300 172644
rect 359700 172604 376300 172632
rect 359700 172592 359706 172604
rect 376294 172592 376300 172604
rect 376352 172592 376358 172644
rect 386506 172592 386512 172644
rect 386564 172632 386570 172644
rect 403342 172632 403348 172644
rect 386564 172604 403348 172632
rect 386564 172592 386570 172604
rect 403342 172592 403348 172604
rect 403400 172592 403406 172644
rect 421282 172592 421288 172644
rect 421340 172632 421346 172644
rect 443638 172632 443644 172644
rect 421340 172604 443644 172632
rect 421340 172592 421346 172604
rect 443638 172592 443644 172604
rect 443696 172592 443702 172644
rect 494514 172592 494520 172644
rect 494572 172632 494578 172644
rect 511350 172632 511356 172644
rect 494572 172604 511356 172632
rect 494572 172592 494578 172604
rect 511350 172592 511356 172604
rect 511408 172592 511414 172644
rect 522298 172592 522304 172644
rect 522356 172632 522362 172644
rect 538398 172632 538404 172644
rect 522356 172604 538404 172632
rect 522356 172592 522362 172604
rect 538398 172592 538404 172604
rect 538456 172592 538462 172644
rect 43346 172524 43352 172576
rect 43404 172564 43410 172576
rect 62758 172564 62764 172576
rect 43404 172536 62764 172564
rect 43404 172524 43410 172536
rect 62758 172524 62764 172536
rect 62816 172524 62822 172576
rect 144270 172524 144276 172576
rect 144328 172564 144334 172576
rect 160278 172564 160284 172576
rect 144328 172536 160284 172564
rect 144328 172524 144334 172536
rect 160278 172524 160284 172536
rect 160336 172524 160342 172576
rect 171778 172524 171784 172576
rect 171836 172564 171842 172576
rect 197446 172564 197452 172576
rect 171836 172536 197452 172564
rect 171836 172524 171842 172536
rect 197446 172524 197452 172536
rect 197504 172524 197510 172576
rect 199378 172524 199384 172576
rect 199436 172564 199442 172576
rect 223942 172564 223948 172576
rect 199436 172536 223948 172564
rect 199436 172524 199442 172536
rect 223942 172524 223948 172536
rect 224000 172524 224006 172576
rect 225598 172524 225604 172576
rect 225656 172564 225662 172576
rect 251266 172564 251272 172576
rect 225656 172536 251272 172564
rect 225656 172524 225662 172536
rect 251266 172524 251272 172536
rect 251324 172524 251330 172576
rect 253198 172524 253204 172576
rect 253256 172564 253262 172576
rect 278038 172564 278044 172576
rect 253256 172536 278044 172564
rect 253256 172524 253262 172536
rect 278038 172524 278044 172536
rect 278096 172524 278102 172576
rect 279510 172524 279516 172576
rect 279568 172564 279574 172576
rect 305454 172564 305460 172576
rect 279568 172536 305460 172564
rect 279568 172524 279574 172536
rect 305454 172524 305460 172536
rect 305512 172524 305518 172576
rect 307018 172524 307024 172576
rect 307076 172564 307082 172576
rect 331950 172564 331956 172576
rect 307076 172536 331956 172564
rect 307076 172524 307082 172536
rect 331950 172524 331956 172536
rect 332008 172524 332014 172576
rect 333238 172524 333244 172576
rect 333296 172564 333302 172576
rect 359458 172564 359464 172576
rect 333296 172536 359464 172564
rect 333296 172524 333302 172536
rect 359458 172524 359464 172536
rect 359516 172524 359522 172576
rect 359550 172524 359556 172576
rect 359608 172564 359614 172576
rect 386046 172564 386052 172576
rect 359608 172536 386052 172564
rect 359608 172524 359614 172536
rect 386046 172524 386052 172536
rect 386104 172524 386110 172576
rect 387058 172524 387064 172576
rect 387116 172564 387122 172576
rect 412910 172564 412916 172576
rect 387116 172536 412916 172564
rect 387116 172524 387122 172536
rect 412910 172524 412916 172536
rect 412968 172524 412974 172576
rect 414658 172524 414664 172576
rect 414716 172564 414722 172576
rect 440234 172564 440240 172576
rect 414716 172536 440240 172564
rect 414716 172524 414722 172536
rect 440234 172524 440240 172536
rect 440292 172524 440298 172576
rect 442258 172524 442264 172576
rect 442316 172564 442322 172576
rect 467006 172564 467012 172576
rect 442316 172536 467012 172564
rect 442316 172524 442322 172536
rect 467006 172524 467012 172536
rect 467064 172524 467070 172576
rect 468570 172524 468576 172576
rect 468628 172564 468634 172576
rect 494054 172564 494060 172576
rect 468628 172536 494060 172564
rect 468628 172524 468634 172536
rect 494054 172524 494060 172536
rect 494112 172524 494118 172576
rect 496078 172524 496084 172576
rect 496136 172564 496142 172576
rect 520918 172564 520924 172576
rect 496136 172536 520924 172564
rect 496136 172524 496142 172536
rect 520918 172524 520924 172536
rect 520976 172524 520982 172576
rect 522390 172524 522396 172576
rect 522448 172564 522454 172576
rect 547966 172564 547972 172576
rect 522448 172536 547972 172564
rect 522448 172524 522454 172536
rect 547966 172524 547972 172536
rect 548024 172524 548030 172576
rect 37918 170348 37924 170400
rect 37976 170388 37982 170400
rect 526438 170388 526444 170400
rect 37976 170360 526444 170388
rect 37976 170348 37982 170360
rect 526438 170348 526444 170360
rect 526496 170348 526502 170400
rect 285766 170280 285772 170332
rect 285824 170320 285830 170332
rect 286134 170320 286140 170332
rect 285824 170292 286140 170320
rect 285824 170280 285830 170292
rect 286134 170280 286140 170292
rect 286192 170280 286198 170332
rect 339586 170280 339592 170332
rect 339644 170320 339650 170332
rect 340138 170320 340144 170332
rect 339644 170292 340144 170320
rect 339644 170280 339650 170292
rect 340138 170280 340144 170292
rect 340196 170280 340202 170332
rect 35618 169736 35624 169788
rect 35676 169776 35682 169788
rect 36630 169776 36636 169788
rect 35676 169748 36636 169776
rect 35676 169736 35682 169748
rect 36630 169736 36636 169748
rect 36688 169736 36694 169788
rect 359550 166336 359556 166388
rect 359608 166336 359614 166388
rect 359568 166184 359596 166336
rect 359550 166132 359556 166184
rect 359608 166132 359614 166184
rect 89714 156612 89720 156664
rect 89772 156652 89778 156664
rect 90450 156652 90456 156664
rect 89772 156624 90456 156652
rect 89772 156612 89778 156624
rect 90450 156612 90456 156624
rect 90508 156612 90514 156664
rect 143626 154300 143632 154352
rect 143684 154340 143690 154352
rect 144270 154340 144276 154352
rect 143684 154312 144276 154340
rect 143684 154300 143690 154312
rect 144270 154300 144276 154312
rect 144328 154300 144334 154352
rect 13722 151716 13728 151768
rect 13780 151756 13786 151768
rect 64874 151756 64880 151768
rect 13780 151728 64880 151756
rect 13780 151716 13786 151728
rect 64874 151716 64880 151728
rect 64932 151716 64938 151768
rect 95142 151716 95148 151768
rect 95200 151756 95206 151768
rect 146294 151756 146300 151768
rect 95200 151728 146300 151756
rect 95200 151716 95206 151728
rect 146294 151716 146300 151728
rect 146352 151716 146358 151768
rect 148962 151716 148968 151768
rect 149020 151756 149026 151768
rect 200114 151756 200120 151768
rect 149020 151728 200120 151756
rect 149020 151716 149026 151728
rect 200114 151716 200120 151728
rect 200172 151716 200178 151768
rect 202782 151716 202788 151768
rect 202840 151756 202846 151768
rect 253934 151756 253940 151768
rect 202840 151728 253940 151756
rect 202840 151716 202846 151728
rect 253934 151716 253940 151728
rect 253992 151716 253998 151768
rect 256602 151716 256608 151768
rect 256660 151756 256666 151768
rect 307754 151756 307760 151768
rect 256660 151728 307760 151756
rect 256660 151716 256666 151728
rect 307754 151716 307760 151728
rect 307812 151716 307818 151768
rect 332502 151716 332508 151768
rect 332560 151756 332566 151768
rect 334618 151756 334624 151768
rect 332560 151728 334624 151756
rect 332560 151716 332566 151728
rect 334618 151716 334624 151728
rect 334676 151716 334682 151768
rect 338022 151716 338028 151768
rect 338080 151756 338086 151768
rect 389174 151756 389180 151768
rect 338080 151728 389180 151756
rect 338080 151716 338086 151728
rect 389174 151716 389180 151728
rect 389232 151716 389238 151768
rect 391842 151716 391848 151768
rect 391900 151756 391906 151768
rect 442994 151756 443000 151768
rect 391900 151728 443000 151756
rect 391900 151716 391906 151728
rect 442994 151716 443000 151728
rect 443052 151716 443058 151768
rect 445662 151716 445668 151768
rect 445720 151756 445726 151768
rect 496814 151756 496820 151768
rect 445720 151728 496820 151756
rect 445720 151716 445726 151728
rect 496814 151716 496820 151728
rect 496872 151716 496878 151768
rect 500862 151716 500868 151768
rect 500920 151756 500926 151768
rect 550634 151756 550640 151768
rect 500920 151728 550640 151756
rect 500920 151716 500926 151728
rect 550634 151716 550640 151728
rect 550692 151716 550698 151768
rect 35618 151648 35624 151700
rect 35676 151688 35682 151700
rect 36722 151688 36728 151700
rect 35676 151660 36728 151688
rect 35676 151648 35682 151660
rect 36722 151648 36728 151660
rect 36780 151648 36786 151700
rect 41322 151648 41328 151700
rect 41380 151688 41386 151700
rect 91094 151688 91100 151700
rect 41380 151660 91100 151688
rect 41380 151648 41386 151660
rect 91094 151648 91100 151660
rect 91152 151648 91158 151700
rect 122742 151648 122748 151700
rect 122800 151688 122806 151700
rect 172514 151688 172520 151700
rect 122800 151660 172520 151688
rect 122800 151648 122806 151660
rect 172514 151648 172520 151660
rect 172572 151648 172578 151700
rect 176562 151648 176568 151700
rect 176620 151688 176626 151700
rect 226334 151688 226340 151700
rect 176620 151660 226340 151688
rect 176620 151648 176626 151660
rect 226334 151648 226340 151660
rect 226392 151648 226398 151700
rect 230382 151648 230388 151700
rect 230440 151688 230446 151700
rect 280154 151688 280160 151700
rect 230440 151660 280160 151688
rect 230440 151648 230446 151660
rect 280154 151648 280160 151660
rect 280212 151648 280218 151700
rect 284202 151648 284208 151700
rect 284260 151688 284266 151700
rect 335354 151688 335360 151700
rect 284260 151660 335360 151688
rect 284260 151648 284266 151660
rect 335354 151648 335360 151660
rect 335412 151648 335418 151700
rect 365622 151648 365628 151700
rect 365680 151688 365686 151700
rect 415394 151688 415400 151700
rect 365680 151660 415400 151688
rect 365680 151648 365686 151660
rect 415394 151648 415400 151660
rect 415452 151648 415458 151700
rect 419442 151648 419448 151700
rect 419500 151688 419506 151700
rect 469214 151688 469220 151700
rect 419500 151660 469220 151688
rect 419500 151648 419506 151660
rect 469214 151648 469220 151660
rect 469272 151648 469278 151700
rect 473262 151648 473268 151700
rect 473320 151688 473326 151700
rect 523034 151688 523040 151700
rect 473320 151660 523040 151688
rect 473320 151648 473326 151660
rect 523034 151648 523040 151660
rect 523092 151648 523098 151700
rect 68922 151580 68928 151632
rect 68980 151620 68986 151632
rect 118694 151620 118700 151632
rect 68980 151592 118700 151620
rect 68980 151580 68986 151592
rect 118694 151580 118700 151592
rect 118752 151580 118758 151632
rect 200758 151580 200764 151632
rect 200816 151620 200822 151632
rect 204622 151620 204628 151632
rect 200816 151592 204628 151620
rect 200816 151580 200822 151592
rect 204622 151580 204628 151592
rect 204680 151580 204686 151632
rect 311802 151580 311808 151632
rect 311860 151620 311866 151632
rect 361574 151620 361580 151632
rect 311860 151592 361580 151620
rect 311860 151580 311866 151592
rect 361574 151580 361580 151592
rect 361632 151580 361638 151632
rect 443638 151580 443644 151632
rect 443696 151620 443702 151632
rect 447686 151620 447692 151632
rect 443696 151592 447692 151620
rect 443696 151580 443702 151592
rect 447686 151580 447692 151592
rect 447744 151580 447750 151632
rect 52730 148996 52736 149048
rect 52788 149036 52794 149048
rect 64138 149036 64144 149048
rect 52788 149008 64144 149036
rect 52788 148996 52794 149008
rect 64138 148996 64144 149008
rect 64196 148996 64202 149048
rect 69106 148996 69112 149048
rect 69164 149036 69170 149048
rect 69164 149008 74534 149036
rect 69164 148996 69170 149008
rect 15194 148928 15200 148980
rect 15252 148968 15258 148980
rect 42978 148968 42984 148980
rect 15252 148940 42984 148968
rect 15252 148928 15258 148940
rect 42978 148928 42984 148940
rect 43036 148928 43042 148980
rect 62758 148928 62764 148980
rect 62816 148968 62822 148980
rect 70026 148968 70032 148980
rect 62816 148940 70032 148968
rect 62816 148928 62822 148940
rect 70026 148928 70032 148940
rect 70084 148928 70090 148980
rect 74506 148968 74534 149008
rect 96706 148996 96712 149048
rect 96764 149036 96770 149048
rect 96764 149008 103514 149036
rect 96764 148996 96770 149008
rect 96982 148968 96988 148980
rect 74506 148940 96988 148968
rect 96982 148928 96988 148940
rect 97040 148928 97046 148980
rect 103486 148968 103514 149008
rect 251818 148996 251824 149048
rect 251876 149036 251882 149048
rect 258994 149036 259000 149048
rect 251876 149008 259000 149036
rect 251876 148996 251882 149008
rect 258994 148996 259000 149008
rect 259052 148996 259058 149048
rect 494698 148996 494704 149048
rect 494756 149036 494762 149048
rect 501966 149036 501972 149048
rect 494756 149008 501972 149036
rect 494756 148996 494762 149008
rect 501966 148996 501972 149008
rect 502024 148996 502030 149048
rect 124030 148968 124036 148980
rect 103486 148940 124036 148968
rect 124030 148928 124036 148940
rect 124088 148928 124094 148980
rect 149698 148928 149704 148980
rect 149756 148968 149762 148980
rect 548334 148968 548340 148980
rect 149756 148940 548340 148968
rect 149756 148928 149762 148940
rect 548334 148928 548340 148940
rect 548392 148928 548398 148980
rect 25682 148860 25688 148912
rect 25740 148900 25746 148912
rect 36814 148900 36820 148912
rect 25740 148872 36820 148900
rect 25740 148860 25746 148872
rect 36814 148860 36820 148872
rect 36872 148860 36878 148912
rect 79686 148860 79692 148912
rect 79744 148900 79750 148912
rect 90358 148900 90364 148912
rect 79744 148872 90364 148900
rect 79744 148860 79750 148872
rect 90358 148860 90364 148872
rect 90416 148860 90422 148912
rect 106642 148860 106648 148912
rect 106700 148900 106706 148912
rect 116578 148900 116584 148912
rect 106700 148872 116584 148900
rect 106700 148860 106706 148872
rect 116578 148860 116584 148872
rect 116636 148860 116642 148912
rect 133690 148860 133696 148912
rect 133748 148900 133754 148912
rect 144178 148900 144184 148912
rect 133748 148872 144184 148900
rect 133748 148860 133754 148872
rect 144178 148860 144184 148872
rect 144236 148860 144242 148912
rect 150526 148860 150532 148912
rect 150584 148900 150590 148912
rect 178034 148900 178040 148912
rect 150584 148872 178040 148900
rect 150584 148860 150590 148872
rect 178034 148860 178040 148872
rect 178092 148860 178098 148912
rect 187694 148860 187700 148912
rect 187752 148900 187758 148912
rect 199378 148900 199384 148912
rect 187752 148872 199384 148900
rect 187752 148860 187758 148872
rect 199378 148860 199384 148872
rect 199436 148860 199442 148912
rect 204346 148860 204352 148912
rect 204404 148900 204410 148912
rect 232038 148900 232044 148912
rect 204404 148872 232044 148900
rect 204404 148860 204410 148872
rect 232038 148860 232044 148872
rect 232096 148860 232102 148912
rect 241698 148860 241704 148912
rect 241756 148900 241762 148912
rect 253198 148900 253204 148912
rect 241756 148872 253204 148900
rect 241756 148860 241762 148872
rect 253198 148860 253204 148872
rect 253256 148860 253262 148912
rect 258166 148860 258172 148912
rect 258224 148900 258230 148912
rect 286042 148900 286048 148912
rect 258224 148872 286048 148900
rect 258224 148860 258230 148872
rect 286042 148860 286048 148872
rect 286100 148860 286106 148912
rect 312998 148900 313004 148912
rect 287026 148872 313004 148900
rect 122926 148792 122932 148844
rect 122984 148832 122990 148844
rect 150986 148832 150992 148844
rect 122984 148804 150992 148832
rect 122984 148792 122990 148804
rect 150986 148792 150992 148804
rect 151044 148792 151050 148844
rect 160646 148792 160652 148844
rect 160704 148832 160710 148844
rect 171778 148832 171784 148844
rect 160704 148804 171784 148832
rect 160704 148792 160710 148804
rect 171778 148792 171784 148804
rect 171836 148792 171842 148844
rect 214650 148792 214656 148844
rect 214708 148832 214714 148844
rect 225598 148832 225604 148844
rect 214708 148804 225604 148832
rect 214708 148792 214714 148804
rect 225598 148792 225604 148804
rect 225656 148792 225662 148844
rect 268654 148792 268660 148844
rect 268712 148832 268718 148844
rect 279510 148832 279516 148844
rect 268712 148804 279516 148832
rect 268712 148792 268718 148804
rect 279510 148792 279516 148804
rect 279568 148792 279574 148844
rect 285766 148792 285772 148844
rect 285824 148832 285830 148844
rect 287026 148832 287054 148872
rect 312998 148860 313004 148872
rect 313056 148860 313062 148912
rect 340046 148900 340052 148912
rect 316006 148872 340052 148900
rect 285824 148804 287054 148832
rect 285824 148792 285830 148804
rect 295702 148792 295708 148844
rect 295760 148832 295766 148844
rect 307018 148832 307024 148844
rect 295760 148804 307024 148832
rect 295760 148792 295766 148804
rect 307018 148792 307024 148804
rect 307076 148792 307082 148844
rect 311986 148792 311992 148844
rect 312044 148832 312050 148844
rect 316006 148832 316034 148872
rect 340046 148860 340052 148872
rect 340104 148860 340110 148912
rect 367002 148900 367008 148912
rect 344986 148872 367008 148900
rect 312044 148804 316034 148832
rect 312044 148792 312050 148804
rect 322658 148792 322664 148844
rect 322716 148832 322722 148844
rect 333238 148832 333244 148844
rect 322716 148804 333244 148832
rect 322716 148792 322722 148804
rect 333238 148792 333244 148804
rect 333296 148792 333302 148844
rect 339586 148792 339592 148844
rect 339644 148832 339650 148844
rect 344986 148832 345014 148872
rect 367002 148860 367008 148872
rect 367060 148860 367066 148912
rect 393958 148900 393964 148912
rect 373966 148872 393964 148900
rect 339644 148804 345014 148832
rect 339644 148792 339650 148804
rect 349706 148792 349712 148844
rect 349764 148832 349770 148844
rect 359550 148832 359556 148844
rect 349764 148804 359556 148832
rect 349764 148792 349770 148804
rect 359550 148792 359556 148804
rect 359608 148792 359614 148844
rect 365806 148792 365812 148844
rect 365864 148832 365870 148844
rect 373966 148832 373994 148872
rect 393958 148860 393964 148872
rect 394016 148860 394022 148912
rect 421006 148900 421012 148912
rect 402946 148872 421012 148900
rect 365864 148804 373994 148832
rect 365864 148792 365870 148804
rect 376662 148792 376668 148844
rect 376720 148832 376726 148844
rect 387058 148832 387064 148844
rect 376720 148804 387064 148832
rect 376720 148792 376726 148804
rect 387058 148792 387064 148804
rect 387116 148792 387122 148844
rect 393406 148792 393412 148844
rect 393464 148832 393470 148844
rect 402946 148832 402974 148872
rect 421006 148860 421012 148872
rect 421064 148860 421070 148912
rect 430666 148860 430672 148912
rect 430724 148900 430730 148912
rect 442258 148900 442264 148912
rect 430724 148872 442264 148900
rect 430724 148860 430730 148872
rect 442258 148860 442264 148872
rect 442316 148860 442322 148912
rect 447226 148860 447232 148912
rect 447284 148900 447290 148912
rect 475010 148900 475016 148912
rect 447284 148872 475016 148900
rect 447284 148860 447290 148872
rect 475010 148860 475016 148872
rect 475068 148860 475074 148912
rect 484670 148860 484676 148912
rect 484728 148900 484734 148912
rect 496078 148900 496084 148912
rect 484728 148872 496084 148900
rect 484728 148860 484734 148872
rect 496078 148860 496084 148872
rect 496136 148860 496142 148912
rect 501046 148860 501052 148912
rect 501104 148900 501110 148912
rect 529014 148900 529020 148912
rect 501104 148872 529020 148900
rect 501104 148860 501110 148872
rect 529014 148860 529020 148872
rect 529072 148860 529078 148912
rect 393464 148804 402974 148832
rect 393464 148792 393470 148804
rect 403710 148792 403716 148844
rect 403768 148832 403774 148844
rect 414658 148832 414664 148844
rect 403768 148804 414664 148832
rect 403768 148792 403774 148804
rect 414658 148792 414664 148804
rect 414716 148792 414722 148844
rect 457714 148792 457720 148844
rect 457772 148832 457778 148844
rect 468570 148832 468576 148844
rect 457772 148804 468576 148832
rect 457772 148792 457778 148804
rect 468570 148792 468576 148804
rect 468628 148792 468634 148844
rect 511718 148792 511724 148844
rect 511776 148832 511782 148844
rect 522390 148832 522396 148844
rect 511776 148804 522396 148832
rect 511776 148792 511782 148804
rect 522390 148792 522396 148804
rect 522448 148792 522454 148844
rect 36538 148724 36544 148776
rect 36596 148764 36602 148776
rect 538674 148764 538680 148776
rect 36596 148736 538680 148764
rect 36596 148724 36602 148736
rect 538674 148724 538680 148736
rect 538732 148724 538738 148776
rect 16022 146888 16028 146940
rect 16080 146928 16086 146940
rect 529014 146928 529020 146940
rect 16080 146900 529020 146928
rect 16080 146888 16086 146900
rect 529014 146888 529020 146900
rect 529072 146888 529078 146940
rect 25682 146548 25688 146600
rect 25740 146588 25746 146600
rect 149698 146588 149704 146600
rect 25740 146560 149704 146588
rect 25740 146548 25746 146560
rect 149698 146548 149704 146560
rect 149756 146548 149762 146600
rect 36722 146480 36728 146532
rect 36780 146520 36786 146532
rect 52638 146520 52644 146532
rect 36780 146492 52644 146520
rect 36780 146480 36786 146492
rect 52638 146480 52644 146492
rect 52696 146480 52702 146532
rect 232038 146480 232044 146532
rect 232096 146520 232102 146532
rect 251818 146520 251824 146532
rect 232096 146492 251824 146520
rect 232096 146480 232102 146492
rect 251818 146480 251824 146492
rect 251876 146480 251882 146532
rect 475010 146480 475016 146532
rect 475068 146520 475074 146532
rect 494698 146520 494704 146532
rect 475068 146492 494704 146520
rect 475068 146480 475074 146492
rect 494698 146480 494704 146492
rect 494756 146480 494762 146532
rect 62482 146412 62488 146464
rect 62540 146452 62546 146464
rect 79686 146452 79692 146464
rect 62540 146424 79692 146452
rect 62540 146412 62546 146424
rect 79686 146412 79692 146424
rect 79744 146412 79750 146464
rect 90450 146412 90456 146464
rect 90508 146452 90514 146464
rect 106642 146452 106648 146464
rect 90508 146424 106648 146452
rect 90508 146412 90514 146424
rect 106642 146412 106648 146424
rect 106700 146412 106706 146464
rect 116486 146412 116492 146464
rect 116544 146452 116550 146464
rect 133690 146452 133696 146464
rect 116544 146424 133696 146452
rect 116544 146412 116550 146424
rect 133690 146412 133696 146424
rect 133748 146412 133754 146464
rect 144178 146412 144184 146464
rect 144236 146452 144242 146464
rect 160646 146452 160652 146464
rect 144236 146424 160652 146452
rect 144236 146412 144242 146424
rect 160646 146412 160652 146424
rect 160704 146412 160710 146464
rect 170490 146412 170496 146464
rect 170548 146452 170554 146464
rect 187694 146452 187700 146464
rect 170548 146424 187700 146452
rect 170548 146412 170554 146424
rect 187694 146412 187700 146424
rect 187752 146412 187758 146464
rect 197446 146412 197452 146464
rect 197504 146452 197510 146464
rect 214650 146452 214656 146464
rect 197504 146424 214656 146452
rect 197504 146412 197510 146424
rect 214650 146412 214656 146424
rect 214708 146412 214714 146464
rect 224494 146412 224500 146464
rect 224552 146452 224558 146464
rect 241698 146452 241704 146464
rect 224552 146424 241704 146452
rect 224552 146412 224558 146424
rect 241698 146412 241704 146424
rect 241756 146412 241762 146464
rect 413462 146412 413468 146464
rect 413520 146452 413526 146464
rect 430666 146452 430672 146464
rect 413520 146424 430672 146452
rect 413520 146412 413526 146424
rect 430666 146412 430672 146424
rect 430724 146412 430730 146464
rect 440510 146412 440516 146464
rect 440568 146452 440574 146464
rect 457622 146452 457628 146464
rect 440568 146424 457628 146452
rect 440568 146412 440574 146424
rect 457622 146412 457628 146424
rect 457680 146412 457686 146464
rect 468478 146412 468484 146464
rect 468536 146452 468542 146464
rect 484670 146452 484676 146464
rect 468536 146424 484676 146452
rect 468536 146412 468542 146424
rect 484670 146412 484676 146424
rect 484728 146412 484734 146464
rect 36814 146344 36820 146396
rect 36872 146384 36878 146396
rect 62298 146384 62304 146396
rect 36872 146356 62304 146384
rect 36872 146344 36878 146356
rect 62298 146344 62304 146356
rect 62356 146344 62362 146396
rect 64138 146344 64144 146396
rect 64196 146384 64202 146396
rect 89346 146384 89352 146396
rect 64196 146356 89352 146384
rect 64196 146344 64202 146356
rect 89346 146344 89352 146356
rect 89404 146344 89410 146396
rect 90358 146344 90364 146396
rect 90416 146384 90422 146396
rect 116302 146384 116308 146396
rect 90416 146356 116308 146384
rect 90416 146344 90422 146356
rect 116302 146344 116308 146356
rect 116360 146344 116366 146396
rect 116578 146344 116584 146396
rect 116636 146384 116642 146396
rect 143350 146384 143356 146396
rect 116636 146356 143356 146384
rect 116636 146344 116642 146356
rect 143350 146344 143356 146356
rect 143408 146344 143414 146396
rect 144270 146344 144276 146396
rect 144328 146384 144334 146396
rect 170306 146384 170312 146396
rect 144328 146356 170312 146384
rect 144328 146344 144334 146356
rect 170306 146344 170312 146356
rect 170364 146344 170370 146396
rect 178034 146344 178040 146396
rect 178092 146384 178098 146396
rect 200758 146384 200764 146396
rect 178092 146356 200764 146384
rect 178092 146344 178098 146356
rect 200758 146344 200764 146356
rect 200816 146344 200822 146396
rect 251450 146344 251456 146396
rect 251508 146384 251514 146396
rect 268654 146384 268660 146396
rect 251508 146356 268660 146384
rect 251508 146344 251514 146356
rect 268654 146344 268660 146356
rect 268712 146344 268718 146396
rect 279510 146344 279516 146396
rect 279568 146384 279574 146396
rect 295702 146384 295708 146396
rect 279568 146356 295708 146384
rect 279568 146344 279574 146356
rect 295702 146344 295708 146356
rect 295760 146344 295766 146396
rect 305454 146344 305460 146396
rect 305512 146384 305518 146396
rect 322658 146384 322664 146396
rect 305512 146356 322664 146384
rect 305512 146344 305518 146356
rect 322658 146344 322664 146356
rect 322716 146344 322722 146396
rect 335998 146344 336004 146396
rect 336056 146384 336062 146396
rect 349706 146384 349712 146396
rect 336056 146356 349712 146384
rect 336056 146344 336062 146356
rect 349706 146344 349712 146356
rect 349764 146344 349770 146396
rect 359458 146344 359464 146396
rect 359516 146384 359522 146396
rect 376662 146384 376668 146396
rect 359516 146356 376668 146384
rect 359516 146344 359522 146356
rect 376662 146344 376668 146356
rect 376720 146344 376726 146396
rect 386506 146344 386512 146396
rect 386564 146384 386570 146396
rect 403618 146384 403624 146396
rect 386564 146356 403624 146384
rect 386564 146344 386570 146356
rect 403618 146344 403624 146356
rect 403676 146344 403682 146396
rect 421006 146344 421012 146396
rect 421064 146384 421070 146396
rect 445018 146384 445024 146396
rect 421064 146356 445024 146384
rect 421064 146344 421070 146356
rect 445018 146344 445024 146356
rect 445076 146344 445082 146396
rect 494514 146344 494520 146396
rect 494572 146384 494578 146396
rect 511626 146384 511632 146396
rect 494572 146356 511632 146384
rect 494572 146344 494578 146356
rect 511626 146344 511632 146356
rect 511684 146344 511690 146396
rect 522390 146344 522396 146396
rect 522448 146384 522454 146396
rect 538674 146384 538680 146396
rect 522448 146356 538680 146384
rect 522448 146344 522454 146356
rect 538674 146344 538680 146356
rect 538732 146344 538738 146396
rect 43070 146276 43076 146328
rect 43128 146316 43134 146328
rect 62758 146316 62764 146328
rect 43128 146288 62764 146316
rect 43128 146276 43134 146288
rect 62758 146276 62764 146288
rect 62816 146276 62822 146328
rect 171778 146276 171784 146328
rect 171836 146316 171842 146328
rect 197354 146316 197360 146328
rect 171836 146288 197360 146316
rect 171836 146276 171842 146288
rect 197354 146276 197360 146288
rect 197412 146276 197418 146328
rect 199378 146276 199384 146328
rect 199436 146316 199442 146328
rect 224310 146316 224316 146328
rect 199436 146288 224316 146316
rect 199436 146276 199442 146288
rect 224310 146276 224316 146288
rect 224368 146276 224374 146328
rect 225598 146276 225604 146328
rect 225656 146316 225662 146328
rect 251358 146316 251364 146328
rect 225656 146288 251364 146316
rect 225656 146276 225662 146288
rect 251358 146276 251364 146288
rect 251416 146276 251422 146328
rect 253198 146276 253204 146328
rect 253256 146316 253262 146328
rect 278314 146316 278320 146328
rect 253256 146288 278320 146316
rect 253256 146276 253262 146288
rect 278314 146276 278320 146288
rect 278372 146276 278378 146328
rect 279418 146276 279424 146328
rect 279476 146316 279482 146328
rect 305362 146316 305368 146328
rect 279476 146288 305368 146316
rect 279476 146276 279482 146288
rect 305362 146276 305368 146288
rect 305420 146276 305426 146328
rect 307018 146276 307024 146328
rect 307076 146316 307082 146328
rect 332318 146316 332324 146328
rect 307076 146288 332324 146316
rect 307076 146276 307082 146288
rect 332318 146276 332324 146288
rect 332376 146276 332382 146328
rect 333238 146276 333244 146328
rect 333296 146316 333302 146328
rect 359366 146316 359372 146328
rect 333296 146288 359372 146316
rect 333296 146276 333302 146288
rect 359366 146276 359372 146288
rect 359424 146276 359430 146328
rect 359550 146276 359556 146328
rect 359608 146316 359614 146328
rect 386322 146316 386328 146328
rect 359608 146288 386328 146316
rect 359608 146276 359614 146288
rect 386322 146276 386328 146288
rect 386380 146276 386386 146328
rect 387058 146276 387064 146328
rect 387116 146316 387122 146328
rect 413278 146316 413284 146328
rect 387116 146288 413284 146316
rect 387116 146276 387122 146288
rect 413278 146276 413284 146288
rect 413336 146276 413342 146328
rect 414658 146276 414664 146328
rect 414716 146316 414722 146328
rect 440326 146316 440332 146328
rect 414716 146288 440332 146316
rect 414716 146276 414722 146288
rect 440326 146276 440332 146288
rect 440384 146276 440390 146328
rect 442258 146276 442264 146328
rect 442316 146316 442322 146328
rect 467282 146316 467288 146328
rect 442316 146288 467288 146316
rect 442316 146276 442322 146288
rect 467282 146276 467288 146288
rect 467340 146276 467346 146328
rect 468570 146276 468576 146328
rect 468628 146316 468634 146328
rect 494330 146316 494336 146328
rect 468628 146288 494336 146316
rect 468628 146276 468634 146288
rect 494330 146276 494336 146288
rect 494388 146276 494394 146328
rect 496078 146276 496084 146328
rect 496136 146316 496142 146328
rect 521286 146316 521292 146328
rect 496136 146288 521292 146316
rect 496136 146276 496142 146288
rect 521286 146276 521292 146288
rect 521344 146276 521350 146328
rect 522298 146276 522304 146328
rect 522356 146316 522362 146328
rect 548334 146316 548340 146328
rect 522356 146288 548340 146316
rect 522356 146276 522362 146288
rect 548334 146276 548340 146288
rect 548392 146276 548398 146328
rect 37918 144168 37924 144220
rect 37976 144208 37982 144220
rect 526438 144208 526444 144220
rect 37976 144180 526444 144208
rect 37976 144168 37982 144180
rect 526438 144168 526444 144180
rect 526496 144168 526502 144220
rect 89714 128256 89720 128308
rect 89772 128296 89778 128308
rect 90450 128296 90456 128308
rect 89772 128268 90456 128296
rect 89772 128256 89778 128268
rect 90450 128256 90456 128268
rect 90508 128256 90514 128308
rect 13722 125536 13728 125588
rect 13780 125576 13786 125588
rect 64874 125576 64880 125588
rect 13780 125548 64880 125576
rect 13780 125536 13786 125548
rect 64874 125536 64880 125548
rect 64932 125536 64938 125588
rect 95142 125536 95148 125588
rect 95200 125576 95206 125588
rect 146294 125576 146300 125588
rect 95200 125548 146300 125576
rect 95200 125536 95206 125548
rect 146294 125536 146300 125548
rect 146352 125536 146358 125588
rect 148962 125536 148968 125588
rect 149020 125576 149026 125588
rect 200114 125576 200120 125588
rect 149020 125548 200120 125576
rect 149020 125536 149026 125548
rect 200114 125536 200120 125548
rect 200172 125536 200178 125588
rect 202782 125536 202788 125588
rect 202840 125576 202846 125588
rect 253934 125576 253940 125588
rect 202840 125548 253940 125576
rect 202840 125536 202846 125548
rect 253934 125536 253940 125548
rect 253992 125536 253998 125588
rect 256602 125536 256608 125588
rect 256660 125576 256666 125588
rect 307754 125576 307760 125588
rect 256660 125548 307760 125576
rect 256660 125536 256666 125548
rect 307754 125536 307760 125548
rect 307812 125536 307818 125588
rect 338022 125536 338028 125588
rect 338080 125576 338086 125588
rect 389174 125576 389180 125588
rect 338080 125548 389180 125576
rect 338080 125536 338086 125548
rect 389174 125536 389180 125548
rect 389232 125536 389238 125588
rect 391842 125536 391848 125588
rect 391900 125576 391906 125588
rect 442994 125576 443000 125588
rect 391900 125548 443000 125576
rect 391900 125536 391906 125548
rect 442994 125536 443000 125548
rect 443052 125536 443058 125588
rect 445662 125536 445668 125588
rect 445720 125576 445726 125588
rect 496814 125576 496820 125588
rect 445720 125548 496820 125576
rect 445720 125536 445726 125548
rect 496814 125536 496820 125548
rect 496872 125536 496878 125588
rect 500862 125536 500868 125588
rect 500920 125576 500926 125588
rect 550634 125576 550640 125588
rect 500920 125548 550640 125576
rect 500920 125536 500926 125548
rect 550634 125536 550640 125548
rect 550692 125536 550698 125588
rect 41322 125468 41328 125520
rect 41380 125508 41386 125520
rect 91094 125508 91100 125520
rect 41380 125480 91100 125508
rect 41380 125468 41386 125480
rect 91094 125468 91100 125480
rect 91152 125468 91158 125520
rect 122742 125468 122748 125520
rect 122800 125508 122806 125520
rect 172514 125508 172520 125520
rect 122800 125480 172520 125508
rect 122800 125468 122806 125480
rect 172514 125468 172520 125480
rect 172572 125468 172578 125520
rect 176562 125468 176568 125520
rect 176620 125508 176626 125520
rect 226334 125508 226340 125520
rect 176620 125480 226340 125508
rect 176620 125468 176626 125480
rect 226334 125468 226340 125480
rect 226392 125468 226398 125520
rect 230382 125468 230388 125520
rect 230440 125508 230446 125520
rect 230440 125480 277394 125508
rect 230440 125468 230446 125480
rect 68922 125400 68928 125452
rect 68980 125440 68986 125452
rect 118694 125440 118700 125452
rect 68980 125412 118700 125440
rect 68980 125400 68986 125412
rect 118694 125400 118700 125412
rect 118752 125400 118758 125452
rect 277366 125440 277394 125480
rect 278682 125468 278688 125520
rect 278740 125508 278746 125520
rect 279510 125508 279516 125520
rect 278740 125480 279516 125508
rect 278740 125468 278746 125480
rect 279510 125468 279516 125480
rect 279568 125468 279574 125520
rect 284202 125468 284208 125520
rect 284260 125508 284266 125520
rect 335354 125508 335360 125520
rect 284260 125480 335360 125508
rect 284260 125468 284266 125480
rect 335354 125468 335360 125480
rect 335412 125468 335418 125520
rect 365622 125468 365628 125520
rect 365680 125508 365686 125520
rect 415394 125508 415400 125520
rect 365680 125480 415400 125508
rect 365680 125468 365686 125480
rect 415394 125468 415400 125480
rect 415452 125468 415458 125520
rect 419442 125468 419448 125520
rect 419500 125508 419506 125520
rect 469214 125508 469220 125520
rect 419500 125480 469220 125508
rect 419500 125468 419506 125480
rect 469214 125468 469220 125480
rect 469272 125468 469278 125520
rect 473262 125468 473268 125520
rect 473320 125508 473326 125520
rect 523034 125508 523040 125520
rect 473320 125480 523040 125508
rect 473320 125468 473326 125480
rect 523034 125468 523040 125480
rect 523092 125468 523098 125520
rect 280154 125440 280160 125452
rect 277366 125412 280160 125440
rect 280154 125400 280160 125412
rect 280212 125400 280218 125452
rect 311802 125400 311808 125452
rect 311860 125440 311866 125452
rect 361574 125440 361580 125452
rect 311860 125412 361580 125440
rect 311860 125400 311866 125412
rect 361574 125400 361580 125412
rect 361632 125400 361638 125452
rect 445018 125400 445024 125452
rect 445076 125440 445082 125452
rect 447686 125440 447692 125452
rect 445076 125412 447692 125440
rect 445076 125400 445082 125412
rect 447686 125400 447692 125412
rect 447744 125400 447750 125452
rect 35618 124788 35624 124840
rect 35676 124828 35682 124840
rect 36722 124828 36728 124840
rect 35676 124800 36728 124828
rect 35676 124788 35682 124800
rect 36722 124788 36728 124800
rect 36780 124788 36786 124840
rect 116210 124584 116216 124636
rect 116268 124624 116274 124636
rect 116486 124624 116492 124636
rect 116268 124596 116492 124624
rect 116268 124584 116274 124596
rect 116486 124584 116492 124596
rect 116544 124584 116550 124636
rect 170214 124584 170220 124636
rect 170272 124624 170278 124636
rect 170490 124624 170496 124636
rect 170272 124596 170496 124624
rect 170272 124584 170278 124596
rect 170490 124584 170496 124596
rect 170548 124584 170554 124636
rect 62758 122748 62764 122800
rect 62816 122788 62822 122800
rect 69750 122788 69756 122800
rect 62816 122760 69756 122788
rect 62816 122748 62822 122760
rect 69750 122748 69756 122760
rect 69808 122748 69814 122800
rect 96614 122748 96620 122800
rect 96672 122788 96678 122800
rect 96672 122760 103514 122788
rect 96672 122748 96678 122760
rect 15194 122680 15200 122732
rect 15252 122720 15258 122732
rect 42794 122720 42800 122732
rect 15252 122692 42800 122720
rect 15252 122680 15258 122692
rect 42794 122680 42800 122692
rect 42852 122680 42858 122732
rect 53098 122680 53104 122732
rect 53156 122720 53162 122732
rect 64138 122720 64144 122732
rect 53156 122692 64144 122720
rect 53156 122680 53162 122692
rect 64138 122680 64144 122692
rect 64196 122680 64202 122732
rect 69106 122680 69112 122732
rect 69164 122720 69170 122732
rect 96706 122720 96712 122732
rect 69164 122692 96712 122720
rect 69164 122680 69170 122692
rect 96706 122680 96712 122692
rect 96764 122680 96770 122732
rect 103486 122720 103514 122760
rect 200758 122748 200764 122800
rect 200816 122788 200822 122800
rect 204622 122788 204628 122800
rect 200816 122760 204628 122788
rect 200816 122748 200822 122760
rect 204622 122748 204628 122760
rect 204680 122748 204686 122800
rect 251818 122748 251824 122800
rect 251876 122788 251882 122800
rect 258718 122788 258724 122800
rect 251876 122760 258724 122788
rect 251876 122748 251882 122760
rect 258718 122748 258724 122760
rect 258776 122748 258782 122800
rect 332502 122748 332508 122800
rect 332560 122788 332566 122800
rect 335998 122788 336004 122800
rect 332560 122760 336004 122788
rect 332560 122748 332566 122760
rect 335998 122748 336004 122760
rect 336056 122748 336062 122800
rect 494698 122748 494704 122800
rect 494756 122788 494762 122800
rect 501598 122788 501604 122800
rect 494756 122760 501604 122788
rect 494756 122748 494762 122760
rect 501598 122748 501604 122760
rect 501656 122748 501662 122800
rect 521470 122748 521476 122800
rect 521528 122788 521534 122800
rect 522390 122788 522396 122800
rect 521528 122760 522396 122788
rect 521528 122748 521534 122760
rect 522390 122748 522396 122760
rect 522448 122748 522454 122800
rect 123662 122720 123668 122732
rect 103486 122692 123668 122720
rect 123662 122680 123668 122692
rect 123720 122680 123726 122732
rect 133782 122680 133788 122732
rect 133840 122720 133846 122732
rect 144270 122720 144276 122732
rect 133840 122692 144276 122720
rect 133840 122680 133846 122692
rect 144270 122680 144276 122692
rect 144328 122680 144334 122732
rect 146938 122680 146944 122732
rect 146996 122720 147002 122732
rect 547966 122720 547972 122732
rect 146996 122692 547972 122720
rect 146996 122680 147002 122692
rect 547966 122680 547972 122692
rect 548024 122680 548030 122732
rect 26050 122612 26056 122664
rect 26108 122652 26114 122664
rect 36814 122652 36820 122664
rect 26108 122624 36820 122652
rect 26108 122612 26114 122624
rect 36814 122612 36820 122624
rect 36872 122612 36878 122664
rect 79962 122612 79968 122664
rect 80020 122652 80026 122664
rect 90358 122652 90364 122664
rect 80020 122624 90364 122652
rect 80020 122612 80026 122624
rect 90358 122612 90364 122624
rect 90416 122612 90422 122664
rect 106550 122612 106556 122664
rect 106608 122652 106614 122664
rect 116578 122652 116584 122664
rect 106608 122624 116584 122652
rect 106608 122612 106614 122624
rect 116578 122612 116584 122624
rect 116636 122612 116642 122664
rect 122926 122612 122932 122664
rect 122984 122652 122990 122664
rect 122984 122624 142154 122652
rect 122984 122612 122990 122624
rect 142126 122584 142154 122624
rect 150526 122612 150532 122664
rect 150584 122652 150590 122664
rect 178126 122652 178132 122664
rect 150584 122624 178132 122652
rect 150584 122612 150590 122624
rect 178126 122612 178132 122624
rect 178184 122612 178190 122664
rect 187970 122612 187976 122664
rect 188028 122652 188034 122664
rect 199378 122652 199384 122664
rect 188028 122624 199384 122652
rect 188028 122612 188034 122624
rect 199378 122612 199384 122624
rect 199436 122612 199442 122664
rect 204346 122612 204352 122664
rect 204404 122652 204410 122664
rect 231946 122652 231952 122664
rect 204404 122624 231952 122652
rect 204404 122612 204410 122624
rect 231946 122612 231952 122624
rect 232004 122612 232010 122664
rect 242066 122612 242072 122664
rect 242124 122652 242130 122664
rect 253198 122652 253204 122664
rect 242124 122624 253204 122652
rect 242124 122612 242130 122624
rect 253198 122612 253204 122624
rect 253256 122612 253262 122664
rect 258166 122612 258172 122664
rect 258224 122652 258230 122664
rect 258224 122624 281764 122652
rect 258224 122612 258230 122624
rect 150710 122584 150716 122596
rect 142126 122556 150716 122584
rect 150710 122544 150716 122556
rect 150768 122544 150774 122596
rect 160554 122544 160560 122596
rect 160612 122584 160618 122596
rect 171778 122584 171784 122596
rect 160612 122556 171784 122584
rect 160612 122544 160618 122556
rect 171778 122544 171784 122556
rect 171836 122544 171842 122596
rect 215018 122544 215024 122596
rect 215076 122584 215082 122596
rect 225598 122584 225604 122596
rect 215076 122556 225604 122584
rect 215076 122544 215082 122556
rect 225598 122544 225604 122556
rect 225656 122544 225662 122596
rect 268930 122544 268936 122596
rect 268988 122584 268994 122596
rect 279418 122584 279424 122596
rect 268988 122556 279424 122584
rect 268988 122544 268994 122556
rect 279418 122544 279424 122556
rect 279476 122544 279482 122596
rect 281736 122584 281764 122624
rect 285766 122612 285772 122664
rect 285824 122652 285830 122664
rect 312630 122652 312636 122664
rect 285824 122624 312636 122652
rect 285824 122612 285830 122624
rect 312630 122612 312636 122624
rect 312688 122612 312694 122664
rect 316006 122624 335354 122652
rect 286134 122584 286140 122596
rect 281736 122556 286140 122584
rect 286134 122544 286140 122556
rect 286192 122544 286198 122596
rect 295978 122544 295984 122596
rect 296036 122584 296042 122596
rect 307018 122584 307024 122596
rect 296036 122556 307024 122584
rect 296036 122544 296042 122556
rect 307018 122544 307024 122556
rect 307076 122544 307082 122596
rect 311986 122544 311992 122596
rect 312044 122584 312050 122596
rect 316006 122584 316034 122624
rect 312044 122556 316034 122584
rect 312044 122544 312050 122556
rect 322842 122544 322848 122596
rect 322900 122584 322906 122596
rect 333238 122584 333244 122596
rect 322900 122556 333244 122584
rect 322900 122544 322906 122556
rect 333238 122544 333244 122556
rect 333296 122544 333302 122596
rect 335326 122584 335354 122624
rect 339586 122612 339592 122664
rect 339644 122652 339650 122664
rect 366726 122652 366732 122664
rect 339644 122624 366732 122652
rect 339644 122612 339650 122624
rect 366726 122612 366732 122624
rect 366784 122612 366790 122664
rect 393590 122652 393596 122664
rect 373966 122624 393596 122652
rect 340138 122584 340144 122596
rect 335326 122556 340144 122584
rect 340138 122544 340144 122556
rect 340196 122544 340202 122596
rect 350074 122544 350080 122596
rect 350132 122584 350138 122596
rect 359550 122584 359556 122596
rect 350132 122556 359556 122584
rect 350132 122544 350138 122556
rect 359550 122544 359556 122556
rect 359608 122544 359614 122596
rect 365806 122544 365812 122596
rect 365864 122584 365870 122596
rect 373966 122584 373994 122624
rect 393590 122612 393596 122624
rect 393648 122612 393654 122664
rect 420914 122652 420920 122664
rect 402946 122624 420920 122652
rect 365864 122556 373994 122584
rect 365864 122544 365870 122556
rect 376570 122544 376576 122596
rect 376628 122584 376634 122596
rect 387058 122584 387064 122596
rect 376628 122556 387064 122584
rect 376628 122544 376634 122556
rect 387058 122544 387064 122556
rect 387116 122544 387122 122596
rect 393406 122544 393412 122596
rect 393464 122584 393470 122596
rect 402946 122584 402974 122624
rect 420914 122612 420920 122624
rect 420972 122612 420978 122664
rect 431034 122612 431040 122664
rect 431092 122652 431098 122664
rect 442258 122652 442264 122664
rect 431092 122624 442264 122652
rect 431092 122612 431098 122624
rect 442258 122612 442264 122624
rect 442316 122612 442322 122664
rect 447226 122612 447232 122664
rect 447284 122652 447290 122664
rect 474734 122652 474740 122664
rect 447284 122624 474740 122652
rect 447284 122612 447290 122624
rect 474734 122612 474740 122624
rect 474792 122612 474798 122664
rect 484946 122612 484952 122664
rect 485004 122652 485010 122664
rect 496078 122652 496084 122664
rect 485004 122624 496084 122652
rect 485004 122612 485010 122624
rect 496078 122612 496084 122624
rect 496136 122612 496142 122664
rect 501046 122612 501052 122664
rect 501104 122652 501110 122664
rect 528646 122652 528652 122664
rect 501104 122624 528652 122652
rect 501104 122612 501110 122624
rect 528646 122612 528652 122624
rect 528704 122612 528710 122664
rect 393464 122556 402974 122584
rect 393464 122544 393470 122556
rect 403986 122544 403992 122596
rect 404044 122584 404050 122596
rect 414658 122584 414664 122596
rect 404044 122556 414664 122584
rect 404044 122544 404050 122556
rect 414658 122544 414664 122556
rect 414716 122544 414722 122596
rect 458082 122544 458088 122596
rect 458140 122584 458146 122596
rect 468570 122584 468576 122596
rect 458140 122556 468576 122584
rect 458140 122544 458146 122556
rect 468570 122544 468576 122556
rect 468628 122544 468634 122596
rect 511810 122544 511816 122596
rect 511868 122584 511874 122596
rect 522298 122584 522304 122596
rect 511868 122556 522304 122584
rect 511868 122544 511874 122556
rect 522298 122544 522304 122556
rect 522356 122544 522362 122596
rect 36630 122476 36636 122528
rect 36688 122516 36694 122528
rect 538398 122516 538404 122528
rect 36688 122488 538404 122516
rect 36688 122476 36694 122488
rect 538398 122476 538404 122488
rect 538456 122476 538462 122528
rect 16298 119348 16304 119400
rect 16356 119388 16362 119400
rect 528738 119388 528744 119400
rect 16356 119360 528744 119388
rect 16356 119348 16362 119360
rect 528738 119348 528744 119360
rect 528796 119348 528802 119400
rect 25958 118940 25964 118992
rect 26016 118980 26022 118992
rect 146938 118980 146944 118992
rect 26016 118952 146944 118980
rect 26016 118940 26022 118952
rect 146938 118940 146944 118952
rect 146996 118940 147002 118992
rect 36814 118872 36820 118924
rect 36872 118912 36878 118924
rect 52454 118912 52460 118924
rect 36872 118884 52460 118912
rect 36872 118872 36878 118884
rect 52454 118872 52460 118884
rect 52512 118872 52518 118924
rect 232314 118872 232320 118924
rect 232372 118912 232378 118924
rect 251818 118912 251824 118924
rect 232372 118884 251824 118912
rect 232372 118872 232378 118884
rect 251818 118872 251824 118884
rect 251876 118872 251882 118924
rect 62482 118804 62488 118856
rect 62540 118844 62546 118856
rect 79318 118844 79324 118856
rect 62540 118816 79324 118844
rect 62540 118804 62546 118816
rect 79318 118804 79324 118816
rect 79376 118804 79382 118856
rect 90450 118804 90456 118856
rect 90508 118844 90514 118856
rect 106366 118844 106372 118856
rect 90508 118816 106372 118844
rect 90508 118804 90514 118816
rect 106366 118804 106372 118816
rect 106424 118804 106430 118856
rect 116486 118804 116492 118856
rect 116544 118844 116550 118856
rect 133414 118844 133420 118856
rect 116544 118816 133420 118844
rect 116544 118804 116550 118816
rect 133414 118804 133420 118816
rect 133472 118804 133478 118856
rect 170490 118804 170496 118856
rect 170548 118844 170554 118856
rect 187786 118844 187792 118856
rect 170548 118816 187792 118844
rect 170548 118804 170554 118816
rect 187786 118804 187792 118816
rect 187844 118804 187850 118856
rect 197538 118804 197544 118856
rect 197596 118844 197602 118856
rect 214374 118844 214380 118856
rect 197596 118816 214380 118844
rect 197596 118804 197602 118816
rect 214374 118804 214380 118816
rect 214432 118804 214438 118856
rect 224494 118804 224500 118856
rect 224552 118844 224558 118856
rect 241514 118844 241520 118856
rect 224552 118816 241520 118844
rect 224552 118804 224558 118816
rect 241514 118804 241520 118816
rect 241572 118804 241578 118856
rect 413462 118804 413468 118856
rect 413520 118844 413526 118856
rect 430574 118844 430580 118856
rect 413520 118816 430580 118844
rect 413520 118804 413526 118816
rect 430574 118804 430580 118816
rect 430632 118804 430638 118856
rect 440510 118804 440516 118856
rect 440568 118844 440574 118856
rect 457254 118844 457260 118856
rect 440568 118816 457260 118844
rect 440568 118804 440574 118816
rect 457254 118804 457260 118816
rect 457312 118804 457318 118856
rect 468570 118804 468576 118856
rect 468628 118844 468634 118856
rect 484394 118844 484400 118856
rect 468628 118816 484400 118844
rect 468628 118804 468634 118816
rect 484394 118804 484400 118816
rect 484452 118804 484458 118856
rect 494514 118804 494520 118856
rect 494572 118844 494578 118856
rect 511350 118844 511356 118856
rect 494572 118816 511356 118844
rect 494572 118804 494578 118816
rect 511350 118804 511356 118816
rect 511408 118804 511414 118856
rect 36630 118736 36636 118788
rect 36688 118776 36694 118788
rect 62114 118776 62120 118788
rect 36688 118748 62120 118776
rect 36688 118736 36694 118748
rect 62114 118736 62120 118748
rect 62172 118736 62178 118788
rect 64138 118736 64144 118788
rect 64196 118776 64202 118788
rect 89070 118776 89076 118788
rect 64196 118748 89076 118776
rect 64196 118736 64202 118748
rect 89070 118736 89076 118748
rect 89128 118736 89134 118788
rect 90358 118736 90364 118788
rect 90416 118776 90422 118788
rect 115934 118776 115940 118788
rect 90416 118748 115940 118776
rect 90416 118736 90422 118748
rect 115934 118736 115940 118748
rect 115992 118736 115998 118788
rect 116578 118736 116584 118788
rect 116636 118776 116642 118788
rect 142982 118776 142988 118788
rect 116636 118748 142988 118776
rect 116636 118736 116642 118748
rect 142982 118736 142988 118748
rect 143040 118736 143046 118788
rect 144178 118736 144184 118788
rect 144236 118776 144242 118788
rect 170030 118776 170036 118788
rect 144236 118748 170036 118776
rect 144236 118736 144242 118748
rect 170030 118736 170036 118748
rect 170088 118736 170094 118788
rect 178402 118736 178408 118788
rect 178460 118776 178466 118788
rect 200758 118776 200764 118788
rect 178460 118748 200764 118776
rect 178460 118736 178466 118748
rect 200758 118736 200764 118748
rect 200816 118736 200822 118788
rect 251450 118736 251456 118788
rect 251508 118776 251514 118788
rect 268286 118776 268292 118788
rect 251508 118748 268292 118776
rect 251508 118736 251514 118748
rect 268286 118736 268292 118748
rect 268344 118736 268350 118788
rect 279418 118736 279424 118788
rect 279476 118776 279482 118788
rect 295794 118776 295800 118788
rect 279476 118748 295800 118776
rect 279476 118736 279482 118748
rect 295794 118736 295800 118748
rect 295852 118736 295858 118788
rect 305638 118736 305644 118788
rect 305696 118776 305702 118788
rect 322382 118776 322388 118788
rect 305696 118748 322388 118776
rect 305696 118736 305702 118748
rect 322382 118736 322388 118748
rect 322440 118736 322446 118788
rect 334618 118736 334624 118788
rect 334676 118776 334682 118788
rect 349798 118776 349804 118788
rect 334676 118748 349804 118776
rect 334676 118736 334682 118748
rect 349798 118736 349804 118748
rect 349856 118736 349862 118788
rect 359550 118736 359556 118788
rect 359608 118776 359614 118788
rect 376294 118776 376300 118788
rect 359608 118748 376300 118776
rect 359608 118736 359614 118748
rect 376294 118736 376300 118748
rect 376352 118736 376358 118788
rect 386506 118736 386512 118788
rect 386564 118776 386570 118788
rect 403342 118776 403348 118788
rect 386564 118748 403348 118776
rect 386564 118736 386570 118748
rect 403342 118736 403348 118748
rect 403400 118736 403406 118788
rect 421282 118736 421288 118788
rect 421340 118776 421346 118788
rect 443638 118776 443644 118788
rect 421340 118748 443644 118776
rect 421340 118736 421346 118748
rect 443638 118736 443644 118748
rect 443696 118736 443702 118788
rect 475378 118736 475384 118788
rect 475436 118776 475442 118788
rect 494698 118776 494704 118788
rect 475436 118748 494704 118776
rect 475436 118736 475442 118748
rect 494698 118736 494704 118748
rect 494756 118736 494762 118788
rect 522390 118736 522396 118788
rect 522448 118776 522454 118788
rect 538398 118776 538404 118788
rect 522448 118748 538404 118776
rect 522448 118736 522454 118748
rect 538398 118736 538404 118748
rect 538456 118736 538462 118788
rect 43346 118668 43352 118720
rect 43404 118708 43410 118720
rect 62758 118708 62764 118720
rect 43404 118680 62764 118708
rect 43404 118668 43410 118680
rect 62758 118668 62764 118680
rect 62816 118668 62822 118720
rect 144270 118668 144276 118720
rect 144328 118708 144334 118720
rect 160278 118708 160284 118720
rect 144328 118680 160284 118708
rect 144328 118668 144334 118680
rect 160278 118668 160284 118680
rect 160336 118668 160342 118720
rect 171778 118668 171784 118720
rect 171836 118708 171842 118720
rect 197446 118708 197452 118720
rect 171836 118680 197452 118708
rect 171836 118668 171842 118680
rect 197446 118668 197452 118680
rect 197504 118668 197510 118720
rect 199378 118668 199384 118720
rect 199436 118708 199442 118720
rect 223942 118708 223948 118720
rect 199436 118680 223948 118708
rect 199436 118668 199442 118680
rect 223942 118668 223948 118680
rect 224000 118668 224006 118720
rect 225598 118668 225604 118720
rect 225656 118708 225662 118720
rect 251174 118708 251180 118720
rect 225656 118680 251180 118708
rect 225656 118668 225662 118680
rect 251174 118668 251180 118680
rect 251232 118668 251238 118720
rect 253198 118668 253204 118720
rect 253256 118708 253262 118720
rect 278038 118708 278044 118720
rect 253256 118680 278044 118708
rect 253256 118668 253262 118680
rect 278038 118668 278044 118680
rect 278096 118668 278102 118720
rect 279510 118668 279516 118720
rect 279568 118708 279574 118720
rect 305546 118708 305552 118720
rect 279568 118680 305552 118708
rect 279568 118668 279574 118680
rect 305546 118668 305552 118680
rect 305604 118668 305610 118720
rect 307018 118668 307024 118720
rect 307076 118708 307082 118720
rect 331950 118708 331956 118720
rect 307076 118680 331956 118708
rect 307076 118668 307082 118680
rect 331950 118668 331956 118680
rect 332008 118668 332014 118720
rect 333238 118668 333244 118720
rect 333296 118708 333302 118720
rect 359458 118708 359464 118720
rect 333296 118680 359464 118708
rect 333296 118668 333302 118680
rect 359458 118668 359464 118680
rect 359516 118668 359522 118720
rect 359734 118668 359740 118720
rect 359792 118708 359798 118720
rect 386046 118708 386052 118720
rect 359792 118680 386052 118708
rect 359792 118668 359798 118680
rect 386046 118668 386052 118680
rect 386104 118668 386110 118720
rect 387058 118668 387064 118720
rect 387116 118708 387122 118720
rect 412910 118708 412916 118720
rect 387116 118680 412916 118708
rect 387116 118668 387122 118680
rect 412910 118668 412916 118680
rect 412968 118668 412974 118720
rect 414658 118668 414664 118720
rect 414716 118708 414722 118720
rect 440234 118708 440240 118720
rect 414716 118680 440240 118708
rect 414716 118668 414722 118680
rect 440234 118668 440240 118680
rect 440292 118668 440298 118720
rect 442258 118668 442264 118720
rect 442316 118708 442322 118720
rect 467006 118708 467012 118720
rect 442316 118680 467012 118708
rect 442316 118668 442322 118680
rect 467006 118668 467012 118680
rect 467064 118668 467070 118720
rect 468478 118668 468484 118720
rect 468536 118708 468542 118720
rect 494054 118708 494060 118720
rect 468536 118680 494060 118708
rect 468536 118668 468542 118680
rect 494054 118668 494060 118680
rect 494112 118668 494118 118720
rect 496078 118668 496084 118720
rect 496136 118708 496142 118720
rect 520918 118708 520924 118720
rect 496136 118680 520924 118708
rect 496136 118668 496142 118680
rect 520918 118668 520924 118680
rect 520976 118668 520982 118720
rect 522298 118668 522304 118720
rect 522356 118708 522362 118720
rect 548058 118708 548064 118720
rect 522356 118680 548064 118708
rect 522356 118668 522362 118680
rect 548058 118668 548064 118680
rect 548116 118668 548122 118720
rect 37918 116560 37924 116612
rect 37976 116600 37982 116612
rect 526438 116600 526444 116612
rect 37976 116572 526444 116600
rect 37976 116560 37982 116572
rect 526438 116560 526444 116572
rect 526496 116560 526502 116612
rect 285766 116356 285772 116408
rect 285824 116396 285830 116408
rect 286134 116396 286140 116408
rect 285824 116368 286140 116396
rect 285824 116356 285830 116368
rect 286134 116356 286140 116368
rect 286192 116356 286198 116408
rect 339586 116288 339592 116340
rect 339644 116328 339650 116340
rect 340138 116328 340144 116340
rect 339644 116300 340144 116328
rect 339644 116288 339650 116300
rect 340138 116288 340144 116300
rect 340196 116288 340202 116340
rect 35618 116084 35624 116136
rect 35676 116124 35682 116136
rect 36722 116124 36728 116136
rect 35676 116096 36728 116124
rect 35676 116084 35682 116096
rect 36722 116084 36728 116096
rect 36780 116084 36786 116136
rect 89714 100240 89720 100292
rect 89772 100280 89778 100292
rect 90450 100280 90456 100292
rect 89772 100252 90456 100280
rect 89772 100240 89778 100252
rect 90450 100240 90456 100252
rect 90508 100240 90514 100292
rect 143626 100240 143632 100292
rect 143684 100280 143690 100292
rect 144270 100280 144276 100292
rect 143684 100252 144276 100280
rect 143684 100240 143690 100252
rect 144270 100240 144276 100252
rect 144328 100240 144334 100292
rect 521746 100240 521752 100292
rect 521804 100280 521810 100292
rect 522390 100280 522396 100292
rect 521804 100252 522396 100280
rect 521804 100240 521810 100252
rect 522390 100240 522396 100252
rect 522448 100240 522454 100292
rect 13722 97928 13728 97980
rect 13780 97968 13786 97980
rect 64874 97968 64880 97980
rect 13780 97940 64880 97968
rect 13780 97928 13786 97940
rect 64874 97928 64880 97940
rect 64932 97928 64938 97980
rect 95142 97928 95148 97980
rect 95200 97968 95206 97980
rect 146294 97968 146300 97980
rect 95200 97940 146300 97968
rect 95200 97928 95206 97940
rect 146294 97928 146300 97940
rect 146352 97928 146358 97980
rect 148962 97928 148968 97980
rect 149020 97968 149026 97980
rect 200114 97968 200120 97980
rect 149020 97940 200120 97968
rect 149020 97928 149026 97940
rect 200114 97928 200120 97940
rect 200172 97928 200178 97980
rect 202782 97928 202788 97980
rect 202840 97968 202846 97980
rect 253934 97968 253940 97980
rect 202840 97940 253940 97968
rect 202840 97928 202846 97940
rect 253934 97928 253940 97940
rect 253992 97928 253998 97980
rect 284202 97928 284208 97980
rect 284260 97968 284266 97980
rect 335354 97968 335360 97980
rect 284260 97940 335360 97968
rect 284260 97928 284266 97940
rect 335354 97928 335360 97940
rect 335412 97928 335418 97980
rect 338022 97928 338028 97980
rect 338080 97968 338086 97980
rect 389174 97968 389180 97980
rect 338080 97940 389180 97968
rect 338080 97928 338086 97940
rect 389174 97928 389180 97940
rect 389232 97928 389238 97980
rect 391842 97928 391848 97980
rect 391900 97968 391906 97980
rect 442994 97968 443000 97980
rect 391900 97940 443000 97968
rect 391900 97928 391906 97940
rect 442994 97928 443000 97940
rect 443052 97928 443058 97980
rect 445662 97928 445668 97980
rect 445720 97968 445726 97980
rect 496814 97968 496820 97980
rect 445720 97940 496820 97968
rect 445720 97928 445726 97940
rect 496814 97928 496820 97940
rect 496872 97928 496878 97980
rect 500862 97928 500868 97980
rect 500920 97968 500926 97980
rect 550634 97968 550640 97980
rect 500920 97940 550640 97968
rect 500920 97928 500926 97940
rect 550634 97928 550640 97940
rect 550692 97928 550698 97980
rect 41322 97860 41328 97912
rect 41380 97900 41386 97912
rect 91094 97900 91100 97912
rect 41380 97872 91100 97900
rect 41380 97860 41386 97872
rect 91094 97860 91100 97872
rect 91152 97860 91158 97912
rect 122742 97860 122748 97912
rect 122800 97900 122806 97912
rect 172514 97900 172520 97912
rect 122800 97872 172520 97900
rect 122800 97860 122806 97872
rect 172514 97860 172520 97872
rect 172572 97860 172578 97912
rect 176562 97860 176568 97912
rect 176620 97900 176626 97912
rect 226334 97900 226340 97912
rect 176620 97872 226340 97900
rect 176620 97860 176626 97872
rect 226334 97860 226340 97872
rect 226392 97860 226398 97912
rect 256602 97860 256608 97912
rect 256660 97900 256666 97912
rect 307754 97900 307760 97912
rect 256660 97872 307760 97900
rect 256660 97860 256666 97872
rect 307754 97860 307760 97872
rect 307812 97860 307818 97912
rect 311802 97860 311808 97912
rect 311860 97900 311866 97912
rect 361574 97900 361580 97912
rect 311860 97872 361580 97900
rect 311860 97860 311866 97872
rect 361574 97860 361580 97872
rect 361632 97860 361638 97912
rect 365622 97860 365628 97912
rect 365680 97900 365686 97912
rect 415394 97900 415400 97912
rect 365680 97872 415400 97900
rect 365680 97860 365686 97872
rect 415394 97860 415400 97872
rect 415452 97860 415458 97912
rect 419442 97860 419448 97912
rect 419500 97900 419506 97912
rect 469214 97900 469220 97912
rect 419500 97872 469220 97900
rect 419500 97860 419506 97872
rect 469214 97860 469220 97872
rect 469272 97860 469278 97912
rect 473262 97860 473268 97912
rect 473320 97900 473326 97912
rect 523034 97900 523040 97912
rect 473320 97872 523040 97900
rect 473320 97860 473326 97872
rect 523034 97860 523040 97872
rect 523092 97860 523098 97912
rect 68922 97792 68928 97844
rect 68980 97832 68986 97844
rect 118694 97832 118700 97844
rect 68980 97804 118700 97832
rect 68980 97792 68986 97804
rect 118694 97792 118700 97804
rect 118752 97792 118758 97844
rect 200758 97792 200764 97844
rect 200816 97832 200822 97844
rect 204622 97832 204628 97844
rect 200816 97804 204628 97832
rect 200816 97792 200822 97804
rect 204622 97792 204628 97804
rect 204680 97792 204686 97844
rect 230382 97792 230388 97844
rect 230440 97832 230446 97844
rect 280154 97832 280160 97844
rect 230440 97804 280160 97832
rect 230440 97792 230446 97804
rect 280154 97792 280160 97804
rect 280212 97792 280218 97844
rect 332502 97792 332508 97844
rect 332560 97832 332566 97844
rect 334618 97832 334624 97844
rect 332560 97804 334624 97832
rect 332560 97792 332566 97804
rect 334618 97792 334624 97804
rect 334676 97792 334682 97844
rect 443638 97792 443644 97844
rect 443696 97832 443702 97844
rect 447686 97832 447692 97844
rect 443696 97804 447692 97832
rect 443696 97792 443702 97804
rect 447686 97792 447692 97804
rect 447744 97792 447750 97844
rect 467650 97792 467656 97844
rect 467708 97832 467714 97844
rect 468570 97832 468576 97844
rect 467708 97804 468576 97832
rect 467708 97792 467714 97804
rect 468570 97792 468576 97804
rect 468628 97792 468634 97844
rect 35618 97656 35624 97708
rect 35676 97696 35682 97708
rect 36814 97696 36820 97708
rect 35676 97668 36820 97696
rect 35676 97656 35682 97668
rect 36814 97656 36820 97668
rect 36872 97656 36878 97708
rect 257982 96636 257988 96688
rect 258040 96676 258046 96688
rect 258718 96676 258724 96688
rect 258040 96648 258724 96676
rect 258040 96636 258046 96648
rect 258718 96636 258724 96648
rect 258776 96636 258782 96688
rect 494698 96636 494704 96688
rect 494756 96676 494762 96688
rect 501598 96676 501604 96688
rect 494756 96648 501604 96676
rect 494756 96636 494762 96648
rect 501598 96636 501604 96648
rect 501656 96636 501662 96688
rect 62758 95140 62764 95192
rect 62816 95180 62822 95192
rect 70026 95180 70032 95192
rect 62816 95152 70032 95180
rect 62816 95140 62822 95152
rect 70026 95140 70032 95152
rect 70084 95140 70090 95192
rect 96706 95140 96712 95192
rect 96764 95180 96770 95192
rect 96764 95152 103514 95180
rect 96764 95140 96770 95152
rect 15194 95072 15200 95124
rect 15252 95112 15258 95124
rect 42978 95112 42984 95124
rect 15252 95084 42984 95112
rect 15252 95072 15258 95084
rect 42978 95072 42984 95084
rect 43036 95072 43042 95124
rect 52730 95072 52736 95124
rect 52788 95112 52794 95124
rect 64138 95112 64144 95124
rect 52788 95084 64144 95112
rect 52788 95072 52794 95084
rect 64138 95072 64144 95084
rect 64196 95072 64202 95124
rect 69106 95072 69112 95124
rect 69164 95112 69170 95124
rect 96982 95112 96988 95124
rect 69164 95084 96988 95112
rect 69164 95072 69170 95084
rect 96982 95072 96988 95084
rect 97040 95072 97046 95124
rect 103486 95112 103514 95152
rect 251818 95140 251824 95192
rect 251876 95180 251882 95192
rect 257982 95180 257988 95192
rect 251876 95152 257988 95180
rect 251876 95140 251882 95152
rect 257982 95140 257988 95152
rect 258040 95140 258046 95192
rect 124030 95112 124036 95124
rect 103486 95084 124036 95112
rect 124030 95072 124036 95084
rect 124088 95072 124094 95124
rect 149698 95072 149704 95124
rect 149756 95112 149762 95124
rect 548334 95112 548340 95124
rect 149756 95084 548340 95112
rect 149756 95072 149762 95084
rect 548334 95072 548340 95084
rect 548392 95072 548398 95124
rect 25682 95004 25688 95056
rect 25740 95044 25746 95056
rect 36630 95044 36636 95056
rect 25740 95016 36636 95044
rect 25740 95004 25746 95016
rect 36630 95004 36636 95016
rect 36688 95004 36694 95056
rect 79686 95004 79692 95056
rect 79744 95044 79750 95056
rect 90358 95044 90364 95056
rect 79744 95016 90364 95044
rect 79744 95004 79750 95016
rect 90358 95004 90364 95016
rect 90416 95004 90422 95056
rect 106642 95004 106648 95056
rect 106700 95044 106706 95056
rect 116578 95044 116584 95056
rect 106700 95016 116584 95044
rect 106700 95004 106706 95016
rect 116578 95004 116584 95016
rect 116636 95004 116642 95056
rect 133690 95004 133696 95056
rect 133748 95044 133754 95056
rect 144178 95044 144184 95056
rect 133748 95016 144184 95044
rect 133748 95004 133754 95016
rect 144178 95004 144184 95016
rect 144236 95004 144242 95056
rect 150526 95004 150532 95056
rect 150584 95044 150590 95056
rect 178034 95044 178040 95056
rect 150584 95016 178040 95044
rect 150584 95004 150590 95016
rect 178034 95004 178040 95016
rect 178092 95004 178098 95056
rect 187694 95004 187700 95056
rect 187752 95044 187758 95056
rect 199378 95044 199384 95056
rect 187752 95016 199384 95044
rect 187752 95004 187758 95016
rect 199378 95004 199384 95016
rect 199436 95004 199442 95056
rect 204346 95004 204352 95056
rect 204404 95044 204410 95056
rect 232038 95044 232044 95056
rect 204404 95016 232044 95044
rect 204404 95004 204410 95016
rect 232038 95004 232044 95016
rect 232096 95004 232102 95056
rect 241698 95004 241704 95056
rect 241756 95044 241762 95056
rect 253198 95044 253204 95056
rect 241756 95016 253204 95044
rect 241756 95004 241762 95016
rect 253198 95004 253204 95016
rect 253256 95004 253262 95056
rect 258166 95004 258172 95056
rect 258224 95044 258230 95056
rect 286042 95044 286048 95056
rect 258224 95016 286048 95044
rect 258224 95004 258230 95016
rect 286042 95004 286048 95016
rect 286100 95004 286106 95056
rect 312998 95044 313004 95056
rect 287026 95016 313004 95044
rect 122926 94936 122932 94988
rect 122984 94976 122990 94988
rect 150986 94976 150992 94988
rect 122984 94948 150992 94976
rect 122984 94936 122990 94948
rect 150986 94936 150992 94948
rect 151044 94936 151050 94988
rect 160646 94936 160652 94988
rect 160704 94976 160710 94988
rect 171778 94976 171784 94988
rect 160704 94948 171784 94976
rect 160704 94936 160710 94948
rect 171778 94936 171784 94948
rect 171836 94936 171842 94988
rect 214650 94936 214656 94988
rect 214708 94976 214714 94988
rect 225598 94976 225604 94988
rect 214708 94948 225604 94976
rect 214708 94936 214714 94948
rect 225598 94936 225604 94948
rect 225656 94936 225662 94988
rect 268654 94936 268660 94988
rect 268712 94976 268718 94988
rect 279510 94976 279516 94988
rect 268712 94948 279516 94976
rect 268712 94936 268718 94948
rect 279510 94936 279516 94948
rect 279568 94936 279574 94988
rect 285766 94936 285772 94988
rect 285824 94976 285830 94988
rect 287026 94976 287054 95016
rect 312998 95004 313004 95016
rect 313056 95004 313062 95056
rect 340046 95044 340052 95056
rect 316006 95016 340052 95044
rect 285824 94948 287054 94976
rect 285824 94936 285830 94948
rect 295702 94936 295708 94988
rect 295760 94976 295766 94988
rect 307018 94976 307024 94988
rect 295760 94948 307024 94976
rect 295760 94936 295766 94948
rect 307018 94936 307024 94948
rect 307076 94936 307082 94988
rect 311986 94936 311992 94988
rect 312044 94976 312050 94988
rect 316006 94976 316034 95016
rect 340046 95004 340052 95016
rect 340104 95004 340110 95056
rect 367002 95044 367008 95056
rect 344986 95016 367008 95044
rect 312044 94948 316034 94976
rect 312044 94936 312050 94948
rect 322658 94936 322664 94988
rect 322716 94976 322722 94988
rect 333238 94976 333244 94988
rect 322716 94948 333244 94976
rect 322716 94936 322722 94948
rect 333238 94936 333244 94948
rect 333296 94936 333302 94988
rect 339586 94936 339592 94988
rect 339644 94976 339650 94988
rect 344986 94976 345014 95016
rect 367002 95004 367008 95016
rect 367060 95004 367066 95056
rect 393958 95044 393964 95056
rect 373966 95016 393964 95044
rect 339644 94948 345014 94976
rect 339644 94936 339650 94948
rect 349706 94936 349712 94988
rect 349764 94976 349770 94988
rect 359550 94976 359556 94988
rect 349764 94948 359556 94976
rect 349764 94936 349770 94948
rect 359550 94936 359556 94948
rect 359608 94936 359614 94988
rect 365806 94936 365812 94988
rect 365864 94976 365870 94988
rect 373966 94976 373994 95016
rect 393958 95004 393964 95016
rect 394016 95004 394022 95056
rect 421006 95044 421012 95056
rect 402946 95016 421012 95044
rect 365864 94948 373994 94976
rect 365864 94936 365870 94948
rect 376662 94936 376668 94988
rect 376720 94976 376726 94988
rect 387058 94976 387064 94988
rect 376720 94948 387064 94976
rect 376720 94936 376726 94948
rect 387058 94936 387064 94948
rect 387116 94936 387122 94988
rect 393406 94936 393412 94988
rect 393464 94976 393470 94988
rect 402946 94976 402974 95016
rect 421006 95004 421012 95016
rect 421064 95004 421070 95056
rect 430666 95004 430672 95056
rect 430724 95044 430730 95056
rect 442258 95044 442264 95056
rect 430724 95016 442264 95044
rect 430724 95004 430730 95016
rect 442258 95004 442264 95016
rect 442316 95004 442322 95056
rect 447226 95004 447232 95056
rect 447284 95044 447290 95056
rect 475010 95044 475016 95056
rect 447284 95016 475016 95044
rect 447284 95004 447290 95016
rect 475010 95004 475016 95016
rect 475068 95004 475074 95056
rect 484670 95004 484676 95056
rect 484728 95044 484734 95056
rect 496078 95044 496084 95056
rect 484728 95016 496084 95044
rect 484728 95004 484734 95016
rect 496078 95004 496084 95016
rect 496136 95004 496142 95056
rect 501046 95004 501052 95056
rect 501104 95044 501110 95056
rect 529014 95044 529020 95056
rect 501104 95016 529020 95044
rect 501104 95004 501110 95016
rect 529014 95004 529020 95016
rect 529072 95004 529078 95056
rect 393464 94948 402974 94976
rect 393464 94936 393470 94948
rect 403710 94936 403716 94988
rect 403768 94976 403774 94988
rect 414658 94976 414664 94988
rect 403768 94948 414664 94976
rect 403768 94936 403774 94948
rect 414658 94936 414664 94948
rect 414716 94936 414722 94988
rect 457714 94936 457720 94988
rect 457772 94976 457778 94988
rect 468478 94976 468484 94988
rect 457772 94948 468484 94976
rect 457772 94936 457778 94948
rect 468478 94936 468484 94948
rect 468536 94936 468542 94988
rect 511718 94936 511724 94988
rect 511776 94976 511782 94988
rect 522298 94976 522304 94988
rect 511776 94948 522304 94976
rect 511776 94936 511782 94948
rect 522298 94936 522304 94948
rect 522356 94936 522362 94988
rect 36538 94868 36544 94920
rect 36596 94908 36602 94920
rect 538674 94908 538680 94920
rect 36596 94880 538680 94908
rect 36596 94868 36602 94880
rect 538674 94868 538680 94880
rect 538732 94868 538738 94920
rect 15286 91740 15292 91792
rect 15344 91780 15350 91792
rect 529014 91780 529020 91792
rect 15344 91752 529020 91780
rect 15344 91740 15350 91752
rect 529014 91740 529020 91752
rect 529072 91740 529078 91792
rect 25682 91332 25688 91384
rect 25740 91372 25746 91384
rect 149698 91372 149704 91384
rect 25740 91344 149704 91372
rect 25740 91332 25746 91344
rect 149698 91332 149704 91344
rect 149756 91332 149762 91384
rect 36538 91264 36544 91316
rect 36596 91304 36602 91316
rect 52638 91304 52644 91316
rect 36596 91276 52644 91304
rect 36596 91264 36602 91276
rect 52638 91264 52644 91276
rect 52696 91264 52702 91316
rect 475010 91264 475016 91316
rect 475068 91304 475074 91316
rect 494698 91304 494704 91316
rect 475068 91276 494704 91304
rect 475068 91264 475074 91276
rect 494698 91264 494704 91276
rect 494756 91264 494762 91316
rect 43070 91196 43076 91248
rect 43128 91236 43134 91248
rect 62758 91236 62764 91248
rect 43128 91208 62764 91236
rect 43128 91196 43134 91208
rect 62758 91196 62764 91208
rect 62816 91196 62822 91248
rect 90450 91196 90456 91248
rect 90508 91236 90514 91248
rect 106642 91236 106648 91248
rect 90508 91208 106648 91236
rect 90508 91196 90514 91208
rect 106642 91196 106648 91208
rect 106700 91196 106706 91248
rect 116486 91196 116492 91248
rect 116544 91236 116550 91248
rect 133690 91236 133696 91248
rect 116544 91208 133696 91236
rect 116544 91196 116550 91208
rect 133690 91196 133696 91208
rect 133748 91196 133754 91248
rect 144270 91196 144276 91248
rect 144328 91236 144334 91248
rect 160646 91236 160652 91248
rect 144328 91208 160652 91236
rect 144328 91196 144334 91208
rect 160646 91196 160652 91208
rect 160704 91196 160710 91248
rect 170490 91196 170496 91248
rect 170548 91236 170554 91248
rect 187694 91236 187700 91248
rect 170548 91208 187700 91236
rect 170548 91196 170554 91208
rect 187694 91196 187700 91208
rect 187752 91196 187758 91248
rect 197446 91196 197452 91248
rect 197504 91236 197510 91248
rect 214650 91236 214656 91248
rect 197504 91208 214656 91236
rect 197504 91196 197510 91208
rect 214650 91196 214656 91208
rect 214708 91196 214714 91248
rect 224494 91196 224500 91248
rect 224552 91236 224558 91248
rect 241698 91236 241704 91248
rect 224552 91208 241704 91236
rect 224552 91196 224558 91208
rect 241698 91196 241704 91208
rect 241756 91196 241762 91248
rect 251450 91196 251456 91248
rect 251508 91236 251514 91248
rect 268654 91236 268660 91248
rect 251508 91208 268660 91236
rect 251508 91196 251514 91208
rect 268654 91196 268660 91208
rect 268712 91196 268718 91248
rect 413462 91196 413468 91248
rect 413520 91236 413526 91248
rect 430666 91236 430672 91248
rect 413520 91208 430672 91236
rect 413520 91196 413526 91208
rect 430666 91196 430672 91208
rect 430724 91196 430730 91248
rect 440510 91196 440516 91248
rect 440568 91236 440574 91248
rect 457622 91236 457628 91248
rect 440568 91208 457628 91236
rect 440568 91196 440574 91208
rect 457622 91196 457628 91208
rect 457680 91196 457686 91248
rect 468478 91196 468484 91248
rect 468536 91236 468542 91248
rect 484670 91236 484676 91248
rect 468536 91208 484676 91236
rect 468536 91196 468542 91208
rect 484670 91196 484676 91208
rect 484728 91196 484734 91248
rect 36814 91128 36820 91180
rect 36872 91168 36878 91180
rect 62298 91168 62304 91180
rect 36872 91140 62304 91168
rect 36872 91128 36878 91140
rect 62298 91128 62304 91140
rect 62356 91128 62362 91180
rect 64138 91128 64144 91180
rect 64196 91168 64202 91180
rect 89346 91168 89352 91180
rect 64196 91140 89352 91168
rect 64196 91128 64202 91140
rect 89346 91128 89352 91140
rect 89404 91128 89410 91180
rect 90358 91128 90364 91180
rect 90416 91168 90422 91180
rect 116302 91168 116308 91180
rect 90416 91140 116308 91168
rect 90416 91128 90422 91140
rect 116302 91128 116308 91140
rect 116360 91128 116366 91180
rect 116578 91128 116584 91180
rect 116636 91168 116642 91180
rect 143350 91168 143356 91180
rect 116636 91140 143356 91168
rect 116636 91128 116642 91140
rect 143350 91128 143356 91140
rect 143408 91128 143414 91180
rect 144178 91128 144184 91180
rect 144236 91168 144242 91180
rect 170306 91168 170312 91180
rect 144236 91140 170312 91168
rect 144236 91128 144242 91140
rect 170306 91128 170312 91140
rect 170364 91128 170370 91180
rect 178034 91128 178040 91180
rect 178092 91168 178098 91180
rect 200758 91168 200764 91180
rect 178092 91140 200764 91168
rect 178092 91128 178098 91140
rect 200758 91128 200764 91140
rect 200816 91128 200822 91180
rect 232038 91128 232044 91180
rect 232096 91168 232102 91180
rect 251818 91168 251824 91180
rect 232096 91140 251824 91168
rect 232096 91128 232102 91140
rect 251818 91128 251824 91140
rect 251876 91128 251882 91180
rect 279418 91128 279424 91180
rect 279476 91168 279482 91180
rect 295702 91168 295708 91180
rect 279476 91140 295708 91168
rect 279476 91128 279482 91140
rect 295702 91128 295708 91140
rect 295760 91128 295766 91180
rect 305454 91128 305460 91180
rect 305512 91168 305518 91180
rect 322658 91168 322664 91180
rect 305512 91140 322664 91168
rect 305512 91128 305518 91140
rect 322658 91128 322664 91140
rect 322716 91128 322722 91180
rect 334618 91128 334624 91180
rect 334676 91168 334682 91180
rect 349706 91168 349712 91180
rect 334676 91140 349712 91168
rect 334676 91128 334682 91140
rect 349706 91128 349712 91140
rect 349764 91128 349770 91180
rect 359458 91128 359464 91180
rect 359516 91168 359522 91180
rect 376662 91168 376668 91180
rect 359516 91140 376668 91168
rect 359516 91128 359522 91140
rect 376662 91128 376668 91140
rect 376720 91128 376726 91180
rect 386506 91128 386512 91180
rect 386564 91168 386570 91180
rect 403618 91168 403624 91180
rect 386564 91140 403624 91168
rect 386564 91128 386570 91140
rect 403618 91128 403624 91140
rect 403676 91128 403682 91180
rect 421006 91128 421012 91180
rect 421064 91168 421070 91180
rect 443638 91168 443644 91180
rect 421064 91140 443644 91168
rect 421064 91128 421070 91140
rect 443638 91128 443644 91140
rect 443696 91128 443702 91180
rect 494514 91128 494520 91180
rect 494572 91168 494578 91180
rect 511626 91168 511632 91180
rect 494572 91140 511632 91168
rect 494572 91128 494578 91140
rect 511626 91128 511632 91140
rect 511684 91128 511690 91180
rect 522298 91128 522304 91180
rect 522356 91168 522362 91180
rect 538674 91168 538680 91180
rect 522356 91140 538680 91168
rect 522356 91128 522362 91140
rect 538674 91128 538680 91140
rect 538732 91128 538738 91180
rect 62482 91060 62488 91112
rect 62540 91100 62546 91112
rect 79686 91100 79692 91112
rect 62540 91072 79692 91100
rect 62540 91060 62546 91072
rect 79686 91060 79692 91072
rect 79744 91060 79750 91112
rect 171778 91060 171784 91112
rect 171836 91100 171842 91112
rect 197354 91100 197360 91112
rect 171836 91072 197360 91100
rect 171836 91060 171842 91072
rect 197354 91060 197360 91072
rect 197412 91060 197418 91112
rect 199378 91060 199384 91112
rect 199436 91100 199442 91112
rect 224310 91100 224316 91112
rect 199436 91072 224316 91100
rect 199436 91060 199442 91072
rect 224310 91060 224316 91072
rect 224368 91060 224374 91112
rect 225598 91060 225604 91112
rect 225656 91100 225662 91112
rect 251358 91100 251364 91112
rect 225656 91072 251364 91100
rect 225656 91060 225662 91072
rect 251358 91060 251364 91072
rect 251416 91060 251422 91112
rect 253198 91060 253204 91112
rect 253256 91100 253262 91112
rect 278314 91100 278320 91112
rect 253256 91072 278320 91100
rect 253256 91060 253262 91072
rect 278314 91060 278320 91072
rect 278372 91060 278378 91112
rect 279510 91060 279516 91112
rect 279568 91100 279574 91112
rect 305362 91100 305368 91112
rect 279568 91072 305368 91100
rect 279568 91060 279574 91072
rect 305362 91060 305368 91072
rect 305420 91060 305426 91112
rect 307018 91060 307024 91112
rect 307076 91100 307082 91112
rect 332318 91100 332324 91112
rect 307076 91072 332324 91100
rect 307076 91060 307082 91072
rect 332318 91060 332324 91072
rect 332376 91060 332382 91112
rect 333238 91060 333244 91112
rect 333296 91100 333302 91112
rect 359366 91100 359372 91112
rect 333296 91072 359372 91100
rect 333296 91060 333302 91072
rect 359366 91060 359372 91072
rect 359424 91060 359430 91112
rect 359550 91060 359556 91112
rect 359608 91100 359614 91112
rect 386322 91100 386328 91112
rect 359608 91072 386328 91100
rect 359608 91060 359614 91072
rect 386322 91060 386328 91072
rect 386380 91060 386386 91112
rect 387058 91060 387064 91112
rect 387116 91100 387122 91112
rect 413278 91100 413284 91112
rect 387116 91072 413284 91100
rect 387116 91060 387122 91072
rect 413278 91060 413284 91072
rect 413336 91060 413342 91112
rect 414658 91060 414664 91112
rect 414716 91100 414722 91112
rect 440326 91100 440332 91112
rect 414716 91072 440332 91100
rect 414716 91060 414722 91072
rect 440326 91060 440332 91072
rect 440384 91060 440390 91112
rect 442258 91060 442264 91112
rect 442316 91100 442322 91112
rect 467282 91100 467288 91112
rect 442316 91072 467288 91100
rect 442316 91060 442322 91072
rect 467282 91060 467288 91072
rect 467340 91060 467346 91112
rect 468570 91060 468576 91112
rect 468628 91100 468634 91112
rect 494330 91100 494336 91112
rect 468628 91072 494336 91100
rect 468628 91060 468634 91072
rect 494330 91060 494336 91072
rect 494388 91060 494394 91112
rect 496078 91060 496084 91112
rect 496136 91100 496142 91112
rect 521286 91100 521292 91112
rect 496136 91072 521292 91100
rect 496136 91060 496142 91072
rect 521286 91060 521292 91072
rect 521344 91060 521350 91112
rect 522390 91060 522396 91112
rect 522448 91100 522454 91112
rect 548334 91100 548340 91112
rect 522448 91072 548340 91100
rect 522448 91060 522454 91072
rect 548334 91060 548340 91072
rect 548392 91060 548398 91112
rect 37918 90312 37924 90364
rect 37976 90352 37982 90364
rect 526438 90352 526444 90364
rect 37976 90324 526444 90352
rect 37976 90312 37982 90324
rect 526438 90312 526444 90324
rect 526496 90312 526502 90364
rect 68922 88476 68928 88528
rect 68980 88516 68986 88528
rect 118694 88516 118700 88528
rect 68980 88488 118700 88516
rect 68980 88476 68986 88488
rect 118694 88476 118700 88488
rect 118752 88476 118758 88528
rect 230382 88476 230388 88528
rect 230440 88516 230446 88528
rect 280154 88516 280160 88528
rect 230440 88488 280160 88516
rect 230440 88476 230446 88488
rect 280154 88476 280160 88488
rect 280212 88476 280218 88528
rect 35618 88408 35624 88460
rect 35676 88448 35682 88460
rect 36630 88448 36636 88460
rect 35676 88420 36636 88448
rect 35676 88408 35682 88420
rect 36630 88408 36636 88420
rect 36688 88408 36694 88460
rect 41322 88408 41328 88460
rect 41380 88448 41386 88460
rect 91094 88448 91100 88460
rect 41380 88420 91100 88448
rect 41380 88408 41386 88420
rect 91094 88408 91100 88420
rect 91152 88408 91158 88460
rect 122742 88408 122748 88460
rect 122800 88448 122806 88460
rect 172514 88448 172520 88460
rect 122800 88420 172520 88448
rect 122800 88408 122806 88420
rect 172514 88408 172520 88420
rect 172572 88408 172578 88460
rect 176562 88408 176568 88460
rect 176620 88448 176626 88460
rect 226334 88448 226340 88460
rect 176620 88420 226340 88448
rect 176620 88408 176626 88420
rect 226334 88408 226340 88420
rect 226392 88408 226398 88460
rect 256602 88408 256608 88460
rect 256660 88448 256666 88460
rect 307754 88448 307760 88460
rect 256660 88420 307760 88448
rect 256660 88408 256666 88420
rect 307754 88408 307760 88420
rect 307812 88408 307818 88460
rect 311802 88408 311808 88460
rect 311860 88448 311866 88460
rect 361574 88448 361580 88460
rect 311860 88420 361580 88448
rect 311860 88408 311866 88420
rect 361574 88408 361580 88420
rect 361632 88408 361638 88460
rect 365622 88408 365628 88460
rect 365680 88448 365686 88460
rect 415394 88448 415400 88460
rect 365680 88420 415400 88448
rect 365680 88408 365686 88420
rect 415394 88408 415400 88420
rect 415452 88408 415458 88460
rect 419442 88408 419448 88460
rect 419500 88448 419506 88460
rect 469214 88448 469220 88460
rect 419500 88420 469220 88448
rect 419500 88408 419506 88420
rect 469214 88408 469220 88420
rect 469272 88408 469278 88460
rect 473262 88408 473268 88460
rect 473320 88448 473326 88460
rect 523034 88448 523040 88460
rect 473320 88420 523040 88448
rect 473320 88408 473326 88420
rect 523034 88408 523040 88420
rect 523092 88408 523098 88460
rect 13722 88340 13728 88392
rect 13780 88380 13786 88392
rect 64874 88380 64880 88392
rect 13780 88352 64880 88380
rect 13780 88340 13786 88352
rect 64874 88340 64880 88352
rect 64932 88340 64938 88392
rect 95142 88340 95148 88392
rect 95200 88380 95206 88392
rect 146294 88380 146300 88392
rect 95200 88352 146300 88380
rect 95200 88340 95206 88352
rect 146294 88340 146300 88352
rect 146352 88340 146358 88392
rect 148962 88340 148968 88392
rect 149020 88380 149026 88392
rect 200114 88380 200120 88392
rect 149020 88352 200120 88380
rect 149020 88340 149026 88352
rect 200114 88340 200120 88352
rect 200172 88340 200178 88392
rect 202782 88340 202788 88392
rect 202840 88380 202846 88392
rect 253934 88380 253940 88392
rect 202840 88352 253940 88380
rect 202840 88340 202846 88352
rect 253934 88340 253940 88352
rect 253992 88340 253998 88392
rect 284202 88340 284208 88392
rect 284260 88380 284266 88392
rect 335354 88380 335360 88392
rect 284260 88352 335360 88380
rect 284260 88340 284266 88352
rect 335354 88340 335360 88352
rect 335412 88340 335418 88392
rect 338022 88340 338028 88392
rect 338080 88380 338086 88392
rect 389174 88380 389180 88392
rect 338080 88352 389180 88380
rect 338080 88340 338086 88352
rect 389174 88340 389180 88352
rect 389232 88340 389238 88392
rect 391842 88340 391848 88392
rect 391900 88380 391906 88392
rect 442994 88380 443000 88392
rect 391900 88352 443000 88380
rect 391900 88340 391906 88352
rect 442994 88340 443000 88352
rect 443052 88340 443058 88392
rect 445662 88340 445668 88392
rect 445720 88380 445726 88392
rect 496814 88380 496820 88392
rect 445720 88352 496820 88380
rect 445720 88340 445726 88352
rect 496814 88340 496820 88352
rect 496872 88340 496878 88392
rect 500862 88340 500868 88392
rect 500920 88380 500926 88392
rect 550634 88380 550640 88392
rect 500920 88352 550640 88380
rect 500920 88340 500926 88352
rect 550634 88340 550640 88352
rect 550692 88340 550698 88392
rect 89714 72292 89720 72344
rect 89772 72332 89778 72344
rect 90450 72332 90456 72344
rect 89772 72304 90456 72332
rect 89772 72292 89778 72304
rect 90450 72292 90456 72304
rect 90508 72292 90514 72344
rect 143626 72292 143632 72344
rect 143684 72332 143690 72344
rect 144270 72332 144276 72344
rect 143684 72304 144276 72332
rect 143684 72292 143690 72304
rect 144270 72292 144276 72304
rect 144328 72292 144334 72344
rect 332502 71680 332508 71732
rect 332560 71720 332566 71732
rect 334618 71720 334624 71732
rect 332560 71692 334624 71720
rect 332560 71680 332566 71692
rect 334618 71680 334624 71692
rect 334676 71680 334682 71732
rect 116210 70592 116216 70644
rect 116268 70632 116274 70644
rect 116486 70632 116492 70644
rect 116268 70604 116492 70632
rect 116268 70592 116274 70604
rect 116486 70592 116492 70604
rect 116544 70592 116550 70644
rect 170214 70592 170220 70644
rect 170272 70632 170278 70644
rect 170490 70632 170496 70644
rect 170272 70604 170496 70632
rect 170272 70592 170278 70604
rect 170490 70592 170496 70604
rect 170548 70592 170554 70644
rect 53098 68960 53104 69012
rect 53156 69000 53162 69012
rect 64138 69000 64144 69012
rect 53156 68972 64144 69000
rect 53156 68960 53162 68972
rect 64138 68960 64144 68972
rect 64196 68960 64202 69012
rect 69106 68960 69112 69012
rect 69164 69000 69170 69012
rect 69164 68972 74534 69000
rect 69164 68960 69170 68972
rect 15194 68892 15200 68944
rect 15252 68932 15258 68944
rect 42794 68932 42800 68944
rect 15252 68904 42800 68932
rect 15252 68892 15258 68904
rect 42794 68892 42800 68904
rect 42852 68892 42858 68944
rect 62758 68892 62764 68944
rect 62816 68932 62822 68944
rect 69750 68932 69756 68944
rect 62816 68904 69756 68932
rect 62816 68892 62822 68904
rect 69750 68892 69756 68904
rect 69808 68892 69814 68944
rect 74506 68932 74534 68972
rect 96706 68960 96712 69012
rect 96764 69000 96770 69012
rect 96764 68972 103514 69000
rect 96764 68960 96770 68972
rect 96798 68932 96804 68944
rect 74506 68904 96804 68932
rect 96798 68892 96804 68904
rect 96856 68892 96862 68944
rect 103486 68932 103514 68972
rect 146938 68960 146944 69012
rect 146996 69000 147002 69012
rect 146996 68972 151814 69000
rect 146996 68960 147002 68972
rect 123662 68932 123668 68944
rect 103486 68904 123668 68932
rect 123662 68892 123668 68904
rect 123720 68892 123726 68944
rect 133782 68892 133788 68944
rect 133840 68932 133846 68944
rect 144178 68932 144184 68944
rect 133840 68904 144184 68932
rect 133840 68892 133846 68904
rect 144178 68892 144184 68904
rect 144236 68892 144242 68944
rect 150710 68932 150716 68944
rect 146588 68904 150716 68932
rect 25958 68824 25964 68876
rect 26016 68864 26022 68876
rect 36814 68864 36820 68876
rect 26016 68836 36820 68864
rect 26016 68824 26022 68836
rect 36814 68824 36820 68836
rect 36872 68824 36878 68876
rect 79962 68824 79968 68876
rect 80020 68864 80026 68876
rect 90358 68864 90364 68876
rect 80020 68836 90364 68864
rect 80020 68824 80026 68836
rect 90358 68824 90364 68836
rect 90416 68824 90422 68876
rect 106550 68824 106556 68876
rect 106608 68864 106614 68876
rect 116578 68864 116584 68876
rect 106608 68836 116584 68864
rect 106608 68824 106614 68836
rect 116578 68824 116584 68836
rect 116636 68824 116642 68876
rect 122926 68824 122932 68876
rect 122984 68864 122990 68876
rect 146588 68864 146616 68904
rect 150710 68892 150716 68904
rect 150768 68892 150774 68944
rect 151786 68932 151814 68972
rect 200758 68960 200764 69012
rect 200816 69000 200822 69012
rect 204622 69000 204628 69012
rect 200816 68972 204628 69000
rect 200816 68960 200822 68972
rect 204622 68960 204628 68972
rect 204680 68960 204686 69012
rect 251818 68960 251824 69012
rect 251876 69000 251882 69012
rect 258718 69000 258724 69012
rect 251876 68972 258724 69000
rect 251876 68960 251882 68972
rect 258718 68960 258724 68972
rect 258776 68960 258782 69012
rect 443638 68960 443644 69012
rect 443696 69000 443702 69012
rect 447686 69000 447692 69012
rect 443696 68972 447692 69000
rect 443696 68960 443702 68972
rect 447686 68960 447692 68972
rect 447744 68960 447750 69012
rect 494698 68960 494704 69012
rect 494756 69000 494762 69012
rect 501598 69000 501604 69012
rect 494756 68972 501604 69000
rect 494756 68960 494762 68972
rect 501598 68960 501604 68972
rect 501656 68960 501662 69012
rect 548058 68932 548064 68944
rect 151786 68904 548064 68932
rect 548058 68892 548064 68904
rect 548116 68892 548122 68944
rect 122984 68836 146616 68864
rect 122984 68824 122990 68836
rect 150526 68824 150532 68876
rect 150584 68864 150590 68876
rect 178126 68864 178132 68876
rect 150584 68836 178132 68864
rect 150584 68824 150590 68836
rect 178126 68824 178132 68836
rect 178184 68824 178190 68876
rect 187970 68824 187976 68876
rect 188028 68864 188034 68876
rect 199378 68864 199384 68876
rect 188028 68836 199384 68864
rect 188028 68824 188034 68836
rect 199378 68824 199384 68836
rect 199436 68824 199442 68876
rect 204346 68824 204352 68876
rect 204404 68864 204410 68876
rect 231854 68864 231860 68876
rect 204404 68836 231860 68864
rect 204404 68824 204410 68836
rect 231854 68824 231860 68836
rect 231912 68824 231918 68876
rect 242066 68824 242072 68876
rect 242124 68864 242130 68876
rect 253198 68864 253204 68876
rect 242124 68836 253204 68864
rect 242124 68824 242130 68836
rect 253198 68824 253204 68836
rect 253256 68824 253262 68876
rect 258166 68824 258172 68876
rect 258224 68864 258230 68876
rect 258224 68836 281764 68864
rect 258224 68824 258230 68836
rect 160554 68756 160560 68808
rect 160612 68796 160618 68808
rect 171778 68796 171784 68808
rect 160612 68768 171784 68796
rect 160612 68756 160618 68768
rect 171778 68756 171784 68768
rect 171836 68756 171842 68808
rect 215018 68756 215024 68808
rect 215076 68796 215082 68808
rect 225598 68796 225604 68808
rect 215076 68768 225604 68796
rect 215076 68756 215082 68768
rect 225598 68756 225604 68768
rect 225656 68756 225662 68808
rect 268930 68756 268936 68808
rect 268988 68796 268994 68808
rect 279510 68796 279516 68808
rect 268988 68768 279516 68796
rect 268988 68756 268994 68768
rect 279510 68756 279516 68768
rect 279568 68756 279574 68808
rect 281736 68796 281764 68836
rect 285766 68824 285772 68876
rect 285824 68864 285830 68876
rect 312630 68864 312636 68876
rect 285824 68836 312636 68864
rect 285824 68824 285830 68836
rect 312630 68824 312636 68836
rect 312688 68824 312694 68876
rect 340138 68864 340144 68876
rect 316006 68836 340144 68864
rect 286134 68796 286140 68808
rect 281736 68768 286140 68796
rect 286134 68756 286140 68768
rect 286192 68756 286198 68808
rect 295978 68756 295984 68808
rect 296036 68796 296042 68808
rect 307018 68796 307024 68808
rect 296036 68768 307024 68796
rect 296036 68756 296042 68768
rect 307018 68756 307024 68768
rect 307076 68756 307082 68808
rect 311986 68756 311992 68808
rect 312044 68796 312050 68808
rect 316006 68796 316034 68836
rect 340138 68824 340144 68836
rect 340196 68824 340202 68876
rect 344986 68836 364334 68864
rect 312044 68768 316034 68796
rect 312044 68756 312050 68768
rect 322842 68756 322848 68808
rect 322900 68796 322906 68808
rect 333238 68796 333244 68808
rect 322900 68768 333244 68796
rect 322900 68756 322906 68768
rect 333238 68756 333244 68768
rect 333296 68756 333302 68808
rect 339586 68756 339592 68808
rect 339644 68796 339650 68808
rect 344986 68796 345014 68836
rect 339644 68768 345014 68796
rect 339644 68756 339650 68768
rect 350074 68756 350080 68808
rect 350132 68796 350138 68808
rect 359550 68796 359556 68808
rect 350132 68768 359556 68796
rect 350132 68756 350138 68768
rect 359550 68756 359556 68768
rect 359608 68756 359614 68808
rect 364306 68796 364334 68836
rect 365806 68824 365812 68876
rect 365864 68864 365870 68876
rect 393590 68864 393596 68876
rect 365864 68836 393596 68864
rect 365864 68824 365870 68836
rect 393590 68824 393596 68836
rect 393648 68824 393654 68876
rect 420914 68864 420920 68876
rect 402946 68836 420920 68864
rect 366726 68796 366732 68808
rect 364306 68768 366732 68796
rect 366726 68756 366732 68768
rect 366784 68756 366790 68808
rect 376570 68756 376576 68808
rect 376628 68796 376634 68808
rect 387058 68796 387064 68808
rect 376628 68768 387064 68796
rect 376628 68756 376634 68768
rect 387058 68756 387064 68768
rect 387116 68756 387122 68808
rect 393406 68756 393412 68808
rect 393464 68796 393470 68808
rect 402946 68796 402974 68836
rect 420914 68824 420920 68836
rect 420972 68824 420978 68876
rect 431034 68824 431040 68876
rect 431092 68864 431098 68876
rect 442258 68864 442264 68876
rect 431092 68836 442264 68864
rect 431092 68824 431098 68836
rect 442258 68824 442264 68836
rect 442316 68824 442322 68876
rect 447226 68824 447232 68876
rect 447284 68864 447290 68876
rect 474734 68864 474740 68876
rect 447284 68836 474740 68864
rect 447284 68824 447290 68836
rect 474734 68824 474740 68836
rect 474792 68824 474798 68876
rect 484946 68824 484952 68876
rect 485004 68864 485010 68876
rect 496078 68864 496084 68876
rect 485004 68836 496084 68864
rect 485004 68824 485010 68836
rect 496078 68824 496084 68836
rect 496136 68824 496142 68876
rect 501046 68824 501052 68876
rect 501104 68864 501110 68876
rect 528738 68864 528744 68876
rect 501104 68836 528744 68864
rect 501104 68824 501110 68836
rect 528738 68824 528744 68836
rect 528796 68824 528802 68876
rect 393464 68768 402974 68796
rect 393464 68756 393470 68768
rect 403986 68756 403992 68808
rect 404044 68796 404050 68808
rect 414658 68796 414664 68808
rect 404044 68768 414664 68796
rect 404044 68756 404050 68768
rect 414658 68756 414664 68768
rect 414716 68756 414722 68808
rect 458082 68756 458088 68808
rect 458140 68796 458146 68808
rect 468570 68796 468576 68808
rect 458140 68768 468576 68796
rect 458140 68756 458146 68768
rect 468570 68756 468576 68768
rect 468628 68756 468634 68808
rect 511902 68756 511908 68808
rect 511960 68796 511966 68808
rect 522390 68796 522396 68808
rect 511960 68768 522396 68796
rect 511960 68756 511966 68768
rect 522390 68756 522396 68768
rect 522448 68756 522454 68808
rect 36722 68688 36728 68740
rect 36780 68728 36786 68740
rect 538398 68728 538404 68740
rect 36780 68700 538404 68728
rect 36780 68688 36786 68700
rect 538398 68688 538404 68700
rect 538456 68688 538462 68740
rect 16298 65492 16304 65544
rect 16356 65532 16362 65544
rect 528646 65532 528652 65544
rect 16356 65504 528652 65532
rect 16356 65492 16362 65504
rect 528646 65492 528652 65504
rect 528704 65492 528710 65544
rect 26050 65152 26056 65204
rect 26108 65192 26114 65204
rect 146938 65192 146944 65204
rect 26108 65164 146944 65192
rect 26108 65152 26114 65164
rect 146938 65152 146944 65164
rect 146996 65152 147002 65204
rect 36722 65084 36728 65136
rect 36780 65124 36786 65136
rect 52454 65124 52460 65136
rect 36780 65096 52460 65124
rect 36780 65084 36786 65096
rect 52454 65084 52460 65096
rect 52512 65084 52518 65136
rect 232314 65084 232320 65136
rect 232372 65124 232378 65136
rect 251818 65124 251824 65136
rect 232372 65096 251824 65124
rect 232372 65084 232378 65096
rect 251818 65084 251824 65096
rect 251876 65084 251882 65136
rect 475378 65084 475384 65136
rect 475436 65124 475442 65136
rect 494698 65124 494704 65136
rect 475436 65096 494704 65124
rect 475436 65084 475442 65096
rect 494698 65084 494704 65096
rect 494756 65084 494762 65136
rect 43346 65016 43352 65068
rect 43404 65056 43410 65068
rect 62758 65056 62764 65068
rect 43404 65028 62764 65056
rect 43404 65016 43410 65028
rect 62758 65016 62764 65028
rect 62816 65016 62822 65068
rect 90450 65016 90456 65068
rect 90508 65056 90514 65068
rect 106458 65056 106464 65068
rect 90508 65028 106464 65056
rect 90508 65016 90514 65028
rect 106458 65016 106464 65028
rect 106516 65016 106522 65068
rect 116486 65016 116492 65068
rect 116544 65056 116550 65068
rect 133414 65056 133420 65068
rect 116544 65028 133420 65056
rect 116544 65016 116550 65028
rect 133414 65016 133420 65028
rect 133472 65016 133478 65068
rect 170490 65016 170496 65068
rect 170548 65056 170554 65068
rect 187786 65056 187792 65068
rect 170548 65028 187792 65056
rect 170548 65016 170554 65028
rect 187786 65016 187792 65028
rect 187844 65016 187850 65068
rect 197538 65016 197544 65068
rect 197596 65056 197602 65068
rect 214374 65056 214380 65068
rect 197596 65028 214380 65056
rect 197596 65016 197602 65028
rect 214374 65016 214380 65028
rect 214432 65016 214438 65068
rect 224494 65016 224500 65068
rect 224552 65056 224558 65068
rect 241606 65056 241612 65068
rect 224552 65028 241612 65056
rect 224552 65016 224558 65028
rect 241606 65016 241612 65028
rect 241664 65016 241670 65068
rect 413462 65016 413468 65068
rect 413520 65056 413526 65068
rect 430574 65056 430580 65068
rect 413520 65028 430580 65056
rect 413520 65016 413526 65028
rect 430574 65016 430580 65028
rect 430632 65016 430638 65068
rect 440510 65016 440516 65068
rect 440568 65056 440574 65068
rect 457254 65056 457260 65068
rect 440568 65028 457260 65056
rect 440568 65016 440574 65028
rect 457254 65016 457260 65028
rect 457312 65016 457318 65068
rect 468570 65016 468576 65068
rect 468628 65056 468634 65068
rect 484394 65056 484400 65068
rect 468628 65028 484400 65056
rect 468628 65016 468634 65028
rect 484394 65016 484400 65028
rect 484452 65016 484458 65068
rect 36814 64948 36820 65000
rect 36872 64988 36878 65000
rect 62114 64988 62120 65000
rect 36872 64960 62120 64988
rect 36872 64948 36878 64960
rect 62114 64948 62120 64960
rect 62172 64948 62178 65000
rect 64138 64948 64144 65000
rect 64196 64988 64202 65000
rect 89070 64988 89076 65000
rect 64196 64960 89076 64988
rect 64196 64948 64202 64960
rect 89070 64948 89076 64960
rect 89128 64948 89134 65000
rect 90358 64948 90364 65000
rect 90416 64988 90422 65000
rect 116118 64988 116124 65000
rect 90416 64960 116124 64988
rect 90416 64948 90422 64960
rect 116118 64948 116124 64960
rect 116176 64948 116182 65000
rect 116578 64948 116584 65000
rect 116636 64988 116642 65000
rect 142982 64988 142988 65000
rect 116636 64960 142988 64988
rect 116636 64948 116642 64960
rect 142982 64948 142988 64960
rect 143040 64948 143046 65000
rect 144270 64948 144276 65000
rect 144328 64988 144334 65000
rect 170030 64988 170036 65000
rect 144328 64960 170036 64988
rect 144328 64948 144334 64960
rect 170030 64948 170036 64960
rect 170088 64948 170094 65000
rect 178402 64948 178408 65000
rect 178460 64988 178466 65000
rect 200758 64988 200764 65000
rect 178460 64960 200764 64988
rect 178460 64948 178466 64960
rect 200758 64948 200764 64960
rect 200816 64948 200822 65000
rect 251450 64948 251456 65000
rect 251508 64988 251514 65000
rect 268286 64988 268292 65000
rect 251508 64960 268292 64988
rect 251508 64948 251514 64960
rect 268286 64948 268292 64960
rect 268344 64948 268350 65000
rect 279418 64948 279424 65000
rect 279476 64988 279482 65000
rect 295794 64988 295800 65000
rect 279476 64960 295800 64988
rect 279476 64948 279482 64960
rect 295794 64948 295800 64960
rect 295852 64948 295858 65000
rect 305546 64948 305552 65000
rect 305604 64988 305610 65000
rect 322382 64988 322388 65000
rect 305604 64960 322388 64988
rect 305604 64948 305610 64960
rect 322382 64948 322388 64960
rect 322440 64948 322446 65000
rect 334618 64948 334624 65000
rect 334676 64988 334682 65000
rect 349798 64988 349804 65000
rect 334676 64960 349804 64988
rect 334676 64948 334682 64960
rect 349798 64948 349804 64960
rect 349856 64948 349862 65000
rect 359642 64948 359648 65000
rect 359700 64988 359706 65000
rect 376294 64988 376300 65000
rect 359700 64960 376300 64988
rect 359700 64948 359706 64960
rect 376294 64948 376300 64960
rect 376352 64948 376358 65000
rect 386506 64948 386512 65000
rect 386564 64988 386570 65000
rect 403342 64988 403348 65000
rect 386564 64960 403348 64988
rect 386564 64948 386570 64960
rect 403342 64948 403348 64960
rect 403400 64948 403406 65000
rect 421282 64948 421288 65000
rect 421340 64988 421346 65000
rect 443638 64988 443644 65000
rect 421340 64960 443644 64988
rect 421340 64948 421346 64960
rect 443638 64948 443644 64960
rect 443696 64948 443702 65000
rect 494514 64948 494520 65000
rect 494572 64988 494578 65000
rect 511350 64988 511356 65000
rect 494572 64960 511356 64988
rect 494572 64948 494578 64960
rect 511350 64948 511356 64960
rect 511408 64948 511414 65000
rect 522298 64948 522304 65000
rect 522356 64988 522362 65000
rect 538398 64988 538404 65000
rect 522356 64960 538404 64988
rect 522356 64948 522362 64960
rect 538398 64948 538404 64960
rect 538456 64948 538462 65000
rect 62482 64880 62488 64932
rect 62540 64920 62546 64932
rect 79318 64920 79324 64932
rect 62540 64892 79324 64920
rect 62540 64880 62546 64892
rect 79318 64880 79324 64892
rect 79376 64880 79382 64932
rect 144178 64880 144184 64932
rect 144236 64920 144242 64932
rect 160278 64920 160284 64932
rect 144236 64892 160284 64920
rect 144236 64880 144242 64892
rect 160278 64880 160284 64892
rect 160336 64880 160342 64932
rect 171778 64880 171784 64932
rect 171836 64920 171842 64932
rect 197446 64920 197452 64932
rect 171836 64892 197452 64920
rect 171836 64880 171842 64892
rect 197446 64880 197452 64892
rect 197504 64880 197510 64932
rect 199378 64880 199384 64932
rect 199436 64920 199442 64932
rect 223942 64920 223948 64932
rect 199436 64892 223948 64920
rect 199436 64880 199442 64892
rect 223942 64880 223948 64892
rect 224000 64880 224006 64932
rect 225598 64880 225604 64932
rect 225656 64920 225662 64932
rect 251266 64920 251272 64932
rect 225656 64892 251272 64920
rect 225656 64880 225662 64892
rect 251266 64880 251272 64892
rect 251324 64880 251330 64932
rect 253198 64880 253204 64932
rect 253256 64920 253262 64932
rect 278038 64920 278044 64932
rect 253256 64892 278044 64920
rect 253256 64880 253262 64892
rect 278038 64880 278044 64892
rect 278096 64880 278102 64932
rect 279510 64880 279516 64932
rect 279568 64920 279574 64932
rect 305454 64920 305460 64932
rect 279568 64892 305460 64920
rect 279568 64880 279574 64892
rect 305454 64880 305460 64892
rect 305512 64880 305518 64932
rect 307018 64880 307024 64932
rect 307076 64920 307082 64932
rect 331950 64920 331956 64932
rect 307076 64892 331956 64920
rect 307076 64880 307082 64892
rect 331950 64880 331956 64892
rect 332008 64880 332014 64932
rect 333238 64880 333244 64932
rect 333296 64920 333302 64932
rect 359458 64920 359464 64932
rect 333296 64892 359464 64920
rect 333296 64880 333302 64892
rect 359458 64880 359464 64892
rect 359516 64880 359522 64932
rect 359550 64880 359556 64932
rect 359608 64920 359614 64932
rect 386046 64920 386052 64932
rect 359608 64892 386052 64920
rect 359608 64880 359614 64892
rect 386046 64880 386052 64892
rect 386104 64880 386110 64932
rect 387058 64880 387064 64932
rect 387116 64920 387122 64932
rect 412910 64920 412916 64932
rect 387116 64892 412916 64920
rect 387116 64880 387122 64892
rect 412910 64880 412916 64892
rect 412968 64880 412974 64932
rect 414658 64880 414664 64932
rect 414716 64920 414722 64932
rect 440234 64920 440240 64932
rect 414716 64892 440240 64920
rect 414716 64880 414722 64892
rect 440234 64880 440240 64892
rect 440292 64880 440298 64932
rect 442258 64880 442264 64932
rect 442316 64920 442322 64932
rect 467006 64920 467012 64932
rect 442316 64892 467012 64920
rect 442316 64880 442322 64892
rect 467006 64880 467012 64892
rect 467064 64880 467070 64932
rect 468478 64880 468484 64932
rect 468536 64920 468542 64932
rect 494054 64920 494060 64932
rect 468536 64892 494060 64920
rect 468536 64880 468542 64892
rect 494054 64880 494060 64892
rect 494112 64880 494118 64932
rect 496078 64880 496084 64932
rect 496136 64920 496142 64932
rect 520918 64920 520924 64932
rect 496136 64892 520924 64920
rect 496136 64880 496142 64892
rect 520918 64880 520924 64892
rect 520976 64880 520982 64932
rect 522390 64880 522396 64932
rect 522448 64920 522454 64932
rect 547966 64920 547972 64932
rect 522448 64892 547972 64920
rect 522448 64880 522454 64892
rect 547966 64880 547972 64892
rect 548024 64880 548030 64932
rect 37918 62772 37924 62824
rect 37976 62812 37982 62824
rect 526438 62812 526444 62824
rect 37976 62784 526444 62812
rect 37976 62772 37982 62784
rect 526438 62772 526444 62784
rect 526496 62772 526502 62824
rect 285766 62364 285772 62416
rect 285824 62404 285830 62416
rect 286134 62404 286140 62416
rect 285824 62376 286140 62404
rect 285824 62364 285830 62376
rect 286134 62364 286140 62376
rect 286192 62364 286198 62416
rect 339586 62296 339592 62348
rect 339644 62336 339650 62348
rect 340138 62336 340144 62348
rect 339644 62308 340144 62336
rect 339644 62296 339650 62308
rect 340138 62296 340144 62308
rect 340196 62296 340202 62348
rect 68922 62160 68928 62212
rect 68980 62200 68986 62212
rect 118694 62200 118700 62212
rect 68980 62172 118700 62200
rect 68980 62160 68986 62172
rect 118694 62160 118700 62172
rect 118752 62160 118758 62212
rect 122742 62160 122748 62212
rect 122800 62200 122806 62212
rect 172514 62200 172520 62212
rect 122800 62172 172520 62200
rect 122800 62160 122806 62172
rect 172514 62160 172520 62172
rect 172572 62160 172578 62212
rect 230382 62160 230388 62212
rect 230440 62200 230446 62212
rect 280154 62200 280160 62212
rect 230440 62172 280160 62200
rect 230440 62160 230446 62172
rect 280154 62160 280160 62172
rect 280212 62160 280218 62212
rect 311802 62160 311808 62212
rect 311860 62200 311866 62212
rect 361574 62200 361580 62212
rect 311860 62172 361580 62200
rect 311860 62160 311866 62172
rect 361574 62160 361580 62172
rect 361632 62160 361638 62212
rect 473262 62160 473268 62212
rect 473320 62200 473326 62212
rect 523034 62200 523040 62212
rect 473320 62172 523040 62200
rect 473320 62160 473326 62172
rect 523034 62160 523040 62172
rect 523092 62160 523098 62212
rect 41322 62092 41328 62144
rect 41380 62132 41386 62144
rect 91094 62132 91100 62144
rect 41380 62104 91100 62132
rect 41380 62092 41386 62104
rect 91094 62092 91100 62104
rect 91152 62092 91158 62144
rect 148962 62092 148968 62144
rect 149020 62132 149026 62144
rect 200114 62132 200120 62144
rect 149020 62104 200120 62132
rect 149020 62092 149026 62104
rect 200114 62092 200120 62104
rect 200172 62092 200178 62144
rect 202782 62092 202788 62144
rect 202840 62132 202846 62144
rect 253934 62132 253940 62144
rect 202840 62104 253940 62132
rect 202840 62092 202846 62104
rect 253934 62092 253940 62104
rect 253992 62092 253998 62144
rect 284202 62092 284208 62144
rect 284260 62132 284266 62144
rect 335354 62132 335360 62144
rect 284260 62104 335360 62132
rect 284260 62092 284266 62104
rect 335354 62092 335360 62104
rect 335412 62092 335418 62144
rect 365622 62092 365628 62144
rect 365680 62132 365686 62144
rect 415394 62132 415400 62144
rect 365680 62104 415400 62132
rect 365680 62092 365686 62104
rect 415394 62092 415400 62104
rect 415452 62092 415458 62144
rect 419442 62092 419448 62144
rect 419500 62132 419506 62144
rect 469214 62132 469220 62144
rect 419500 62104 469220 62132
rect 419500 62092 419506 62104
rect 469214 62092 469220 62104
rect 469272 62092 469278 62144
rect 500862 62092 500868 62144
rect 500920 62132 500926 62144
rect 550634 62132 550640 62144
rect 500920 62104 550640 62132
rect 500920 62092 500926 62104
rect 550634 62092 550640 62104
rect 550692 62092 550698 62144
rect 359550 60120 359556 60172
rect 359608 60120 359614 60172
rect 359568 59968 359596 60120
rect 359550 59916 359556 59968
rect 359608 59916 359614 59968
rect 89714 50328 89720 50380
rect 89772 50368 89778 50380
rect 90450 50368 90456 50380
rect 89772 50340 90456 50368
rect 89772 50328 89778 50340
rect 90450 50328 90456 50340
rect 90508 50328 90514 50380
rect 13722 44072 13728 44124
rect 13780 44112 13786 44124
rect 64874 44112 64880 44124
rect 13780 44084 64880 44112
rect 13780 44072 13786 44084
rect 64874 44072 64880 44084
rect 64932 44072 64938 44124
rect 95142 44072 95148 44124
rect 95200 44112 95206 44124
rect 146294 44112 146300 44124
rect 95200 44084 146300 44112
rect 95200 44072 95206 44084
rect 146294 44072 146300 44084
rect 146352 44072 146358 44124
rect 176562 44072 176568 44124
rect 176620 44112 176626 44124
rect 226334 44112 226340 44124
rect 176620 44084 226340 44112
rect 176620 44072 176626 44084
rect 226334 44072 226340 44084
rect 226392 44072 226398 44124
rect 256602 44072 256608 44124
rect 256660 44112 256666 44124
rect 307754 44112 307760 44124
rect 256660 44084 307760 44112
rect 256660 44072 256666 44084
rect 307754 44072 307760 44084
rect 307812 44072 307818 44124
rect 332502 44072 332508 44124
rect 332560 44112 332566 44124
rect 334618 44112 334624 44124
rect 332560 44084 334624 44112
rect 332560 44072 332566 44084
rect 334618 44072 334624 44084
rect 334676 44072 334682 44124
rect 338022 44072 338028 44124
rect 338080 44112 338086 44124
rect 389174 44112 389180 44124
rect 338080 44084 389180 44112
rect 338080 44072 338086 44084
rect 389174 44072 389180 44084
rect 389232 44072 389238 44124
rect 391842 44072 391848 44124
rect 391900 44112 391906 44124
rect 442994 44112 443000 44124
rect 391900 44084 443000 44112
rect 391900 44072 391906 44084
rect 442994 44072 443000 44084
rect 443052 44072 443058 44124
rect 445662 44072 445668 44124
rect 445720 44112 445726 44124
rect 496814 44112 496820 44124
rect 445720 44084 496820 44112
rect 445720 44072 445726 44084
rect 496814 44072 496820 44084
rect 496872 44072 496878 44124
rect 35618 44004 35624 44056
rect 35676 44044 35682 44056
rect 36722 44044 36728 44056
rect 35676 44016 36728 44044
rect 35676 44004 35682 44016
rect 36722 44004 36728 44016
rect 36780 44004 36786 44056
rect 467650 44004 467656 44056
rect 467708 44044 467714 44056
rect 468570 44044 468576 44056
rect 467708 44016 468576 44044
rect 467708 44004 467714 44016
rect 468570 44004 468576 44016
rect 468628 44004 468634 44056
rect 62758 41352 62764 41404
rect 62816 41392 62822 41404
rect 70026 41392 70032 41404
rect 62816 41364 70032 41392
rect 62816 41352 62822 41364
rect 70026 41352 70032 41364
rect 70084 41352 70090 41404
rect 96706 41352 96712 41404
rect 96764 41392 96770 41404
rect 96764 41364 103514 41392
rect 96764 41352 96770 41364
rect 15194 41284 15200 41336
rect 15252 41324 15258 41336
rect 42978 41324 42984 41336
rect 15252 41296 42984 41324
rect 15252 41284 15258 41296
rect 42978 41284 42984 41296
rect 43036 41284 43042 41336
rect 52730 41284 52736 41336
rect 52788 41324 52794 41336
rect 64138 41324 64144 41336
rect 52788 41296 64144 41324
rect 52788 41284 52794 41296
rect 64138 41284 64144 41296
rect 64196 41284 64202 41336
rect 69106 41284 69112 41336
rect 69164 41324 69170 41336
rect 96982 41324 96988 41336
rect 69164 41296 96988 41324
rect 69164 41284 69170 41296
rect 96982 41284 96988 41296
rect 97040 41284 97046 41336
rect 103486 41324 103514 41364
rect 200758 41352 200764 41404
rect 200816 41392 200822 41404
rect 204990 41392 204996 41404
rect 200816 41364 204996 41392
rect 200816 41352 200822 41364
rect 204990 41352 204996 41364
rect 205048 41352 205054 41404
rect 251818 41352 251824 41404
rect 251876 41392 251882 41404
rect 258994 41392 259000 41404
rect 251876 41364 259000 41392
rect 251876 41352 251882 41364
rect 258994 41352 259000 41364
rect 259052 41352 259058 41404
rect 443638 41352 443644 41404
rect 443696 41392 443702 41404
rect 447962 41392 447968 41404
rect 443696 41364 447968 41392
rect 443696 41352 443702 41364
rect 447962 41352 447968 41364
rect 448020 41352 448026 41404
rect 494698 41352 494704 41404
rect 494756 41392 494762 41404
rect 501966 41392 501972 41404
rect 494756 41364 501972 41392
rect 494756 41352 494762 41364
rect 501966 41352 501972 41364
rect 502024 41352 502030 41404
rect 124030 41324 124036 41336
rect 103486 41296 124036 41324
rect 124030 41284 124036 41296
rect 124088 41284 124094 41336
rect 149698 41284 149704 41336
rect 149756 41324 149762 41336
rect 548334 41324 548340 41336
rect 149756 41296 548340 41324
rect 149756 41284 149762 41296
rect 548334 41284 548340 41296
rect 548392 41284 548398 41336
rect 25682 41216 25688 41268
rect 25740 41256 25746 41268
rect 36814 41256 36820 41268
rect 25740 41228 36820 41256
rect 25740 41216 25746 41228
rect 36814 41216 36820 41228
rect 36872 41216 36878 41268
rect 79686 41216 79692 41268
rect 79744 41256 79750 41268
rect 90358 41256 90364 41268
rect 79744 41228 90364 41256
rect 79744 41216 79750 41228
rect 90358 41216 90364 41228
rect 90416 41216 90422 41268
rect 106642 41216 106648 41268
rect 106700 41256 106706 41268
rect 116578 41256 116584 41268
rect 106700 41228 116584 41256
rect 106700 41216 106706 41228
rect 116578 41216 116584 41228
rect 116636 41216 116642 41268
rect 133690 41216 133696 41268
rect 133748 41256 133754 41268
rect 144270 41256 144276 41268
rect 133748 41228 144276 41256
rect 133748 41216 133754 41228
rect 144270 41216 144276 41228
rect 144328 41216 144334 41268
rect 150526 41216 150532 41268
rect 150584 41256 150590 41268
rect 178034 41256 178040 41268
rect 150584 41228 178040 41256
rect 150584 41216 150590 41228
rect 178034 41216 178040 41228
rect 178092 41216 178098 41268
rect 187694 41216 187700 41268
rect 187752 41256 187758 41268
rect 199378 41256 199384 41268
rect 187752 41228 199384 41256
rect 187752 41216 187758 41228
rect 199378 41216 199384 41228
rect 199436 41216 199442 41268
rect 204346 41216 204352 41268
rect 204404 41256 204410 41268
rect 232038 41256 232044 41268
rect 204404 41228 232044 41256
rect 204404 41216 204410 41228
rect 232038 41216 232044 41228
rect 232096 41216 232102 41268
rect 241698 41216 241704 41268
rect 241756 41256 241762 41268
rect 253198 41256 253204 41268
rect 241756 41228 253204 41256
rect 241756 41216 241762 41228
rect 253198 41216 253204 41228
rect 253256 41216 253262 41268
rect 258166 41216 258172 41268
rect 258224 41256 258230 41268
rect 286042 41256 286048 41268
rect 258224 41228 286048 41256
rect 258224 41216 258230 41228
rect 286042 41216 286048 41228
rect 286100 41216 286106 41268
rect 312998 41256 313004 41268
rect 287026 41228 313004 41256
rect 122926 41148 122932 41200
rect 122984 41188 122990 41200
rect 150986 41188 150992 41200
rect 122984 41160 150992 41188
rect 122984 41148 122990 41160
rect 150986 41148 150992 41160
rect 151044 41148 151050 41200
rect 160646 41148 160652 41200
rect 160704 41188 160710 41200
rect 171778 41188 171784 41200
rect 160704 41160 171784 41188
rect 160704 41148 160710 41160
rect 171778 41148 171784 41160
rect 171836 41148 171842 41200
rect 214650 41148 214656 41200
rect 214708 41188 214714 41200
rect 225598 41188 225604 41200
rect 214708 41160 225604 41188
rect 214708 41148 214714 41160
rect 225598 41148 225604 41160
rect 225656 41148 225662 41200
rect 268654 41148 268660 41200
rect 268712 41188 268718 41200
rect 279510 41188 279516 41200
rect 268712 41160 279516 41188
rect 268712 41148 268718 41160
rect 279510 41148 279516 41160
rect 279568 41148 279574 41200
rect 285766 41148 285772 41200
rect 285824 41188 285830 41200
rect 287026 41188 287054 41228
rect 312998 41216 313004 41228
rect 313056 41216 313062 41268
rect 340046 41256 340052 41268
rect 316006 41228 340052 41256
rect 285824 41160 287054 41188
rect 285824 41148 285830 41160
rect 295702 41148 295708 41200
rect 295760 41188 295766 41200
rect 307018 41188 307024 41200
rect 295760 41160 307024 41188
rect 295760 41148 295766 41160
rect 307018 41148 307024 41160
rect 307076 41148 307082 41200
rect 311986 41148 311992 41200
rect 312044 41188 312050 41200
rect 316006 41188 316034 41228
rect 340046 41216 340052 41228
rect 340104 41216 340110 41268
rect 367002 41256 367008 41268
rect 344986 41228 367008 41256
rect 312044 41160 316034 41188
rect 312044 41148 312050 41160
rect 322658 41148 322664 41200
rect 322716 41188 322722 41200
rect 333238 41188 333244 41200
rect 322716 41160 333244 41188
rect 322716 41148 322722 41160
rect 333238 41148 333244 41160
rect 333296 41148 333302 41200
rect 339586 41148 339592 41200
rect 339644 41188 339650 41200
rect 344986 41188 345014 41228
rect 367002 41216 367008 41228
rect 367060 41216 367066 41268
rect 393958 41256 393964 41268
rect 373966 41228 393964 41256
rect 339644 41160 345014 41188
rect 339644 41148 339650 41160
rect 349706 41148 349712 41200
rect 349764 41188 349770 41200
rect 359550 41188 359556 41200
rect 349764 41160 359556 41188
rect 349764 41148 349770 41160
rect 359550 41148 359556 41160
rect 359608 41148 359614 41200
rect 365806 41148 365812 41200
rect 365864 41188 365870 41200
rect 373966 41188 373994 41228
rect 393958 41216 393964 41228
rect 394016 41216 394022 41268
rect 421006 41256 421012 41268
rect 402946 41228 421012 41256
rect 365864 41160 373994 41188
rect 365864 41148 365870 41160
rect 376662 41148 376668 41200
rect 376720 41188 376726 41200
rect 387058 41188 387064 41200
rect 376720 41160 387064 41188
rect 376720 41148 376726 41160
rect 387058 41148 387064 41160
rect 387116 41148 387122 41200
rect 393406 41148 393412 41200
rect 393464 41188 393470 41200
rect 402946 41188 402974 41228
rect 421006 41216 421012 41228
rect 421064 41216 421070 41268
rect 430666 41216 430672 41268
rect 430724 41256 430730 41268
rect 442258 41256 442264 41268
rect 430724 41228 442264 41256
rect 430724 41216 430730 41228
rect 442258 41216 442264 41228
rect 442316 41216 442322 41268
rect 447226 41216 447232 41268
rect 447284 41256 447290 41268
rect 475010 41256 475016 41268
rect 447284 41228 475016 41256
rect 447284 41216 447290 41228
rect 475010 41216 475016 41228
rect 475068 41216 475074 41268
rect 484670 41216 484676 41268
rect 484728 41256 484734 41268
rect 496078 41256 496084 41268
rect 484728 41228 496084 41256
rect 484728 41216 484734 41228
rect 496078 41216 496084 41228
rect 496136 41216 496142 41268
rect 501046 41216 501052 41268
rect 501104 41256 501110 41268
rect 529014 41256 529020 41268
rect 501104 41228 529020 41256
rect 501104 41216 501110 41228
rect 529014 41216 529020 41228
rect 529072 41216 529078 41268
rect 393464 41160 402974 41188
rect 393464 41148 393470 41160
rect 403710 41148 403716 41200
rect 403768 41188 403774 41200
rect 414658 41188 414664 41200
rect 403768 41160 414664 41188
rect 403768 41148 403774 41160
rect 414658 41148 414664 41160
rect 414716 41148 414722 41200
rect 457714 41148 457720 41200
rect 457772 41188 457778 41200
rect 468478 41188 468484 41200
rect 457772 41160 468484 41188
rect 457772 41148 457778 41160
rect 468478 41148 468484 41160
rect 468536 41148 468542 41200
rect 511718 41148 511724 41200
rect 511776 41188 511782 41200
rect 522390 41188 522396 41200
rect 511776 41160 522396 41188
rect 511776 41148 511782 41160
rect 522390 41148 522396 41160
rect 522448 41148 522454 41200
rect 36630 41080 36636 41132
rect 36688 41120 36694 41132
rect 538674 41120 538680 41132
rect 36688 41092 538680 41120
rect 36688 41080 36694 41092
rect 538674 41080 538680 41092
rect 538732 41080 538738 41132
rect 16022 38020 16028 38072
rect 16080 38060 16086 38072
rect 529014 38060 529020 38072
rect 16080 38032 529020 38060
rect 16080 38020 16086 38032
rect 529014 38020 529020 38032
rect 529072 38020 529078 38072
rect 35342 37952 35348 38004
rect 35400 37992 35406 38004
rect 580534 37992 580540 38004
rect 35400 37964 580540 37992
rect 35400 37952 35406 37964
rect 580534 37952 580540 37964
rect 580592 37952 580598 38004
rect 25682 37884 25688 37936
rect 25740 37924 25746 37936
rect 580350 37924 580356 37936
rect 25740 37896 580356 37924
rect 25740 37884 25746 37896
rect 580350 37884 580356 37896
rect 580408 37884 580414 37936
rect 43070 37476 43076 37528
rect 43128 37516 43134 37528
rect 62758 37516 62764 37528
rect 43128 37488 62764 37516
rect 43128 37476 43134 37488
rect 62758 37476 62764 37488
rect 62816 37476 62822 37528
rect 232038 37476 232044 37528
rect 232096 37516 232102 37528
rect 251818 37516 251824 37528
rect 232096 37488 251824 37516
rect 232096 37476 232102 37488
rect 251818 37476 251824 37488
rect 251876 37476 251882 37528
rect 36630 37408 36636 37460
rect 36688 37448 36694 37460
rect 52638 37448 52644 37460
rect 36688 37420 52644 37448
rect 36688 37408 36694 37420
rect 52638 37408 52644 37420
rect 52696 37408 52702 37460
rect 170490 37408 170496 37460
rect 170548 37448 170554 37460
rect 187694 37448 187700 37460
rect 170548 37420 187700 37448
rect 170548 37408 170554 37420
rect 187694 37408 187700 37420
rect 187752 37408 187758 37460
rect 197446 37408 197452 37460
rect 197504 37448 197510 37460
rect 214650 37448 214656 37460
rect 197504 37420 214656 37448
rect 197504 37408 197510 37420
rect 214650 37408 214656 37420
rect 214708 37408 214714 37460
rect 224494 37408 224500 37460
rect 224552 37448 224558 37460
rect 241698 37448 241704 37460
rect 224552 37420 241704 37448
rect 224552 37408 224558 37420
rect 241698 37408 241704 37420
rect 241756 37408 241762 37460
rect 413462 37408 413468 37460
rect 413520 37448 413526 37460
rect 430666 37448 430672 37460
rect 413520 37420 430672 37448
rect 413520 37408 413526 37420
rect 430666 37408 430672 37420
rect 430724 37408 430730 37460
rect 440510 37408 440516 37460
rect 440568 37448 440574 37460
rect 457622 37448 457628 37460
rect 440568 37420 457628 37448
rect 440568 37408 440574 37420
rect 457622 37408 457628 37420
rect 457680 37408 457686 37460
rect 468478 37408 468484 37460
rect 468536 37448 468542 37460
rect 484670 37448 484676 37460
rect 468536 37420 484676 37448
rect 468536 37408 468542 37420
rect 484670 37408 484676 37420
rect 484728 37408 484734 37460
rect 494514 37408 494520 37460
rect 494572 37448 494578 37460
rect 511626 37448 511632 37460
rect 494572 37420 511632 37448
rect 494572 37408 494578 37420
rect 511626 37408 511632 37420
rect 511684 37408 511690 37460
rect 62482 37340 62488 37392
rect 62540 37380 62546 37392
rect 79686 37380 79692 37392
rect 62540 37352 79692 37380
rect 62540 37340 62546 37352
rect 79686 37340 79692 37352
rect 79744 37340 79750 37392
rect 90358 37340 90364 37392
rect 90416 37380 90422 37392
rect 106642 37380 106648 37392
rect 90416 37352 106648 37380
rect 90416 37340 90422 37352
rect 106642 37340 106648 37352
rect 106700 37340 106706 37392
rect 116486 37340 116492 37392
rect 116544 37380 116550 37392
rect 133690 37380 133696 37392
rect 116544 37352 133696 37380
rect 116544 37340 116550 37352
rect 133690 37340 133696 37352
rect 133748 37340 133754 37392
rect 144178 37340 144184 37392
rect 144236 37380 144242 37392
rect 160646 37380 160652 37392
rect 144236 37352 160652 37380
rect 144236 37340 144242 37352
rect 160646 37340 160652 37352
rect 160704 37340 160710 37392
rect 178034 37340 178040 37392
rect 178092 37380 178098 37392
rect 200758 37380 200764 37392
rect 178092 37352 200764 37380
rect 178092 37340 178098 37352
rect 200758 37340 200764 37352
rect 200816 37340 200822 37392
rect 251450 37340 251456 37392
rect 251508 37380 251514 37392
rect 268654 37380 268660 37392
rect 251508 37352 268660 37380
rect 251508 37340 251514 37352
rect 268654 37340 268660 37352
rect 268712 37340 268718 37392
rect 279418 37340 279424 37392
rect 279476 37380 279482 37392
rect 295702 37380 295708 37392
rect 279476 37352 295708 37380
rect 279476 37340 279482 37352
rect 295702 37340 295708 37352
rect 295760 37340 295766 37392
rect 305454 37340 305460 37392
rect 305512 37380 305518 37392
rect 322658 37380 322664 37392
rect 305512 37352 322664 37380
rect 305512 37340 305518 37352
rect 322658 37340 322664 37352
rect 322716 37340 322722 37392
rect 335998 37340 336004 37392
rect 336056 37380 336062 37392
rect 349706 37380 349712 37392
rect 336056 37352 349712 37380
rect 336056 37340 336062 37352
rect 349706 37340 349712 37352
rect 349764 37340 349770 37392
rect 359458 37340 359464 37392
rect 359516 37380 359522 37392
rect 376662 37380 376668 37392
rect 359516 37352 376668 37380
rect 359516 37340 359522 37352
rect 376662 37340 376668 37352
rect 376720 37340 376726 37392
rect 386506 37340 386512 37392
rect 386564 37380 386570 37392
rect 403618 37380 403624 37392
rect 386564 37352 403624 37380
rect 386564 37340 386570 37352
rect 403618 37340 403624 37352
rect 403676 37340 403682 37392
rect 421006 37340 421012 37392
rect 421064 37380 421070 37392
rect 446398 37380 446404 37392
rect 421064 37352 446404 37380
rect 421064 37340 421070 37352
rect 446398 37340 446404 37352
rect 446456 37340 446462 37392
rect 475010 37340 475016 37392
rect 475068 37380 475074 37392
rect 494698 37380 494704 37392
rect 475068 37352 494704 37380
rect 475068 37340 475074 37352
rect 494698 37340 494704 37352
rect 494756 37340 494762 37392
rect 522390 37340 522396 37392
rect 522448 37380 522454 37392
rect 538674 37380 538680 37392
rect 522448 37352 538680 37380
rect 522448 37340 522454 37352
rect 538674 37340 538680 37352
rect 538732 37340 538738 37392
rect 36722 37272 36728 37324
rect 36780 37312 36786 37324
rect 62298 37312 62304 37324
rect 36780 37284 62304 37312
rect 36780 37272 36786 37284
rect 62298 37272 62304 37284
rect 62356 37272 62362 37324
rect 64138 37272 64144 37324
rect 64196 37312 64202 37324
rect 89346 37312 89352 37324
rect 64196 37284 89352 37312
rect 64196 37272 64202 37284
rect 89346 37272 89352 37284
rect 89404 37272 89410 37324
rect 90450 37272 90456 37324
rect 90508 37312 90514 37324
rect 116302 37312 116308 37324
rect 90508 37284 116308 37312
rect 90508 37272 90514 37284
rect 116302 37272 116308 37284
rect 116360 37272 116366 37324
rect 116578 37272 116584 37324
rect 116636 37312 116642 37324
rect 143350 37312 143356 37324
rect 116636 37284 143356 37312
rect 116636 37272 116642 37284
rect 143350 37272 143356 37284
rect 143408 37272 143414 37324
rect 144270 37272 144276 37324
rect 144328 37312 144334 37324
rect 170306 37312 170312 37324
rect 144328 37284 170312 37312
rect 144328 37272 144334 37284
rect 170306 37272 170312 37284
rect 170364 37272 170370 37324
rect 171778 37272 171784 37324
rect 171836 37312 171842 37324
rect 197354 37312 197360 37324
rect 171836 37284 197360 37312
rect 171836 37272 171842 37284
rect 197354 37272 197360 37284
rect 197412 37272 197418 37324
rect 199378 37272 199384 37324
rect 199436 37312 199442 37324
rect 224310 37312 224316 37324
rect 199436 37284 224316 37312
rect 199436 37272 199442 37284
rect 224310 37272 224316 37284
rect 224368 37272 224374 37324
rect 225598 37272 225604 37324
rect 225656 37312 225662 37324
rect 251358 37312 251364 37324
rect 225656 37284 251364 37312
rect 225656 37272 225662 37284
rect 251358 37272 251364 37284
rect 251416 37272 251422 37324
rect 253198 37272 253204 37324
rect 253256 37312 253262 37324
rect 278314 37312 278320 37324
rect 253256 37284 278320 37312
rect 253256 37272 253262 37284
rect 278314 37272 278320 37284
rect 278372 37272 278378 37324
rect 279510 37272 279516 37324
rect 279568 37312 279574 37324
rect 305362 37312 305368 37324
rect 279568 37284 305368 37312
rect 279568 37272 279574 37284
rect 305362 37272 305368 37284
rect 305420 37272 305426 37324
rect 307018 37272 307024 37324
rect 307076 37312 307082 37324
rect 332318 37312 332324 37324
rect 307076 37284 332324 37312
rect 307076 37272 307082 37284
rect 332318 37272 332324 37284
rect 332376 37272 332382 37324
rect 333238 37272 333244 37324
rect 333296 37312 333302 37324
rect 359366 37312 359372 37324
rect 333296 37284 359372 37312
rect 333296 37272 333302 37284
rect 359366 37272 359372 37284
rect 359424 37272 359430 37324
rect 359550 37272 359556 37324
rect 359608 37312 359614 37324
rect 386322 37312 386328 37324
rect 359608 37284 386328 37312
rect 359608 37272 359614 37284
rect 386322 37272 386328 37284
rect 386380 37272 386386 37324
rect 387058 37272 387064 37324
rect 387116 37312 387122 37324
rect 413278 37312 413284 37324
rect 387116 37284 413284 37312
rect 387116 37272 387122 37284
rect 413278 37272 413284 37284
rect 413336 37272 413342 37324
rect 414658 37272 414664 37324
rect 414716 37312 414722 37324
rect 440326 37312 440332 37324
rect 414716 37284 440332 37312
rect 414716 37272 414722 37284
rect 440326 37272 440332 37284
rect 440384 37272 440390 37324
rect 442258 37272 442264 37324
rect 442316 37312 442322 37324
rect 467282 37312 467288 37324
rect 442316 37284 467288 37312
rect 442316 37272 442322 37284
rect 467282 37272 467288 37284
rect 467340 37272 467346 37324
rect 468570 37272 468576 37324
rect 468628 37312 468634 37324
rect 494330 37312 494336 37324
rect 468628 37284 494336 37312
rect 468628 37272 468634 37284
rect 494330 37272 494336 37284
rect 494388 37272 494394 37324
rect 496078 37272 496084 37324
rect 496136 37312 496142 37324
rect 521286 37312 521292 37324
rect 496136 37284 521292 37312
rect 496136 37272 496142 37284
rect 521286 37272 521292 37284
rect 521344 37272 521350 37324
rect 522298 37272 522304 37324
rect 522356 37312 522362 37324
rect 548334 37312 548340 37324
rect 522356 37284 548340 37312
rect 522356 37272 522362 37284
rect 548334 37272 548340 37284
rect 548392 37272 548398 37324
rect 37918 36592 37924 36644
rect 37976 36632 37982 36644
rect 526438 36632 526444 36644
rect 37976 36604 526444 36632
rect 37976 36592 37982 36604
rect 526438 36592 526444 36604
rect 526496 36592 526502 36644
rect 38010 36524 38016 36576
rect 38068 36564 38074 36576
rect 580442 36564 580448 36576
rect 38068 36536 580448 36564
rect 38068 36524 38074 36536
rect 580442 36524 580448 36536
rect 580500 36524 580506 36576
rect 68922 34620 68928 34672
rect 68980 34660 68986 34672
rect 118694 34660 118700 34672
rect 68980 34632 118700 34660
rect 68980 34620 68986 34632
rect 118694 34620 118700 34632
rect 118752 34620 118758 34672
rect 311802 34620 311808 34672
rect 311860 34660 311866 34672
rect 361574 34660 361580 34672
rect 311860 34632 361580 34660
rect 311860 34620 311866 34632
rect 361574 34620 361580 34632
rect 361632 34620 361638 34672
rect 41322 34552 41328 34604
rect 41380 34592 41386 34604
rect 91094 34592 91100 34604
rect 41380 34564 91100 34592
rect 41380 34552 41386 34564
rect 91094 34552 91100 34564
rect 91152 34552 91158 34604
rect 122742 34552 122748 34604
rect 122800 34592 122806 34604
rect 172514 34592 172520 34604
rect 122800 34564 172520 34592
rect 122800 34552 122806 34564
rect 172514 34552 172520 34564
rect 172572 34552 172578 34604
rect 176562 34552 176568 34604
rect 176620 34592 176626 34604
rect 226334 34592 226340 34604
rect 176620 34564 226340 34592
rect 176620 34552 176626 34564
rect 226334 34552 226340 34564
rect 226392 34552 226398 34604
rect 230382 34552 230388 34604
rect 230440 34592 230446 34604
rect 280154 34592 280160 34604
rect 230440 34564 280160 34592
rect 230440 34552 230446 34564
rect 280154 34552 280160 34564
rect 280212 34552 280218 34604
rect 284202 34552 284208 34604
rect 284260 34592 284266 34604
rect 335354 34592 335360 34604
rect 284260 34564 335360 34592
rect 284260 34552 284266 34564
rect 335354 34552 335360 34564
rect 335412 34552 335418 34604
rect 365622 34552 365628 34604
rect 365680 34592 365686 34604
rect 415394 34592 415400 34604
rect 365680 34564 415400 34592
rect 365680 34552 365686 34564
rect 415394 34552 415400 34564
rect 415452 34552 415458 34604
rect 419442 34552 419448 34604
rect 419500 34592 419506 34604
rect 469214 34592 469220 34604
rect 419500 34564 469220 34592
rect 419500 34552 419506 34564
rect 469214 34552 469220 34564
rect 469272 34552 469278 34604
rect 473262 34552 473268 34604
rect 473320 34592 473326 34604
rect 523034 34592 523040 34604
rect 473320 34564 523040 34592
rect 473320 34552 473326 34564
rect 523034 34552 523040 34564
rect 523092 34552 523098 34604
rect 13722 34484 13728 34536
rect 13780 34524 13786 34536
rect 64874 34524 64880 34536
rect 13780 34496 64880 34524
rect 13780 34484 13786 34496
rect 64874 34484 64880 34496
rect 64932 34484 64938 34536
rect 95142 34484 95148 34536
rect 95200 34524 95206 34536
rect 146294 34524 146300 34536
rect 95200 34496 146300 34524
rect 95200 34484 95206 34496
rect 146294 34484 146300 34496
rect 146352 34484 146358 34536
rect 148962 34484 148968 34536
rect 149020 34524 149026 34536
rect 200114 34524 200120 34536
rect 149020 34496 200120 34524
rect 149020 34484 149026 34496
rect 200114 34484 200120 34496
rect 200172 34484 200178 34536
rect 202782 34484 202788 34536
rect 202840 34524 202846 34536
rect 253934 34524 253940 34536
rect 202840 34496 253940 34524
rect 202840 34484 202846 34496
rect 253934 34484 253940 34496
rect 253992 34484 253998 34536
rect 256602 34484 256608 34536
rect 256660 34524 256666 34536
rect 307754 34524 307760 34536
rect 256660 34496 307760 34524
rect 256660 34484 256666 34496
rect 307754 34484 307760 34496
rect 307812 34484 307818 34536
rect 338022 34484 338028 34536
rect 338080 34524 338086 34536
rect 389174 34524 389180 34536
rect 338080 34496 389180 34524
rect 338080 34484 338086 34496
rect 389174 34484 389180 34496
rect 389232 34484 389238 34536
rect 391842 34484 391848 34536
rect 391900 34524 391906 34536
rect 442994 34524 443000 34536
rect 391900 34496 443000 34524
rect 391900 34484 391906 34496
rect 442994 34484 443000 34496
rect 443052 34484 443058 34536
rect 445662 34484 445668 34536
rect 445720 34524 445726 34536
rect 496814 34524 496820 34536
rect 445720 34496 496820 34524
rect 445720 34484 445726 34496
rect 496814 34484 496820 34496
rect 496872 34484 496878 34536
rect 500862 34484 500868 34536
rect 500920 34524 500926 34536
rect 550634 34524 550640 34536
rect 500920 34496 550640 34524
rect 500920 34484 500926 34496
rect 550634 34484 550640 34496
rect 550692 34484 550698 34536
rect 35618 16532 35624 16584
rect 35676 16572 35682 16584
rect 36630 16572 36636 16584
rect 35676 16544 36636 16572
rect 35676 16532 35682 16544
rect 36630 16532 36636 16544
rect 36688 16532 36694 16584
rect 200758 16532 200764 16584
rect 200816 16572 200822 16584
rect 204622 16572 204628 16584
rect 200816 16544 204628 16572
rect 200816 16532 200822 16544
rect 204622 16532 204628 16544
rect 204680 16532 204686 16584
rect 332502 16532 332508 16584
rect 332560 16572 332566 16584
rect 335998 16572 336004 16584
rect 332560 16544 336004 16572
rect 332560 16532 332566 16544
rect 335998 16532 336004 16544
rect 336056 16532 336062 16584
rect 446398 16532 446404 16584
rect 446456 16572 446462 16584
rect 447686 16572 447692 16584
rect 446456 16544 447692 16572
rect 446456 16532 446462 16544
rect 447686 16532 447692 16544
rect 447744 16532 447750 16584
rect 521746 16532 521752 16584
rect 521804 16572 521810 16584
rect 522390 16572 522396 16584
rect 521804 16544 522396 16572
rect 521804 16532 521810 16544
rect 522390 16532 522396 16544
rect 522448 16532 522454 16584
rect 144886 13824 154574 13852
rect 62758 13744 62764 13796
rect 62816 13784 62822 13796
rect 69750 13784 69756 13796
rect 62816 13756 69756 13784
rect 62816 13744 62822 13756
rect 69750 13744 69756 13756
rect 69808 13744 69814 13796
rect 36538 13676 36544 13728
rect 36596 13716 36602 13728
rect 144886 13716 144914 13824
rect 154546 13784 154574 13824
rect 154546 13756 157334 13784
rect 36596 13688 144914 13716
rect 36596 13676 36602 13688
rect 146938 13676 146944 13728
rect 146996 13716 147002 13728
rect 157306 13716 157334 13756
rect 251818 13744 251824 13796
rect 251876 13784 251882 13796
rect 258718 13784 258724 13796
rect 251876 13756 258724 13784
rect 251876 13744 251882 13756
rect 258718 13744 258724 13756
rect 258776 13744 258782 13796
rect 350074 13744 350080 13796
rect 350132 13784 350138 13796
rect 359550 13784 359556 13796
rect 350132 13756 359556 13784
rect 350132 13744 350138 13756
rect 359550 13744 359556 13756
rect 359608 13744 359614 13796
rect 494698 13744 494704 13796
rect 494756 13784 494762 13796
rect 501598 13784 501604 13796
rect 494756 13756 501604 13784
rect 494756 13744 494762 13756
rect 501598 13744 501604 13756
rect 501656 13744 501662 13796
rect 538398 13716 538404 13728
rect 146996 13688 150848 13716
rect 157306 13688 538404 13716
rect 146996 13676 147002 13688
rect 15194 13608 15200 13660
rect 15252 13648 15258 13660
rect 42794 13648 42800 13660
rect 15252 13620 42800 13648
rect 15252 13608 15258 13620
rect 42794 13608 42800 13620
rect 42852 13608 42858 13660
rect 53098 13608 53104 13660
rect 53156 13648 53162 13660
rect 64138 13648 64144 13660
rect 53156 13620 64144 13648
rect 53156 13608 53162 13620
rect 64138 13608 64144 13620
rect 64196 13608 64202 13660
rect 69106 13608 69112 13660
rect 69164 13648 69170 13660
rect 96798 13648 96804 13660
rect 69164 13620 96804 13648
rect 69164 13608 69170 13620
rect 96798 13608 96804 13620
rect 96856 13608 96862 13660
rect 123662 13648 123668 13660
rect 103486 13620 123668 13648
rect 25958 13540 25964 13592
rect 26016 13580 26022 13592
rect 36722 13580 36728 13592
rect 26016 13552 36728 13580
rect 26016 13540 26022 13552
rect 36722 13540 36728 13552
rect 36780 13540 36786 13592
rect 79962 13540 79968 13592
rect 80020 13580 80026 13592
rect 90450 13580 90456 13592
rect 80020 13552 90456 13580
rect 80020 13540 80026 13552
rect 90450 13540 90456 13552
rect 90508 13540 90514 13592
rect 96706 13540 96712 13592
rect 96764 13580 96770 13592
rect 103486 13580 103514 13620
rect 123662 13608 123668 13620
rect 123720 13608 123726 13660
rect 133782 13608 133788 13660
rect 133840 13648 133846 13660
rect 144270 13648 144276 13660
rect 133840 13620 144276 13648
rect 133840 13608 133846 13620
rect 144270 13608 144276 13620
rect 144328 13608 144334 13660
rect 150710 13648 150716 13660
rect 146588 13620 150716 13648
rect 96764 13552 103514 13580
rect 96764 13540 96770 13552
rect 106550 13540 106556 13592
rect 106608 13580 106614 13592
rect 116578 13580 116584 13592
rect 106608 13552 116584 13580
rect 106608 13540 106614 13552
rect 116578 13540 116584 13552
rect 116636 13540 116642 13592
rect 122926 13540 122932 13592
rect 122984 13580 122990 13592
rect 146588 13580 146616 13620
rect 150710 13608 150716 13620
rect 150768 13608 150774 13660
rect 150820 13648 150848 13688
rect 538398 13676 538404 13688
rect 538456 13676 538462 13728
rect 548058 13648 548064 13660
rect 150820 13620 548064 13648
rect 548058 13608 548064 13620
rect 548116 13608 548122 13660
rect 122984 13552 146616 13580
rect 122984 13540 122990 13552
rect 150526 13540 150532 13592
rect 150584 13580 150590 13592
rect 178126 13580 178132 13592
rect 150584 13552 178132 13580
rect 150584 13540 150590 13552
rect 178126 13540 178132 13552
rect 178184 13540 178190 13592
rect 187970 13540 187976 13592
rect 188028 13580 188034 13592
rect 199378 13580 199384 13592
rect 188028 13552 199384 13580
rect 188028 13540 188034 13552
rect 199378 13540 199384 13552
rect 199436 13540 199442 13592
rect 204346 13540 204352 13592
rect 204404 13580 204410 13592
rect 231854 13580 231860 13592
rect 204404 13552 231860 13580
rect 204404 13540 204410 13552
rect 231854 13540 231860 13552
rect 231912 13540 231918 13592
rect 242066 13540 242072 13592
rect 242124 13580 242130 13592
rect 253198 13580 253204 13592
rect 242124 13552 253204 13580
rect 242124 13540 242130 13552
rect 253198 13540 253204 13552
rect 253256 13540 253262 13592
rect 258166 13540 258172 13592
rect 258224 13580 258230 13592
rect 258224 13552 281764 13580
rect 258224 13540 258230 13552
rect 160554 13472 160560 13524
rect 160612 13512 160618 13524
rect 171778 13512 171784 13524
rect 160612 13484 171784 13512
rect 160612 13472 160618 13484
rect 171778 13472 171784 13484
rect 171836 13472 171842 13524
rect 215018 13472 215024 13524
rect 215076 13512 215082 13524
rect 225598 13512 225604 13524
rect 215076 13484 225604 13512
rect 215076 13472 215082 13484
rect 225598 13472 225604 13484
rect 225656 13472 225662 13524
rect 268930 13472 268936 13524
rect 268988 13512 268994 13524
rect 279510 13512 279516 13524
rect 268988 13484 279516 13512
rect 268988 13472 268994 13484
rect 279510 13472 279516 13484
rect 279568 13472 279574 13524
rect 281736 13512 281764 13552
rect 285766 13540 285772 13592
rect 285824 13580 285830 13592
rect 312630 13580 312636 13592
rect 285824 13552 312636 13580
rect 285824 13540 285830 13552
rect 312630 13540 312636 13552
rect 312688 13540 312694 13592
rect 340138 13580 340144 13592
rect 316006 13552 340144 13580
rect 286134 13512 286140 13524
rect 281736 13484 286140 13512
rect 286134 13472 286140 13484
rect 286192 13472 286198 13524
rect 295978 13472 295984 13524
rect 296036 13512 296042 13524
rect 307018 13512 307024 13524
rect 296036 13484 307024 13512
rect 296036 13472 296042 13484
rect 307018 13472 307024 13484
rect 307076 13472 307082 13524
rect 311986 13472 311992 13524
rect 312044 13512 312050 13524
rect 316006 13512 316034 13552
rect 340138 13540 340144 13552
rect 340196 13540 340202 13592
rect 344986 13552 354674 13580
rect 312044 13484 316034 13512
rect 312044 13472 312050 13484
rect 322842 13472 322848 13524
rect 322900 13512 322906 13524
rect 333238 13512 333244 13524
rect 322900 13484 333244 13512
rect 322900 13472 322906 13484
rect 333238 13472 333244 13484
rect 333296 13472 333302 13524
rect 339586 13472 339592 13524
rect 339644 13512 339650 13524
rect 344986 13512 345014 13552
rect 339644 13484 345014 13512
rect 354646 13512 354674 13552
rect 365806 13540 365812 13592
rect 365864 13580 365870 13592
rect 393590 13580 393596 13592
rect 365864 13552 393596 13580
rect 365864 13540 365870 13552
rect 393590 13540 393596 13552
rect 393648 13540 393654 13592
rect 420914 13580 420920 13592
rect 402946 13552 420920 13580
rect 366726 13512 366732 13524
rect 354646 13484 366732 13512
rect 339644 13472 339650 13484
rect 366726 13472 366732 13484
rect 366784 13472 366790 13524
rect 376570 13472 376576 13524
rect 376628 13512 376634 13524
rect 387058 13512 387064 13524
rect 376628 13484 387064 13512
rect 376628 13472 376634 13484
rect 387058 13472 387064 13484
rect 387116 13472 387122 13524
rect 393406 13472 393412 13524
rect 393464 13512 393470 13524
rect 402946 13512 402974 13552
rect 420914 13540 420920 13552
rect 420972 13540 420978 13592
rect 431034 13540 431040 13592
rect 431092 13580 431098 13592
rect 442258 13580 442264 13592
rect 431092 13552 442264 13580
rect 431092 13540 431098 13552
rect 442258 13540 442264 13552
rect 442316 13540 442322 13592
rect 447226 13540 447232 13592
rect 447284 13580 447290 13592
rect 474734 13580 474740 13592
rect 447284 13552 474740 13580
rect 447284 13540 447290 13552
rect 474734 13540 474740 13552
rect 474792 13540 474798 13592
rect 484946 13540 484952 13592
rect 485004 13580 485010 13592
rect 496078 13580 496084 13592
rect 485004 13552 496084 13580
rect 485004 13540 485010 13552
rect 496078 13540 496084 13552
rect 496136 13540 496142 13592
rect 501046 13540 501052 13592
rect 501104 13580 501110 13592
rect 528738 13580 528744 13592
rect 501104 13552 528744 13580
rect 501104 13540 501110 13552
rect 528738 13540 528744 13552
rect 528796 13540 528802 13592
rect 393464 13484 402974 13512
rect 393464 13472 393470 13484
rect 403986 13472 403992 13524
rect 404044 13512 404050 13524
rect 414658 13512 414664 13524
rect 404044 13484 414664 13512
rect 404044 13472 404050 13484
rect 414658 13472 414664 13484
rect 414716 13472 414722 13524
rect 458082 13472 458088 13524
rect 458140 13512 458146 13524
rect 468570 13512 468576 13524
rect 458140 13484 468576 13512
rect 458140 13472 458146 13484
rect 468570 13472 468576 13484
rect 468628 13472 468634 13524
rect 511902 13472 511908 13524
rect 511960 13512 511966 13524
rect 522298 13512 522304 13524
rect 511960 13484 522304 13512
rect 511960 13472 511966 13484
rect 522298 13472 522304 13484
rect 522356 13472 522362 13524
rect 16298 13404 16304 13456
rect 16356 13444 16362 13456
rect 580258 13444 580264 13456
rect 16356 13416 580264 13444
rect 16356 13404 16362 13416
rect 580258 13404 580264 13416
rect 580316 13404 580322 13456
<< via1 >>
rect 25964 686128 26016 686180
rect 149704 686128 149756 686180
rect 36636 686060 36688 686112
rect 52460 686060 52512 686112
rect 232320 686060 232372 686112
rect 251824 686060 251876 686112
rect 62488 685992 62540 686044
rect 79324 685992 79376 686044
rect 90364 685992 90416 686044
rect 106372 685992 106424 686044
rect 116492 685992 116544 686044
rect 133420 685992 133472 686044
rect 144276 685992 144328 686044
rect 160284 685992 160336 686044
rect 170496 685992 170548 686044
rect 187792 685992 187844 686044
rect 197544 685992 197596 686044
rect 214380 685992 214432 686044
rect 224500 685992 224552 686044
rect 241520 685992 241572 686044
rect 413468 685992 413520 686044
rect 430580 685992 430632 686044
rect 440516 685992 440568 686044
rect 457260 685992 457312 686044
rect 468576 685992 468628 686044
rect 484400 685992 484452 686044
rect 494520 685992 494572 686044
rect 511356 685992 511408 686044
rect 36728 685924 36780 685976
rect 62120 685924 62172 685976
rect 64144 685924 64196 685976
rect 89076 685924 89128 685976
rect 90456 685924 90508 685976
rect 115940 685924 115992 685976
rect 116584 685924 116636 685976
rect 142988 685924 143040 685976
rect 144184 685924 144236 685976
rect 170036 685924 170088 685976
rect 178408 685924 178460 685976
rect 200764 685924 200816 685976
rect 251456 685924 251508 685976
rect 268292 685924 268344 685976
rect 279424 685924 279476 685976
rect 295800 685924 295852 685976
rect 305552 685924 305604 685976
rect 322388 685924 322440 685976
rect 334624 685924 334676 685976
rect 349804 685924 349856 685976
rect 359648 685924 359700 685976
rect 376300 685924 376352 685976
rect 386512 685924 386564 685976
rect 403348 685924 403400 685976
rect 421288 685924 421340 685976
rect 443644 685924 443696 685976
rect 475384 685924 475436 685976
rect 494704 685924 494756 685976
rect 522396 685924 522448 685976
rect 538404 685924 538456 685976
rect 43352 685856 43404 685908
rect 62764 685856 62816 685908
rect 171784 685856 171836 685908
rect 197452 685856 197504 685908
rect 199384 685856 199436 685908
rect 223948 685856 224000 685908
rect 225604 685856 225656 685908
rect 251180 685856 251232 685908
rect 253204 685856 253256 685908
rect 278044 685856 278096 685908
rect 279516 685856 279568 685908
rect 305460 685856 305512 685908
rect 307024 685856 307076 685908
rect 331956 685856 332008 685908
rect 333244 685856 333296 685908
rect 359464 685856 359516 685908
rect 359740 685856 359792 685908
rect 386052 685856 386104 685908
rect 387064 685856 387116 685908
rect 412916 685856 412968 685908
rect 414664 685856 414716 685908
rect 440240 685856 440292 685908
rect 442264 685856 442316 685908
rect 467012 685856 467064 685908
rect 468484 685856 468536 685908
rect 494060 685856 494112 685908
rect 496084 685856 496136 685908
rect 520924 685856 520976 685908
rect 522304 685856 522356 685908
rect 548064 685856 548116 685908
rect 285772 683272 285824 683324
rect 286140 683272 286192 683324
rect 339592 683272 339644 683324
rect 340144 683272 340196 683324
rect 68928 683204 68980 683256
rect 118700 683204 118752 683256
rect 122748 683204 122800 683256
rect 172520 683204 172572 683256
rect 230388 683204 230440 683256
rect 280160 683204 280212 683256
rect 311808 683204 311860 683256
rect 361580 683204 361632 683256
rect 500868 683204 500920 683256
rect 550640 683204 550692 683256
rect 41328 683136 41380 683188
rect 91100 683136 91152 683188
rect 148968 683136 149020 683188
rect 200120 683136 200172 683188
rect 202788 683136 202840 683188
rect 253940 683136 253992 683188
rect 284208 683136 284260 683188
rect 335360 683136 335412 683188
rect 365628 683136 365680 683188
rect 415400 683136 415452 683188
rect 419448 683136 419500 683188
rect 469220 683136 469272 683188
rect 473268 683136 473320 683188
rect 523040 683136 523092 683188
rect 143632 666136 143684 666188
rect 144276 666136 144328 666188
rect 13728 665116 13780 665168
rect 64880 665116 64932 665168
rect 95148 665116 95200 665168
rect 146300 665116 146352 665168
rect 176568 665116 176620 665168
rect 226340 665116 226392 665168
rect 256608 665116 256660 665168
rect 307760 665116 307812 665168
rect 332508 665116 332560 665168
rect 334624 665116 334676 665168
rect 338028 665116 338080 665168
rect 389180 665116 389232 665168
rect 391848 665116 391900 665168
rect 443000 665116 443052 665168
rect 445668 665116 445720 665168
rect 496820 665116 496872 665168
rect 35624 665048 35676 665100
rect 36636 665048 36688 665100
rect 467656 665048 467708 665100
rect 468576 665048 468628 665100
rect 521384 663688 521436 663740
rect 522396 663688 522448 663740
rect 62764 662328 62816 662380
rect 70032 662328 70084 662380
rect 96712 662328 96764 662380
rect 124036 662328 124088 662380
rect 150532 662328 150584 662380
rect 178040 662328 178092 662380
rect 187700 662328 187752 662380
rect 199384 662328 199436 662380
rect 200764 662328 200816 662380
rect 204996 662328 205048 662380
rect 25688 662260 25740 662312
rect 36728 662260 36780 662312
rect 53104 662260 53156 662312
rect 64144 662260 64196 662312
rect 79692 662260 79744 662312
rect 90456 662260 90508 662312
rect 106648 662260 106700 662312
rect 116584 662260 116636 662312
rect 133696 662260 133748 662312
rect 144184 662260 144236 662312
rect 160652 662260 160704 662312
rect 171784 662260 171836 662312
rect 204352 662260 204404 662312
rect 232044 662328 232096 662380
rect 251824 662328 251876 662380
rect 259000 662328 259052 662380
rect 285772 662328 285824 662380
rect 313004 662328 313056 662380
rect 339592 662328 339644 662380
rect 366732 662328 366784 662380
rect 214656 662260 214708 662312
rect 225604 662260 225656 662312
rect 241704 662260 241756 662312
rect 253204 662260 253256 662312
rect 268660 662260 268712 662312
rect 279516 662260 279568 662312
rect 295708 662260 295760 662312
rect 307024 662260 307076 662312
rect 322664 662260 322716 662312
rect 333244 662260 333296 662312
rect 349712 662260 349764 662312
rect 359556 662260 359608 662312
rect 365812 662260 365864 662312
rect 393596 662328 393648 662380
rect 376668 662260 376720 662312
rect 387064 662260 387116 662312
rect 393412 662260 393464 662312
rect 421012 662328 421064 662380
rect 430672 662328 430724 662380
rect 442264 662328 442316 662380
rect 443644 662328 443696 662380
rect 447692 662328 447744 662380
rect 494704 662328 494756 662380
rect 501972 662328 502024 662380
rect 403716 662260 403768 662312
rect 414664 662260 414716 662312
rect 457720 662260 457772 662312
rect 468484 662260 468536 662312
rect 484676 662260 484728 662312
rect 496084 662260 496136 662312
rect 511724 662260 511776 662312
rect 522304 662260 522356 662312
rect 15200 662192 15252 662244
rect 42984 662192 43036 662244
rect 69112 662192 69164 662244
rect 96988 662192 97040 662244
rect 122932 662192 122984 662244
rect 150992 662192 151044 662244
rect 258172 662192 258224 662244
rect 286048 662192 286100 662244
rect 311992 662192 312044 662244
rect 340052 662192 340104 662244
rect 447232 662192 447284 662244
rect 475016 662192 475068 662244
rect 501052 662192 501104 662244
rect 529020 662192 529072 662244
rect 16028 658928 16080 658980
rect 529020 658928 529072 658980
rect 25688 658520 25740 658572
rect 146944 658520 146996 658572
rect 36728 658452 36780 658504
rect 52644 658452 52696 658504
rect 232044 658452 232096 658504
rect 251824 658452 251876 658504
rect 475016 658452 475068 658504
rect 494704 658452 494756 658504
rect 62488 658384 62540 658436
rect 79692 658384 79744 658436
rect 90456 658384 90508 658436
rect 106648 658384 106700 658436
rect 116492 658384 116544 658436
rect 133696 658384 133748 658436
rect 170496 658384 170548 658436
rect 187700 658384 187752 658436
rect 197452 658384 197504 658436
rect 214656 658384 214708 658436
rect 224500 658384 224552 658436
rect 241704 658384 241756 658436
rect 413468 658384 413520 658436
rect 430672 658384 430724 658436
rect 440516 658384 440568 658436
rect 457628 658384 457680 658436
rect 468484 658384 468536 658436
rect 484676 658384 484728 658436
rect 36820 658316 36872 658368
rect 62304 658316 62356 658368
rect 64144 658316 64196 658368
rect 89352 658316 89404 658368
rect 90364 658316 90416 658368
rect 116308 658316 116360 658368
rect 116584 658316 116636 658368
rect 143356 658316 143408 658368
rect 144276 658316 144328 658368
rect 170312 658316 170364 658368
rect 178040 658316 178092 658368
rect 200764 658316 200816 658368
rect 251456 658316 251508 658368
rect 268660 658316 268712 658368
rect 279424 658316 279476 658368
rect 295708 658316 295760 658368
rect 305460 658316 305512 658368
rect 322664 658316 322716 658368
rect 336004 658316 336056 658368
rect 349712 658316 349764 658368
rect 359464 658316 359516 658368
rect 376668 658316 376720 658368
rect 386512 658316 386564 658368
rect 403624 658316 403676 658368
rect 421012 658316 421064 658368
rect 446404 658316 446456 658368
rect 494520 658316 494572 658368
rect 511632 658316 511684 658368
rect 522304 658316 522356 658368
rect 538680 658316 538732 658368
rect 43076 658248 43128 658300
rect 62764 658248 62816 658300
rect 144184 658248 144236 658300
rect 160652 658248 160704 658300
rect 171784 658248 171836 658300
rect 197360 658248 197412 658300
rect 199384 658248 199436 658300
rect 224316 658248 224368 658300
rect 225604 658248 225656 658300
rect 251364 658248 251416 658300
rect 253204 658248 253256 658300
rect 278320 658248 278372 658300
rect 279516 658248 279568 658300
rect 305368 658248 305420 658300
rect 307024 658248 307076 658300
rect 332324 658248 332376 658300
rect 333244 658248 333296 658300
rect 359372 658248 359424 658300
rect 359556 658248 359608 658300
rect 386328 658248 386380 658300
rect 387064 658248 387116 658300
rect 413284 658248 413336 658300
rect 414664 658248 414716 658300
rect 440332 658248 440384 658300
rect 442264 658248 442316 658300
rect 467288 658248 467340 658300
rect 468576 658248 468628 658300
rect 494336 658248 494388 658300
rect 496084 658248 496136 658300
rect 521292 658248 521344 658300
rect 522396 658248 522448 658300
rect 548340 658248 548392 658300
rect 37924 657500 37976 657552
rect 526444 657500 526496 657552
rect 35624 656888 35676 656940
rect 36636 656888 36688 656940
rect 68928 655664 68980 655716
rect 118700 655664 118752 655716
rect 311808 655664 311860 655716
rect 361580 655664 361632 655716
rect 41328 655596 41380 655648
rect 91100 655596 91152 655648
rect 122748 655596 122800 655648
rect 172520 655596 172572 655648
rect 176568 655596 176620 655648
rect 226340 655596 226392 655648
rect 230388 655596 230440 655648
rect 280160 655596 280212 655648
rect 284208 655596 284260 655648
rect 335360 655596 335412 655648
rect 365628 655596 365680 655648
rect 415400 655596 415452 655648
rect 419448 655596 419500 655648
rect 469220 655596 469272 655648
rect 473268 655596 473320 655648
rect 523040 655596 523092 655648
rect 13728 655528 13780 655580
rect 64880 655528 64932 655580
rect 96620 655528 96672 655580
rect 146300 655528 146352 655580
rect 148968 655528 149020 655580
rect 200120 655528 200172 655580
rect 202788 655528 202840 655580
rect 253940 655528 253992 655580
rect 256608 655528 256660 655580
rect 307760 655528 307812 655580
rect 338028 655528 338080 655580
rect 389180 655528 389232 655580
rect 391848 655528 391900 655580
rect 443000 655528 443052 655580
rect 445668 655528 445720 655580
rect 496820 655528 496872 655580
rect 500868 655528 500920 655580
rect 550640 655528 550692 655580
rect 95148 654032 95200 654084
rect 96620 654032 96672 654084
rect 35624 637508 35676 637560
rect 36728 637508 36780 637560
rect 89720 637508 89772 637560
rect 90456 637508 90508 637560
rect 332600 637508 332652 637560
rect 336004 637508 336056 637560
rect 446404 637508 446456 637560
rect 447692 637508 447744 637560
rect 62764 634720 62816 634772
rect 69756 634720 69808 634772
rect 96712 634720 96764 634772
rect 15200 634652 15252 634704
rect 42800 634652 42852 634704
rect 53104 634652 53156 634704
rect 64144 634652 64196 634704
rect 69112 634652 69164 634704
rect 96804 634652 96856 634704
rect 200764 634720 200816 634772
rect 204628 634720 204680 634772
rect 251824 634720 251876 634772
rect 258724 634720 258776 634772
rect 494704 634720 494756 634772
rect 501604 634720 501656 634772
rect 521476 634720 521528 634772
rect 522304 634720 522356 634772
rect 123668 634652 123720 634704
rect 149704 634652 149756 634704
rect 547972 634652 548024 634704
rect 26056 634584 26108 634636
rect 36820 634584 36872 634636
rect 79968 634584 80020 634636
rect 90364 634584 90416 634636
rect 106556 634584 106608 634636
rect 116584 634584 116636 634636
rect 133788 634584 133840 634636
rect 144276 634584 144328 634636
rect 150532 634584 150584 634636
rect 178132 634584 178184 634636
rect 187976 634584 188028 634636
rect 199384 634584 199436 634636
rect 204352 634584 204404 634636
rect 231952 634584 232004 634636
rect 242072 634584 242124 634636
rect 253204 634584 253256 634636
rect 258172 634584 258224 634636
rect 122932 634516 122984 634568
rect 150716 634516 150768 634568
rect 160560 634516 160612 634568
rect 171784 634516 171836 634568
rect 215024 634516 215076 634568
rect 225604 634516 225656 634568
rect 268936 634516 268988 634568
rect 279516 634516 279568 634568
rect 285772 634584 285824 634636
rect 312636 634584 312688 634636
rect 286140 634516 286192 634568
rect 295984 634516 296036 634568
rect 307024 634516 307076 634568
rect 311992 634516 312044 634568
rect 340144 634584 340196 634636
rect 322848 634516 322900 634568
rect 333244 634516 333296 634568
rect 339592 634516 339644 634568
rect 366732 634584 366784 634636
rect 350080 634516 350132 634568
rect 359556 634516 359608 634568
rect 365812 634516 365864 634568
rect 393596 634584 393648 634636
rect 376576 634516 376628 634568
rect 387064 634516 387116 634568
rect 393412 634516 393464 634568
rect 420920 634584 420972 634636
rect 431040 634584 431092 634636
rect 442264 634584 442316 634636
rect 447232 634584 447284 634636
rect 474740 634584 474792 634636
rect 484952 634584 485004 634636
rect 496084 634584 496136 634636
rect 501052 634584 501104 634636
rect 528652 634584 528704 634636
rect 403992 634516 404044 634568
rect 414664 634516 414716 634568
rect 458088 634516 458140 634568
rect 468576 634516 468628 634568
rect 511816 634516 511868 634568
rect 522396 634516 522448 634568
rect 36544 634448 36596 634500
rect 538404 634448 538456 634500
rect 16304 632680 16356 632732
rect 528744 632680 528796 632732
rect 25964 632340 26016 632392
rect 148324 632340 148376 632392
rect 36728 632272 36780 632324
rect 52460 632272 52512 632324
rect 232320 632272 232372 632324
rect 251824 632272 251876 632324
rect 475384 632272 475436 632324
rect 494704 632272 494756 632324
rect 62488 632204 62540 632256
rect 79324 632204 79376 632256
rect 90364 632204 90416 632256
rect 106372 632204 106424 632256
rect 116492 632204 116544 632256
rect 133420 632204 133472 632256
rect 170496 632204 170548 632256
rect 187792 632204 187844 632256
rect 197544 632204 197596 632256
rect 214380 632204 214432 632256
rect 224500 632204 224552 632256
rect 241520 632204 241572 632256
rect 413468 632204 413520 632256
rect 430580 632204 430632 632256
rect 440516 632204 440568 632256
rect 457260 632204 457312 632256
rect 468576 632204 468628 632256
rect 484400 632204 484452 632256
rect 36820 632136 36872 632188
rect 62120 632136 62172 632188
rect 64144 632136 64196 632188
rect 89076 632136 89128 632188
rect 90456 632136 90508 632188
rect 115940 632136 115992 632188
rect 116584 632136 116636 632188
rect 142988 632136 143040 632188
rect 144276 632136 144328 632188
rect 170036 632136 170088 632188
rect 178408 632136 178460 632188
rect 200764 632136 200816 632188
rect 251456 632136 251508 632188
rect 268292 632136 268344 632188
rect 279424 632136 279476 632188
rect 295800 632136 295852 632188
rect 305644 632136 305696 632188
rect 322388 632136 322440 632188
rect 336004 632136 336056 632188
rect 349804 632136 349856 632188
rect 359556 632136 359608 632188
rect 376300 632136 376352 632188
rect 386512 632136 386564 632188
rect 403348 632136 403400 632188
rect 421288 632136 421340 632188
rect 445024 632136 445076 632188
rect 494520 632136 494572 632188
rect 511356 632136 511408 632188
rect 522304 632136 522356 632188
rect 538404 632136 538456 632188
rect 43352 632068 43404 632120
rect 62764 632068 62816 632120
rect 144184 632068 144236 632120
rect 160284 632068 160336 632120
rect 171784 632068 171836 632120
rect 197452 632068 197504 632120
rect 199384 632068 199436 632120
rect 223948 632068 224000 632120
rect 225604 632068 225656 632120
rect 251180 632068 251232 632120
rect 253204 632068 253256 632120
rect 278044 632068 278096 632120
rect 279516 632068 279568 632120
rect 305552 632068 305604 632120
rect 307024 632068 307076 632120
rect 331956 632068 332008 632120
rect 333244 632068 333296 632120
rect 359464 632068 359516 632120
rect 359740 632068 359792 632120
rect 386052 632068 386104 632120
rect 387064 632068 387116 632120
rect 413008 632068 413060 632120
rect 414664 632068 414716 632120
rect 440240 632068 440292 632120
rect 442264 632068 442316 632120
rect 467012 632068 467064 632120
rect 468484 632068 468536 632120
rect 494060 632068 494112 632120
rect 496084 632068 496136 632120
rect 520924 632068 520976 632120
rect 522396 632068 522448 632120
rect 548064 632068 548116 632120
rect 37924 629892 37976 629944
rect 526444 629892 526496 629944
rect 285772 629280 285824 629332
rect 286140 629280 286192 629332
rect 339592 629280 339644 629332
rect 340144 629280 340196 629332
rect 13728 611260 13780 611312
rect 64880 611260 64932 611312
rect 95148 611260 95200 611312
rect 146300 611260 146352 611312
rect 148968 611260 149020 611312
rect 200120 611260 200172 611312
rect 202788 611260 202840 611312
rect 253940 611260 253992 611312
rect 256608 611260 256660 611312
rect 307760 611260 307812 611312
rect 338028 611260 338080 611312
rect 389180 611260 389232 611312
rect 391848 611260 391900 611312
rect 443000 611260 443052 611312
rect 445668 611260 445720 611312
rect 496820 611260 496872 611312
rect 500868 611260 500920 611312
rect 550640 611260 550692 611312
rect 35624 611192 35676 611244
rect 36728 611192 36780 611244
rect 41328 611192 41380 611244
rect 91100 611192 91152 611244
rect 122748 611192 122800 611244
rect 172520 611192 172572 611244
rect 176568 611192 176620 611244
rect 226340 611192 226392 611244
rect 230388 611192 230440 611244
rect 280160 611192 280212 611244
rect 284208 611192 284260 611244
rect 335360 611192 335412 611244
rect 365628 611192 365680 611244
rect 415400 611192 415452 611244
rect 419448 611192 419500 611244
rect 469220 611192 469272 611244
rect 473268 611192 473320 611244
rect 523040 611192 523092 611244
rect 68928 611124 68980 611176
rect 118700 611124 118752 611176
rect 311808 611124 311860 611176
rect 361580 611124 361632 611176
rect 445024 611124 445076 611176
rect 447692 611124 447744 611176
rect 467656 611124 467708 611176
rect 468576 611124 468628 611176
rect 332600 610648 332652 610700
rect 336004 610648 336056 610700
rect 52736 608540 52788 608592
rect 64144 608540 64196 608592
rect 69112 608540 69164 608592
rect 15200 608472 15252 608524
rect 42984 608472 43036 608524
rect 62764 608472 62816 608524
rect 70032 608472 70084 608524
rect 96712 608540 96764 608592
rect 96988 608472 97040 608524
rect 146944 608540 146996 608592
rect 124036 608472 124088 608524
rect 133696 608472 133748 608524
rect 144276 608472 144328 608524
rect 150532 608472 150584 608524
rect 200764 608540 200816 608592
rect 204996 608540 205048 608592
rect 251824 608540 251876 608592
rect 259000 608540 259052 608592
rect 494704 608540 494756 608592
rect 501972 608540 502024 608592
rect 25688 608404 25740 608456
rect 36820 608404 36872 608456
rect 79692 608404 79744 608456
rect 90456 608404 90508 608456
rect 106648 608404 106700 608456
rect 116584 608404 116636 608456
rect 122932 608404 122984 608456
rect 150992 608404 151044 608456
rect 548340 608472 548392 608524
rect 178040 608404 178092 608456
rect 187700 608404 187752 608456
rect 199384 608404 199436 608456
rect 204352 608404 204404 608456
rect 232044 608404 232096 608456
rect 241704 608404 241756 608456
rect 253204 608404 253256 608456
rect 258172 608404 258224 608456
rect 286048 608404 286100 608456
rect 160652 608336 160704 608388
rect 171784 608336 171836 608388
rect 214656 608336 214708 608388
rect 225604 608336 225656 608388
rect 268660 608336 268712 608388
rect 279516 608336 279568 608388
rect 285772 608336 285824 608388
rect 313004 608404 313056 608456
rect 295708 608336 295760 608388
rect 307024 608336 307076 608388
rect 311992 608336 312044 608388
rect 340052 608404 340104 608456
rect 322664 608336 322716 608388
rect 333244 608336 333296 608388
rect 339592 608336 339644 608388
rect 367008 608404 367060 608456
rect 349712 608336 349764 608388
rect 359556 608336 359608 608388
rect 365812 608336 365864 608388
rect 393964 608404 394016 608456
rect 376668 608336 376720 608388
rect 387064 608336 387116 608388
rect 393412 608336 393464 608388
rect 421012 608404 421064 608456
rect 430672 608404 430724 608456
rect 442264 608404 442316 608456
rect 447232 608404 447284 608456
rect 475016 608404 475068 608456
rect 484676 608404 484728 608456
rect 496084 608404 496136 608456
rect 501052 608404 501104 608456
rect 529020 608404 529072 608456
rect 403716 608336 403768 608388
rect 414664 608336 414716 608388
rect 457720 608336 457772 608388
rect 468484 608336 468536 608388
rect 511724 608336 511776 608388
rect 522396 608336 522448 608388
rect 36636 608268 36688 608320
rect 538680 608268 538732 608320
rect 15292 605072 15344 605124
rect 529020 605072 529072 605124
rect 25688 604732 25740 604784
rect 146944 604732 146996 604784
rect 36728 604664 36780 604716
rect 52644 604664 52696 604716
rect 232044 604664 232096 604716
rect 251824 604664 251876 604716
rect 475016 604664 475068 604716
rect 494704 604664 494756 604716
rect 62488 604596 62540 604648
rect 79692 604596 79744 604648
rect 90456 604596 90508 604648
rect 106648 604596 106700 604648
rect 116492 604596 116544 604648
rect 133696 604596 133748 604648
rect 170496 604596 170548 604648
rect 187700 604596 187752 604648
rect 197452 604596 197504 604648
rect 214656 604596 214708 604648
rect 224500 604596 224552 604648
rect 241704 604596 241756 604648
rect 413468 604596 413520 604648
rect 430672 604596 430724 604648
rect 440516 604596 440568 604648
rect 457628 604596 457680 604648
rect 468576 604596 468628 604648
rect 484676 604596 484728 604648
rect 36820 604528 36872 604580
rect 62304 604528 62356 604580
rect 64144 604528 64196 604580
rect 89352 604528 89404 604580
rect 90364 604528 90416 604580
rect 116308 604528 116360 604580
rect 116584 604528 116636 604580
rect 143356 604528 143408 604580
rect 144276 604528 144328 604580
rect 170312 604528 170364 604580
rect 178040 604528 178092 604580
rect 200764 604528 200816 604580
rect 251456 604528 251508 604580
rect 268660 604528 268712 604580
rect 279516 604528 279568 604580
rect 295708 604528 295760 604580
rect 305460 604528 305512 604580
rect 322664 604528 322716 604580
rect 336004 604528 336056 604580
rect 349712 604528 349764 604580
rect 359464 604528 359516 604580
rect 376668 604528 376720 604580
rect 386512 604528 386564 604580
rect 403624 604528 403676 604580
rect 421012 604528 421064 604580
rect 445024 604528 445076 604580
rect 494520 604528 494572 604580
rect 511632 604528 511684 604580
rect 522304 604528 522356 604580
rect 538680 604528 538732 604580
rect 43076 604460 43128 604512
rect 62764 604460 62816 604512
rect 144184 604460 144236 604512
rect 160652 604460 160704 604512
rect 171784 604460 171836 604512
rect 197360 604460 197412 604512
rect 199384 604460 199436 604512
rect 224316 604460 224368 604512
rect 225604 604460 225656 604512
rect 251364 604460 251416 604512
rect 253204 604460 253256 604512
rect 278320 604460 278372 604512
rect 279424 604460 279476 604512
rect 305368 604460 305420 604512
rect 307024 604460 307076 604512
rect 332324 604460 332376 604512
rect 333244 604460 333296 604512
rect 359372 604460 359424 604512
rect 359556 604460 359608 604512
rect 386328 604460 386380 604512
rect 387064 604460 387116 604512
rect 413284 604460 413336 604512
rect 414664 604460 414716 604512
rect 440332 604460 440384 604512
rect 442264 604460 442316 604512
rect 467288 604460 467340 604512
rect 468484 604460 468536 604512
rect 494336 604460 494388 604512
rect 496084 604460 496136 604512
rect 521292 604460 521344 604512
rect 522396 604460 522448 604512
rect 548340 604460 548392 604512
rect 37924 602352 37976 602404
rect 526444 602352 526496 602404
rect 35624 601672 35676 601724
rect 36636 601672 36688 601724
rect 278780 584740 278832 584792
rect 279516 584740 279568 584792
rect 445024 583720 445076 583772
rect 447692 583720 447744 583772
rect 13728 583652 13780 583704
rect 64880 583652 64932 583704
rect 89720 583652 89772 583704
rect 90456 583652 90508 583704
rect 95148 583652 95200 583704
rect 146300 583652 146352 583704
rect 148968 583652 149020 583704
rect 200120 583652 200172 583704
rect 202788 583652 202840 583704
rect 253940 583652 253992 583704
rect 256608 583652 256660 583704
rect 307760 583652 307812 583704
rect 332600 583652 332652 583704
rect 336004 583652 336056 583704
rect 338028 583652 338080 583704
rect 389180 583652 389232 583704
rect 391848 583652 391900 583704
rect 443000 583652 443052 583704
rect 445668 583652 445720 583704
rect 496820 583652 496872 583704
rect 500868 583652 500920 583704
rect 550640 583652 550692 583704
rect 35624 583584 35676 583636
rect 36728 583584 36780 583636
rect 41328 583584 41380 583636
rect 91100 583584 91152 583636
rect 116216 583584 116268 583636
rect 116492 583584 116544 583636
rect 122748 583584 122800 583636
rect 172520 583584 172572 583636
rect 176568 583584 176620 583636
rect 226340 583584 226392 583636
rect 230388 583584 230440 583636
rect 280160 583584 280212 583636
rect 284208 583584 284260 583636
rect 335360 583584 335412 583636
rect 365628 583584 365680 583636
rect 415400 583584 415452 583636
rect 419448 583584 419500 583636
rect 469220 583584 469272 583636
rect 473268 583584 473320 583636
rect 523040 583584 523092 583636
rect 68928 583516 68980 583568
rect 118700 583516 118752 583568
rect 170220 583516 170272 583568
rect 170496 583516 170548 583568
rect 200764 583516 200816 583568
rect 204628 583516 204680 583568
rect 311808 583516 311860 583568
rect 361580 583516 361632 583568
rect 467656 583516 467708 583568
rect 468576 583516 468628 583568
rect 62764 580932 62816 580984
rect 69756 580932 69808 580984
rect 96712 580932 96764 580984
rect 15200 580864 15252 580916
rect 42800 580864 42852 580916
rect 53104 580864 53156 580916
rect 64144 580864 64196 580916
rect 69112 580864 69164 580916
rect 96804 580864 96856 580916
rect 251824 580932 251876 580984
rect 258724 580932 258776 580984
rect 494704 580932 494756 580984
rect 501604 580932 501656 580984
rect 123668 580864 123720 580916
rect 148324 580864 148376 580916
rect 548064 580864 548116 580916
rect 25964 580796 26016 580848
rect 36820 580796 36872 580848
rect 79968 580796 80020 580848
rect 90364 580796 90416 580848
rect 106556 580796 106608 580848
rect 116584 580796 116636 580848
rect 133788 580796 133840 580848
rect 144276 580796 144328 580848
rect 150532 580796 150584 580848
rect 178132 580796 178184 580848
rect 187976 580796 188028 580848
rect 199384 580796 199436 580848
rect 204352 580796 204404 580848
rect 231860 580796 231912 580848
rect 242072 580796 242124 580848
rect 253204 580796 253256 580848
rect 258172 580796 258224 580848
rect 286140 580796 286192 580848
rect 122932 580728 122984 580780
rect 150716 580728 150768 580780
rect 160560 580728 160612 580780
rect 171784 580728 171836 580780
rect 215024 580728 215076 580780
rect 225604 580728 225656 580780
rect 268936 580728 268988 580780
rect 279424 580728 279476 580780
rect 285772 580728 285824 580780
rect 312636 580796 312688 580848
rect 295984 580728 296036 580780
rect 307024 580728 307076 580780
rect 311992 580728 312044 580780
rect 340144 580796 340196 580848
rect 322848 580728 322900 580780
rect 333244 580728 333296 580780
rect 339592 580728 339644 580780
rect 366732 580796 366784 580848
rect 350080 580728 350132 580780
rect 359556 580728 359608 580780
rect 365812 580728 365864 580780
rect 393596 580796 393648 580848
rect 376576 580728 376628 580780
rect 387064 580728 387116 580780
rect 393412 580728 393464 580780
rect 420920 580796 420972 580848
rect 431040 580796 431092 580848
rect 442264 580796 442316 580848
rect 447232 580796 447284 580848
rect 474740 580796 474792 580848
rect 484952 580796 485004 580848
rect 496084 580796 496136 580848
rect 501052 580796 501104 580848
rect 528744 580796 528796 580848
rect 403992 580728 404044 580780
rect 414664 580728 414716 580780
rect 458088 580728 458140 580780
rect 468484 580728 468536 580780
rect 511908 580728 511960 580780
rect 522396 580728 522448 580780
rect 36544 580660 36596 580712
rect 538404 580660 538456 580712
rect 16304 578892 16356 578944
rect 528652 578892 528704 578944
rect 26056 578484 26108 578536
rect 149704 578484 149756 578536
rect 36728 578416 36780 578468
rect 52460 578416 52512 578468
rect 232320 578416 232372 578468
rect 251824 578416 251876 578468
rect 475384 578416 475436 578468
rect 494704 578416 494756 578468
rect 62488 578348 62540 578400
rect 79324 578348 79376 578400
rect 90456 578348 90508 578400
rect 106464 578348 106516 578400
rect 116492 578348 116544 578400
rect 133420 578348 133472 578400
rect 144184 578348 144236 578400
rect 160284 578348 160336 578400
rect 170496 578348 170548 578400
rect 187792 578348 187844 578400
rect 197544 578348 197596 578400
rect 214380 578348 214432 578400
rect 224500 578348 224552 578400
rect 241612 578348 241664 578400
rect 413468 578348 413520 578400
rect 430580 578348 430632 578400
rect 440516 578348 440568 578400
rect 457260 578348 457312 578400
rect 468484 578348 468536 578400
rect 484400 578348 484452 578400
rect 36820 578280 36872 578332
rect 62120 578280 62172 578332
rect 64144 578280 64196 578332
rect 89076 578280 89128 578332
rect 90364 578280 90416 578332
rect 116124 578280 116176 578332
rect 116584 578280 116636 578332
rect 142988 578280 143040 578332
rect 144276 578280 144328 578332
rect 170036 578280 170088 578332
rect 178408 578280 178460 578332
rect 200764 578280 200816 578332
rect 251456 578280 251508 578332
rect 268292 578280 268344 578332
rect 279424 578280 279476 578332
rect 295800 578280 295852 578332
rect 305552 578280 305604 578332
rect 322388 578280 322440 578332
rect 336004 578280 336056 578332
rect 349804 578280 349856 578332
rect 359648 578280 359700 578332
rect 376300 578280 376352 578332
rect 386512 578280 386564 578332
rect 403348 578280 403400 578332
rect 421288 578280 421340 578332
rect 446404 578280 446456 578332
rect 494520 578280 494572 578332
rect 511356 578280 511408 578332
rect 522396 578280 522448 578332
rect 538404 578280 538456 578332
rect 43352 578212 43404 578264
rect 62764 578212 62816 578264
rect 171784 578212 171836 578264
rect 197452 578212 197504 578264
rect 199384 578212 199436 578264
rect 223948 578212 224000 578264
rect 225604 578212 225656 578264
rect 251272 578212 251324 578264
rect 253204 578212 253256 578264
rect 278044 578212 278096 578264
rect 279516 578212 279568 578264
rect 305460 578212 305512 578264
rect 307024 578212 307076 578264
rect 331956 578212 332008 578264
rect 333244 578212 333296 578264
rect 359464 578212 359516 578264
rect 359740 578212 359792 578264
rect 386052 578212 386104 578264
rect 387064 578212 387116 578264
rect 412916 578212 412968 578264
rect 414664 578212 414716 578264
rect 440240 578212 440292 578264
rect 442264 578212 442316 578264
rect 467012 578212 467064 578264
rect 468576 578212 468628 578264
rect 494060 578212 494112 578264
rect 496084 578212 496136 578264
rect 520924 578212 520976 578264
rect 522304 578212 522356 578264
rect 547972 578212 548024 578264
rect 37924 576104 37976 576156
rect 526444 576104 526496 576156
rect 285772 575356 285824 575408
rect 286140 575356 286192 575408
rect 339592 575288 339644 575340
rect 340144 575288 340196 575340
rect 89720 562300 89772 562352
rect 90456 562300 90508 562352
rect 13728 557472 13780 557524
rect 64880 557472 64932 557524
rect 95148 557472 95200 557524
rect 146300 557472 146352 557524
rect 148968 557472 149020 557524
rect 200120 557472 200172 557524
rect 202788 557472 202840 557524
rect 253940 557472 253992 557524
rect 256608 557472 256660 557524
rect 307760 557472 307812 557524
rect 338028 557472 338080 557524
rect 389180 557472 389232 557524
rect 391848 557472 391900 557524
rect 443000 557472 443052 557524
rect 445668 557472 445720 557524
rect 496820 557472 496872 557524
rect 500868 557472 500920 557524
rect 550640 557472 550692 557524
rect 35624 557404 35676 557456
rect 36728 557404 36780 557456
rect 41328 557404 41380 557456
rect 91100 557404 91152 557456
rect 122748 557404 122800 557456
rect 172520 557404 172572 557456
rect 176568 557404 176620 557456
rect 226340 557404 226392 557456
rect 230388 557404 230440 557456
rect 280160 557404 280212 557456
rect 284208 557404 284260 557456
rect 335360 557404 335412 557456
rect 365628 557404 365680 557456
rect 415400 557404 415452 557456
rect 419448 557404 419500 557456
rect 68928 557336 68980 557388
rect 118700 557336 118752 557388
rect 311808 557336 311860 557388
rect 361580 557336 361632 557388
rect 469220 557404 469272 557456
rect 473268 557404 473320 557456
rect 523040 557404 523092 557456
rect 446404 556724 446456 556776
rect 447692 556724 447744 556776
rect 521752 556724 521804 556776
rect 522396 556724 522448 556776
rect 52736 554684 52788 554736
rect 64144 554684 64196 554736
rect 69112 554684 69164 554736
rect 15200 554616 15252 554668
rect 42984 554616 43036 554668
rect 62764 554616 62816 554668
rect 70032 554616 70084 554668
rect 96712 554684 96764 554736
rect 96988 554616 97040 554668
rect 146944 554684 146996 554736
rect 124036 554616 124088 554668
rect 133696 554616 133748 554668
rect 144276 554616 144328 554668
rect 150532 554616 150584 554668
rect 200764 554684 200816 554736
rect 204996 554684 205048 554736
rect 251824 554684 251876 554736
rect 259000 554684 259052 554736
rect 332324 554684 332376 554736
rect 336004 554684 336056 554736
rect 494704 554684 494756 554736
rect 501972 554684 502024 554736
rect 25688 554548 25740 554600
rect 36820 554548 36872 554600
rect 79692 554548 79744 554600
rect 90364 554548 90416 554600
rect 106648 554548 106700 554600
rect 116584 554548 116636 554600
rect 122932 554548 122984 554600
rect 150992 554548 151044 554600
rect 548340 554616 548392 554668
rect 178040 554548 178092 554600
rect 187700 554548 187752 554600
rect 199384 554548 199436 554600
rect 204352 554548 204404 554600
rect 232044 554548 232096 554600
rect 241704 554548 241756 554600
rect 253204 554548 253256 554600
rect 258172 554548 258224 554600
rect 286048 554548 286100 554600
rect 160652 554480 160704 554532
rect 171784 554480 171836 554532
rect 214656 554480 214708 554532
rect 225604 554480 225656 554532
rect 268660 554480 268712 554532
rect 279516 554480 279568 554532
rect 285772 554480 285824 554532
rect 313004 554548 313056 554600
rect 295708 554480 295760 554532
rect 307024 554480 307076 554532
rect 311992 554480 312044 554532
rect 340052 554548 340104 554600
rect 322664 554480 322716 554532
rect 333244 554480 333296 554532
rect 339592 554480 339644 554532
rect 367008 554548 367060 554600
rect 349712 554480 349764 554532
rect 359556 554480 359608 554532
rect 365812 554480 365864 554532
rect 393964 554548 394016 554600
rect 376668 554480 376720 554532
rect 387064 554480 387116 554532
rect 393412 554480 393464 554532
rect 421012 554548 421064 554600
rect 430672 554548 430724 554600
rect 442264 554548 442316 554600
rect 447232 554548 447284 554600
rect 475016 554548 475068 554600
rect 484676 554548 484728 554600
rect 496084 554548 496136 554600
rect 501052 554548 501104 554600
rect 529020 554548 529072 554600
rect 403716 554480 403768 554532
rect 414664 554480 414716 554532
rect 457720 554480 457772 554532
rect 468576 554480 468628 554532
rect 511724 554480 511776 554532
rect 522304 554480 522356 554532
rect 36636 554412 36688 554464
rect 538680 554412 538732 554464
rect 16028 551284 16080 551336
rect 529020 551284 529072 551336
rect 25688 550876 25740 550928
rect 146944 550876 146996 550928
rect 36636 550808 36688 550860
rect 52644 550808 52696 550860
rect 232044 550808 232096 550860
rect 251824 550808 251876 550860
rect 475016 550808 475068 550860
rect 494704 550808 494756 550860
rect 62488 550740 62540 550792
rect 79692 550740 79744 550792
rect 90456 550740 90508 550792
rect 106648 550740 106700 550792
rect 116492 550740 116544 550792
rect 133696 550740 133748 550792
rect 170496 550740 170548 550792
rect 187700 550740 187752 550792
rect 197452 550740 197504 550792
rect 214656 550740 214708 550792
rect 224500 550740 224552 550792
rect 241704 550740 241756 550792
rect 413468 550740 413520 550792
rect 430672 550740 430724 550792
rect 440516 550740 440568 550792
rect 457628 550740 457680 550792
rect 468484 550740 468536 550792
rect 484676 550740 484728 550792
rect 36820 550672 36872 550724
rect 62304 550672 62356 550724
rect 64144 550672 64196 550724
rect 89352 550672 89404 550724
rect 90364 550672 90416 550724
rect 116308 550672 116360 550724
rect 116584 550672 116636 550724
rect 143356 550672 143408 550724
rect 144276 550672 144328 550724
rect 170312 550672 170364 550724
rect 178040 550672 178092 550724
rect 200764 550672 200816 550724
rect 251456 550672 251508 550724
rect 268660 550672 268712 550724
rect 279516 550672 279568 550724
rect 295708 550672 295760 550724
rect 305460 550672 305512 550724
rect 322664 550672 322716 550724
rect 334624 550672 334676 550724
rect 349712 550672 349764 550724
rect 359464 550672 359516 550724
rect 376668 550672 376720 550724
rect 386512 550672 386564 550724
rect 403624 550672 403676 550724
rect 421012 550672 421064 550724
rect 443644 550672 443696 550724
rect 494520 550672 494572 550724
rect 511632 550672 511684 550724
rect 522304 550672 522356 550724
rect 538680 550672 538732 550724
rect 43076 550604 43128 550656
rect 62764 550604 62816 550656
rect 144184 550604 144236 550656
rect 160652 550604 160704 550656
rect 171784 550604 171836 550656
rect 197360 550604 197412 550656
rect 199384 550604 199436 550656
rect 224316 550604 224368 550656
rect 225604 550604 225656 550656
rect 251364 550604 251416 550656
rect 253204 550604 253256 550656
rect 278320 550604 278372 550656
rect 279424 550604 279476 550656
rect 305368 550604 305420 550656
rect 307024 550604 307076 550656
rect 332324 550604 332376 550656
rect 333244 550604 333296 550656
rect 359372 550604 359424 550656
rect 359556 550604 359608 550656
rect 386328 550604 386380 550656
rect 387064 550604 387116 550656
rect 413284 550604 413336 550656
rect 414664 550604 414716 550656
rect 440332 550604 440384 550656
rect 442264 550604 442316 550656
rect 467288 550604 467340 550656
rect 468576 550604 468628 550656
rect 494336 550604 494388 550656
rect 496084 550604 496136 550656
rect 521292 550604 521344 550656
rect 522396 550604 522448 550656
rect 548340 550604 548392 550656
rect 37924 548496 37976 548548
rect 526444 548496 526496 548548
rect 35624 547884 35676 547936
rect 36728 547884 36780 547936
rect 89720 533604 89772 533656
rect 90456 533604 90508 533656
rect 13728 529864 13780 529916
rect 64880 529864 64932 529916
rect 95148 529864 95200 529916
rect 146300 529864 146352 529916
rect 148968 529864 149020 529916
rect 200120 529864 200172 529916
rect 202788 529864 202840 529916
rect 253940 529864 253992 529916
rect 256608 529864 256660 529916
rect 307760 529864 307812 529916
rect 332508 529864 332560 529916
rect 334624 529864 334676 529916
rect 338028 529864 338080 529916
rect 389180 529864 389232 529916
rect 391848 529864 391900 529916
rect 443000 529864 443052 529916
rect 445668 529864 445720 529916
rect 496820 529864 496872 529916
rect 500868 529864 500920 529916
rect 550640 529864 550692 529916
rect 35624 529796 35676 529848
rect 36636 529796 36688 529848
rect 41328 529796 41380 529848
rect 91100 529796 91152 529848
rect 122748 529796 122800 529848
rect 172520 529796 172572 529848
rect 176568 529796 176620 529848
rect 226340 529796 226392 529848
rect 230388 529796 230440 529848
rect 68928 529728 68980 529780
rect 118700 529728 118752 529780
rect 278688 529796 278740 529848
rect 279516 529796 279568 529848
rect 284208 529796 284260 529848
rect 335360 529796 335412 529848
rect 365628 529796 365680 529848
rect 415400 529796 415452 529848
rect 419448 529796 419500 529848
rect 469220 529796 469272 529848
rect 473268 529796 473320 529848
rect 523040 529796 523092 529848
rect 280160 529728 280212 529780
rect 311808 529728 311860 529780
rect 361580 529728 361632 529780
rect 116216 529592 116268 529644
rect 116492 529592 116544 529644
rect 170220 529592 170272 529644
rect 170496 529592 170548 529644
rect 53104 527076 53156 527128
rect 64144 527076 64196 527128
rect 69112 527076 69164 527128
rect 15200 527008 15252 527060
rect 42800 527008 42852 527060
rect 62764 527008 62816 527060
rect 69756 527008 69808 527060
rect 96712 527076 96764 527128
rect 96804 527008 96856 527060
rect 200764 527076 200816 527128
rect 204628 527076 204680 527128
rect 251824 527076 251876 527128
rect 258724 527076 258776 527128
rect 443644 527076 443696 527128
rect 447692 527076 447744 527128
rect 494704 527076 494756 527128
rect 501604 527076 501656 527128
rect 123668 527008 123720 527060
rect 149704 527008 149756 527060
rect 547972 527008 548024 527060
rect 26056 526940 26108 526992
rect 36820 526940 36872 526992
rect 79968 526940 80020 526992
rect 90364 526940 90416 526992
rect 106556 526940 106608 526992
rect 116584 526940 116636 526992
rect 133788 526940 133840 526992
rect 144276 526940 144328 526992
rect 150532 526940 150584 526992
rect 178132 526940 178184 526992
rect 187976 526940 188028 526992
rect 199384 526940 199436 526992
rect 204352 526940 204404 526992
rect 231952 526940 232004 526992
rect 242072 526940 242124 526992
rect 253204 526940 253256 526992
rect 258172 526940 258224 526992
rect 122932 526872 122984 526924
rect 150716 526872 150768 526924
rect 160560 526872 160612 526924
rect 171784 526872 171836 526924
rect 215024 526872 215076 526924
rect 225604 526872 225656 526924
rect 268936 526872 268988 526924
rect 279424 526872 279476 526924
rect 285772 526940 285824 526992
rect 312636 526940 312688 526992
rect 286140 526872 286192 526924
rect 295984 526872 296036 526924
rect 307024 526872 307076 526924
rect 311992 526872 312044 526924
rect 340144 526940 340196 526992
rect 322848 526872 322900 526924
rect 333244 526872 333296 526924
rect 339592 526872 339644 526924
rect 366732 526940 366784 526992
rect 350080 526872 350132 526924
rect 359556 526872 359608 526924
rect 365812 526872 365864 526924
rect 393596 526940 393648 526992
rect 376576 526872 376628 526924
rect 387064 526872 387116 526924
rect 393412 526872 393464 526924
rect 420920 526940 420972 526992
rect 431040 526940 431092 526992
rect 442264 526940 442316 526992
rect 447232 526940 447284 526992
rect 474740 526940 474792 526992
rect 484952 526940 485004 526992
rect 496084 526940 496136 526992
rect 501052 526940 501104 526992
rect 528652 526940 528704 526992
rect 403992 526872 404044 526924
rect 414664 526872 414716 526924
rect 458088 526872 458140 526924
rect 468576 526872 468628 526924
rect 511816 526872 511868 526924
rect 522396 526872 522448 526924
rect 36544 526804 36596 526856
rect 538404 526804 538456 526856
rect 527088 525716 527140 525768
rect 579804 525716 579856 525768
rect 16304 523676 16356 523728
rect 528744 523676 528796 523728
rect 25964 523268 26016 523320
rect 149704 523268 149756 523320
rect 36820 523200 36872 523252
rect 52460 523200 52512 523252
rect 232320 523200 232372 523252
rect 251824 523200 251876 523252
rect 475384 523200 475436 523252
rect 494704 523200 494756 523252
rect 62488 523132 62540 523184
rect 79324 523132 79376 523184
rect 90456 523132 90508 523184
rect 106372 523132 106424 523184
rect 116492 523132 116544 523184
rect 133420 523132 133472 523184
rect 144184 523132 144236 523184
rect 160284 523132 160336 523184
rect 170496 523132 170548 523184
rect 187792 523132 187844 523184
rect 197544 523132 197596 523184
rect 214380 523132 214432 523184
rect 224500 523132 224552 523184
rect 241520 523132 241572 523184
rect 413468 523132 413520 523184
rect 430580 523132 430632 523184
rect 440516 523132 440568 523184
rect 457260 523132 457312 523184
rect 468484 523132 468536 523184
rect 484400 523132 484452 523184
rect 36544 523064 36596 523116
rect 62120 523064 62172 523116
rect 64144 523064 64196 523116
rect 89076 523064 89128 523116
rect 90364 523064 90416 523116
rect 115940 523064 115992 523116
rect 116584 523064 116636 523116
rect 142988 523064 143040 523116
rect 144276 523064 144328 523116
rect 170036 523064 170088 523116
rect 178408 523064 178460 523116
rect 200764 523064 200816 523116
rect 251456 523064 251508 523116
rect 268292 523064 268344 523116
rect 279516 523064 279568 523116
rect 295800 523064 295852 523116
rect 305552 523064 305604 523116
rect 322388 523064 322440 523116
rect 334624 523064 334676 523116
rect 349804 523064 349856 523116
rect 359556 523064 359608 523116
rect 376300 523064 376352 523116
rect 386512 523064 386564 523116
rect 403348 523064 403400 523116
rect 421288 523064 421340 523116
rect 443644 523064 443696 523116
rect 494520 523064 494572 523116
rect 511356 523064 511408 523116
rect 522396 523064 522448 523116
rect 538404 523064 538456 523116
rect 43352 522996 43404 523048
rect 62764 522996 62816 523048
rect 171784 522996 171836 523048
rect 197452 522996 197504 523048
rect 199384 522996 199436 523048
rect 223948 522996 224000 523048
rect 225604 522996 225656 523048
rect 251180 522996 251232 523048
rect 253204 522996 253256 523048
rect 278044 522996 278096 523048
rect 279424 522996 279476 523048
rect 305460 522996 305512 523048
rect 307024 522996 307076 523048
rect 331956 522996 332008 523048
rect 333244 522996 333296 523048
rect 359464 522996 359516 523048
rect 359740 522996 359792 523048
rect 386052 522996 386104 523048
rect 387064 522996 387116 523048
rect 412916 522996 412968 523048
rect 414664 522996 414716 523048
rect 440240 522996 440292 523048
rect 442264 522996 442316 523048
rect 467012 522996 467064 523048
rect 468576 522996 468628 523048
rect 494060 522996 494112 523048
rect 496084 522996 496136 523048
rect 520924 522996 520976 523048
rect 522304 522996 522356 523048
rect 548064 522996 548116 523048
rect 37924 522248 37976 522300
rect 526444 522248 526496 522300
rect 35624 521704 35676 521756
rect 36636 521704 36688 521756
rect 285772 521364 285824 521416
rect 286140 521364 286192 521416
rect 339592 521296 339644 521348
rect 340144 521296 340196 521348
rect 68928 520412 68980 520464
rect 118700 520412 118752 520464
rect 311808 520412 311860 520464
rect 361580 520412 361632 520464
rect 41328 520344 41380 520396
rect 91100 520344 91152 520396
rect 122748 520344 122800 520396
rect 172520 520344 172572 520396
rect 176568 520344 176620 520396
rect 226340 520344 226392 520396
rect 231860 520344 231912 520396
rect 280160 520344 280212 520396
rect 284208 520344 284260 520396
rect 335360 520344 335412 520396
rect 365628 520344 365680 520396
rect 415400 520344 415452 520396
rect 419448 520344 419500 520396
rect 469220 520344 469272 520396
rect 474832 520344 474884 520396
rect 523040 520344 523092 520396
rect 13728 520276 13780 520328
rect 64880 520276 64932 520328
rect 96896 520276 96948 520328
rect 146300 520276 146352 520328
rect 148968 520276 149020 520328
rect 200120 520276 200172 520328
rect 204904 520276 204956 520328
rect 253940 520276 253992 520328
rect 256608 520276 256660 520328
rect 307760 520276 307812 520328
rect 339868 520276 339920 520328
rect 389180 520276 389232 520328
rect 391848 520276 391900 520328
rect 443000 520276 443052 520328
rect 445668 520276 445720 520328
rect 496820 520276 496872 520328
rect 500868 520276 500920 520328
rect 550640 520276 550692 520328
rect 230388 518848 230440 518900
rect 231860 518848 231912 518900
rect 473268 518848 473320 518900
rect 474832 518848 474884 518900
rect 89720 505588 89772 505640
rect 90456 505588 90508 505640
rect 521752 505588 521804 505640
rect 522396 505588 522448 505640
rect 278688 503616 278740 503668
rect 279516 503616 279568 503668
rect 332508 503616 332560 503668
rect 334624 503616 334676 503668
rect 35624 502256 35676 502308
rect 36820 502256 36872 502308
rect 52736 500896 52788 500948
rect 64144 500896 64196 500948
rect 69112 500896 69164 500948
rect 15200 500828 15252 500880
rect 42984 500828 43036 500880
rect 62764 500828 62816 500880
rect 70032 500828 70084 500880
rect 96712 500896 96764 500948
rect 96988 500828 97040 500880
rect 146944 500896 146996 500948
rect 124036 500828 124088 500880
rect 133696 500828 133748 500880
rect 144276 500828 144328 500880
rect 25688 500760 25740 500812
rect 36544 500760 36596 500812
rect 79692 500760 79744 500812
rect 90364 500760 90416 500812
rect 106648 500760 106700 500812
rect 116584 500760 116636 500812
rect 122932 500760 122984 500812
rect 150992 500828 151044 500880
rect 200764 500896 200816 500948
rect 204996 500896 205048 500948
rect 251824 500896 251876 500948
rect 259000 500896 259052 500948
rect 443644 500896 443696 500948
rect 447968 500896 448020 500948
rect 494704 500896 494756 500948
rect 501972 500896 502024 500948
rect 548340 500828 548392 500880
rect 150532 500760 150584 500812
rect 178040 500760 178092 500812
rect 187700 500760 187752 500812
rect 199384 500760 199436 500812
rect 204352 500760 204404 500812
rect 232044 500760 232096 500812
rect 241704 500760 241756 500812
rect 253204 500760 253256 500812
rect 258172 500760 258224 500812
rect 160652 500692 160704 500744
rect 171784 500692 171836 500744
rect 214656 500692 214708 500744
rect 225604 500692 225656 500744
rect 268660 500692 268712 500744
rect 279424 500692 279476 500744
rect 285772 500760 285824 500812
rect 313004 500760 313056 500812
rect 286048 500692 286100 500744
rect 295708 500692 295760 500744
rect 307024 500692 307076 500744
rect 311992 500692 312044 500744
rect 340052 500760 340104 500812
rect 322664 500692 322716 500744
rect 333244 500692 333296 500744
rect 339592 500692 339644 500744
rect 367008 500760 367060 500812
rect 349712 500692 349764 500744
rect 359556 500692 359608 500744
rect 365812 500692 365864 500744
rect 393964 500760 394016 500812
rect 376668 500692 376720 500744
rect 387064 500692 387116 500744
rect 393412 500692 393464 500744
rect 421012 500760 421064 500812
rect 430672 500760 430724 500812
rect 442264 500760 442316 500812
rect 447232 500760 447284 500812
rect 475016 500760 475068 500812
rect 484676 500760 484728 500812
rect 496084 500760 496136 500812
rect 501052 500760 501104 500812
rect 529020 500760 529072 500812
rect 403716 500692 403768 500744
rect 414664 500692 414716 500744
rect 457720 500692 457772 500744
rect 468576 500692 468628 500744
rect 511724 500692 511776 500744
rect 522304 500692 522356 500744
rect 36728 500624 36780 500676
rect 538680 500624 538732 500676
rect 16028 497428 16080 497480
rect 529020 497428 529072 497480
rect 25688 497088 25740 497140
rect 146944 497088 146996 497140
rect 36728 497020 36780 497072
rect 52644 497020 52696 497072
rect 232044 497020 232096 497072
rect 251824 497020 251876 497072
rect 475016 497020 475068 497072
rect 494704 497020 494756 497072
rect 62488 496952 62540 497004
rect 79692 496952 79744 497004
rect 90364 496952 90416 497004
rect 106648 496952 106700 497004
rect 116492 496952 116544 497004
rect 133696 496952 133748 497004
rect 170496 496952 170548 497004
rect 187700 496952 187752 497004
rect 197452 496952 197504 497004
rect 214656 496952 214708 497004
rect 224500 496952 224552 497004
rect 241704 496952 241756 497004
rect 413468 496952 413520 497004
rect 430672 496952 430724 497004
rect 440516 496952 440568 497004
rect 457628 496952 457680 497004
rect 468576 496952 468628 497004
rect 484676 496952 484728 497004
rect 36820 496884 36872 496936
rect 62304 496884 62356 496936
rect 64144 496884 64196 496936
rect 89352 496884 89404 496936
rect 90456 496884 90508 496936
rect 116308 496884 116360 496936
rect 116584 496884 116636 496936
rect 143356 496884 143408 496936
rect 144276 496884 144328 496936
rect 170312 496884 170364 496936
rect 178040 496884 178092 496936
rect 200764 496884 200816 496936
rect 251456 496884 251508 496936
rect 268660 496884 268712 496936
rect 279516 496884 279568 496936
rect 295708 496884 295760 496936
rect 305460 496884 305512 496936
rect 322664 496884 322716 496936
rect 334624 496884 334676 496936
rect 349712 496884 349764 496936
rect 359464 496884 359516 496936
rect 376668 496884 376720 496936
rect 386512 496884 386564 496936
rect 403624 496884 403676 496936
rect 421012 496884 421064 496936
rect 443644 496884 443696 496936
rect 494520 496884 494572 496936
rect 511632 496884 511684 496936
rect 522396 496884 522448 496936
rect 538680 496884 538732 496936
rect 43076 496816 43128 496868
rect 62764 496816 62816 496868
rect 144184 496816 144236 496868
rect 160652 496816 160704 496868
rect 171784 496816 171836 496868
rect 197360 496816 197412 496868
rect 199384 496816 199436 496868
rect 224316 496816 224368 496868
rect 225604 496816 225656 496868
rect 251364 496816 251416 496868
rect 253204 496816 253256 496868
rect 278320 496816 278372 496868
rect 279424 496816 279476 496868
rect 305368 496816 305420 496868
rect 307024 496816 307076 496868
rect 332324 496816 332376 496868
rect 333244 496816 333296 496868
rect 359372 496816 359424 496868
rect 359556 496816 359608 496868
rect 386328 496816 386380 496868
rect 387064 496816 387116 496868
rect 413284 496816 413336 496868
rect 414664 496816 414716 496868
rect 440332 496816 440384 496868
rect 442264 496816 442316 496868
rect 467288 496816 467340 496868
rect 468484 496816 468536 496868
rect 494336 496816 494388 496868
rect 496084 496816 496136 496868
rect 521292 496816 521344 496868
rect 522304 496816 522356 496868
rect 548340 496816 548392 496868
rect 37924 494708 37976 494760
rect 526444 494708 526496 494760
rect 68928 494096 68980 494148
rect 118700 494096 118752 494148
rect 122748 494096 122800 494148
rect 172520 494096 172572 494148
rect 230388 494096 230440 494148
rect 280160 494096 280212 494148
rect 311808 494096 311860 494148
rect 361580 494096 361632 494148
rect 500868 494096 500920 494148
rect 550640 494096 550692 494148
rect 41328 494028 41380 494080
rect 91100 494028 91152 494080
rect 148968 494028 149020 494080
rect 200120 494028 200172 494080
rect 202788 494028 202840 494080
rect 253940 494028 253992 494080
rect 284208 494028 284260 494080
rect 335360 494028 335412 494080
rect 365628 494028 365680 494080
rect 415400 494028 415452 494080
rect 419448 494028 419500 494080
rect 469220 494028 469272 494080
rect 473268 494028 473320 494080
rect 523040 494028 523092 494080
rect 521752 477640 521804 477692
rect 522396 477640 522448 477692
rect 13728 476008 13780 476060
rect 64880 476008 64932 476060
rect 95148 476008 95200 476060
rect 146300 476008 146352 476060
rect 176568 476008 176620 476060
rect 226340 476008 226392 476060
rect 256608 476008 256660 476060
rect 307760 476008 307812 476060
rect 332508 476008 332560 476060
rect 334624 476008 334676 476060
rect 338028 476008 338080 476060
rect 389180 476008 389232 476060
rect 391848 476008 391900 476060
rect 443000 476008 443052 476060
rect 445668 476008 445720 476060
rect 496820 476008 496872 476060
rect 35624 475940 35676 475992
rect 36728 475940 36780 475992
rect 278688 475940 278740 475992
rect 279516 475940 279568 475992
rect 467656 475940 467708 475992
rect 468576 475940 468628 475992
rect 116216 475600 116268 475652
rect 116492 475600 116544 475652
rect 170220 475600 170272 475652
rect 170496 475600 170548 475652
rect 62764 473288 62816 473340
rect 69756 473288 69808 473340
rect 96712 473288 96764 473340
rect 15200 473220 15252 473272
rect 42800 473220 42852 473272
rect 53104 473220 53156 473272
rect 64144 473220 64196 473272
rect 69112 473220 69164 473272
rect 96804 473220 96856 473272
rect 200764 473288 200816 473340
rect 204628 473288 204680 473340
rect 251824 473288 251876 473340
rect 258724 473288 258776 473340
rect 443644 473288 443696 473340
rect 447692 473288 447744 473340
rect 494704 473288 494756 473340
rect 501604 473288 501656 473340
rect 123668 473220 123720 473272
rect 149704 473220 149756 473272
rect 547972 473220 548024 473272
rect 26056 473152 26108 473204
rect 36820 473152 36872 473204
rect 79968 473152 80020 473204
rect 90456 473152 90508 473204
rect 106556 473152 106608 473204
rect 116584 473152 116636 473204
rect 133788 473152 133840 473204
rect 144276 473152 144328 473204
rect 150532 473152 150584 473204
rect 178132 473152 178184 473204
rect 187976 473152 188028 473204
rect 199384 473152 199436 473204
rect 204352 473152 204404 473204
rect 231860 473152 231912 473204
rect 242072 473152 242124 473204
rect 253204 473152 253256 473204
rect 258172 473152 258224 473204
rect 286140 473152 286192 473204
rect 122932 473084 122984 473136
rect 150716 473084 150768 473136
rect 160560 473084 160612 473136
rect 171784 473084 171836 473136
rect 215024 473084 215076 473136
rect 225604 473084 225656 473136
rect 268936 473084 268988 473136
rect 279424 473084 279476 473136
rect 285772 473084 285824 473136
rect 312636 473152 312688 473204
rect 295984 473084 296036 473136
rect 307024 473084 307076 473136
rect 311992 473084 312044 473136
rect 340144 473152 340196 473204
rect 322848 473084 322900 473136
rect 333244 473084 333296 473136
rect 339592 473084 339644 473136
rect 366732 473152 366784 473204
rect 350080 473084 350132 473136
rect 359556 473084 359608 473136
rect 365812 473084 365864 473136
rect 393596 473152 393648 473204
rect 376576 473084 376628 473136
rect 387064 473084 387116 473136
rect 393412 473084 393464 473136
rect 420920 473152 420972 473204
rect 431040 473152 431092 473204
rect 442264 473152 442316 473204
rect 447232 473152 447284 473204
rect 474740 473152 474792 473204
rect 484952 473152 485004 473204
rect 496084 473152 496136 473204
rect 501052 473152 501104 473204
rect 528652 473152 528704 473204
rect 403992 473084 404044 473136
rect 414664 473084 414716 473136
rect 458088 473084 458140 473136
rect 468484 473084 468536 473136
rect 511908 473084 511960 473136
rect 522304 473084 522356 473136
rect 36636 473016 36688 473068
rect 538404 473016 538456 473068
rect 15292 469820 15344 469872
rect 528744 469820 528796 469872
rect 25964 469480 26016 469532
rect 149704 469480 149756 469532
rect 35716 469412 35768 469464
rect 52460 469412 52512 469464
rect 232320 469412 232372 469464
rect 251824 469412 251876 469464
rect 62488 469344 62540 469396
rect 79324 469344 79376 469396
rect 90456 469344 90508 469396
rect 106372 469344 106424 469396
rect 116492 469344 116544 469396
rect 133420 469344 133472 469396
rect 144276 469344 144328 469396
rect 160284 469344 160336 469396
rect 170496 469344 170548 469396
rect 187792 469344 187844 469396
rect 197544 469344 197596 469396
rect 214380 469344 214432 469396
rect 224500 469344 224552 469396
rect 241520 469344 241572 469396
rect 413468 469344 413520 469396
rect 430580 469344 430632 469396
rect 440516 469344 440568 469396
rect 457260 469344 457312 469396
rect 36728 469276 36780 469328
rect 62120 469276 62172 469328
rect 64144 469276 64196 469328
rect 89076 469276 89128 469328
rect 90364 469276 90416 469328
rect 115940 469276 115992 469328
rect 116584 469276 116636 469328
rect 142988 469276 143040 469328
rect 144184 469276 144236 469328
rect 170036 469276 170088 469328
rect 178408 469276 178460 469328
rect 200764 469276 200816 469328
rect 251456 469276 251508 469328
rect 268292 469276 268344 469328
rect 279516 469276 279568 469328
rect 295800 469276 295852 469328
rect 305552 469276 305604 469328
rect 322388 469276 322440 469328
rect 336004 469276 336056 469328
rect 349804 469276 349856 469328
rect 359556 469276 359608 469328
rect 376300 469276 376352 469328
rect 386512 469276 386564 469328
rect 403348 469276 403400 469328
rect 421288 469276 421340 469328
rect 446404 469276 446456 469328
rect 467472 469276 467524 469328
rect 484400 469276 484452 469328
rect 494520 469276 494572 469328
rect 511356 469276 511408 469328
rect 522304 469276 522356 469328
rect 538404 469276 538456 469328
rect 43352 469208 43404 469260
rect 62764 469208 62816 469260
rect 171784 469208 171836 469260
rect 197452 469208 197504 469260
rect 199384 469208 199436 469260
rect 223948 469208 224000 469260
rect 225604 469208 225656 469260
rect 251180 469208 251232 469260
rect 253204 469208 253256 469260
rect 278044 469208 278096 469260
rect 279424 469208 279476 469260
rect 305460 469208 305512 469260
rect 307024 469208 307076 469260
rect 331956 469208 332008 469260
rect 333244 469208 333296 469260
rect 359464 469208 359516 469260
rect 359740 469208 359792 469260
rect 386052 469208 386104 469260
rect 387064 469208 387116 469260
rect 412916 469208 412968 469260
rect 414664 469208 414716 469260
rect 440240 469208 440292 469260
rect 442264 469208 442316 469260
rect 467012 469208 467064 469260
rect 468484 469208 468536 469260
rect 494060 469208 494112 469260
rect 496084 469208 496136 469260
rect 520924 469208 520976 469260
rect 522396 469208 522448 469260
rect 548064 469208 548116 469260
rect 37924 468460 37976 468512
rect 526444 468460 526496 468512
rect 339592 467304 339644 467356
rect 340144 467304 340196 467356
rect 68928 466556 68980 466608
rect 118700 466556 118752 466608
rect 230388 466556 230440 466608
rect 280160 466556 280212 466608
rect 35624 466488 35676 466540
rect 36636 466488 36688 466540
rect 41328 466488 41380 466540
rect 91100 466488 91152 466540
rect 122748 466488 122800 466540
rect 172520 466488 172572 466540
rect 176568 466488 176620 466540
rect 226340 466488 226392 466540
rect 256608 466488 256660 466540
rect 307760 466488 307812 466540
rect 311808 466488 311860 466540
rect 361580 466488 361632 466540
rect 365628 466488 365680 466540
rect 415400 466488 415452 466540
rect 419448 466488 419500 466540
rect 469220 466488 469272 466540
rect 473268 466488 473320 466540
rect 523040 466488 523092 466540
rect 13728 466420 13780 466472
rect 64880 466420 64932 466472
rect 95148 466420 95200 466472
rect 146300 466420 146352 466472
rect 148968 466420 149020 466472
rect 200120 466420 200172 466472
rect 202788 466420 202840 466472
rect 253940 466420 253992 466472
rect 284208 466420 284260 466472
rect 335360 466420 335412 466472
rect 338028 466420 338080 466472
rect 389180 466420 389232 466472
rect 391848 466420 391900 466472
rect 443000 466420 443052 466472
rect 445668 466420 445720 466472
rect 496820 466420 496872 466472
rect 500868 466420 500920 466472
rect 550640 466420 550692 466472
rect 143632 449624 143684 449676
rect 144276 449624 144328 449676
rect 89720 448468 89772 448520
rect 90456 448468 90508 448520
rect 200764 448468 200816 448520
rect 204628 448468 204680 448520
rect 278688 448468 278740 448520
rect 279516 448468 279568 448520
rect 332600 448468 332652 448520
rect 336004 448468 336056 448520
rect 446404 448468 446456 448520
rect 447692 448468 447744 448520
rect 25688 445680 25740 445732
rect 36728 445680 36780 445732
rect 62764 445680 62816 445732
rect 70032 445680 70084 445732
rect 96712 445680 96764 445732
rect 15200 445612 15252 445664
rect 42984 445612 43036 445664
rect 52736 445612 52788 445664
rect 64144 445612 64196 445664
rect 69112 445612 69164 445664
rect 96988 445612 97040 445664
rect 146944 445680 146996 445732
rect 124036 445612 124088 445664
rect 133696 445612 133748 445664
rect 144184 445612 144236 445664
rect 79692 445544 79744 445596
rect 90364 445544 90416 445596
rect 106648 445544 106700 445596
rect 116584 445544 116636 445596
rect 122932 445544 122984 445596
rect 150992 445612 151044 445664
rect 251824 445680 251876 445732
rect 259000 445680 259052 445732
rect 548340 445612 548392 445664
rect 150532 445544 150584 445596
rect 178040 445544 178092 445596
rect 187700 445544 187752 445596
rect 199384 445544 199436 445596
rect 204352 445544 204404 445596
rect 232044 445544 232096 445596
rect 241704 445544 241756 445596
rect 253204 445544 253256 445596
rect 258172 445544 258224 445596
rect 160652 445476 160704 445528
rect 171784 445476 171836 445528
rect 214656 445476 214708 445528
rect 225604 445476 225656 445528
rect 268660 445476 268712 445528
rect 279424 445476 279476 445528
rect 285772 445544 285824 445596
rect 313004 445544 313056 445596
rect 286048 445476 286100 445528
rect 295708 445476 295760 445528
rect 307024 445476 307076 445528
rect 311992 445476 312044 445528
rect 340052 445544 340104 445596
rect 322664 445476 322716 445528
rect 333244 445476 333296 445528
rect 339592 445476 339644 445528
rect 349712 445476 349764 445528
rect 359556 445476 359608 445528
rect 365812 445544 365864 445596
rect 393964 445544 394016 445596
rect 367008 445476 367060 445528
rect 376668 445476 376720 445528
rect 387064 445476 387116 445528
rect 393412 445476 393464 445528
rect 421012 445544 421064 445596
rect 430672 445544 430724 445596
rect 442264 445544 442316 445596
rect 447232 445544 447284 445596
rect 475016 445544 475068 445596
rect 403716 445476 403768 445528
rect 414664 445476 414716 445528
rect 457720 445476 457772 445528
rect 468484 445476 468536 445528
rect 474832 445476 474884 445528
rect 484676 445476 484728 445528
rect 496084 445476 496136 445528
rect 501052 445544 501104 445596
rect 529020 445544 529072 445596
rect 501972 445476 502024 445528
rect 511724 445476 511776 445528
rect 522396 445476 522448 445528
rect 36544 445408 36596 445460
rect 538680 445408 538732 445460
rect 16028 443640 16080 443692
rect 529020 443640 529072 443692
rect 25688 443232 25740 443284
rect 146944 443232 146996 443284
rect 36728 443164 36780 443216
rect 52644 443164 52696 443216
rect 232044 443164 232096 443216
rect 251824 443164 251876 443216
rect 502064 443164 502116 443216
rect 522488 443164 522540 443216
rect 62488 443096 62540 443148
rect 79692 443096 79744 443148
rect 90456 443096 90508 443148
rect 106648 443096 106700 443148
rect 116492 443096 116544 443148
rect 133696 443096 133748 443148
rect 170496 443096 170548 443148
rect 187700 443096 187752 443148
rect 197452 443096 197504 443148
rect 214656 443096 214708 443148
rect 224500 443096 224552 443148
rect 241704 443096 241756 443148
rect 305460 443096 305512 443148
rect 322664 443096 322716 443148
rect 413468 443096 413520 443148
rect 430672 443096 430724 443148
rect 440516 443096 440568 443148
rect 457260 443096 457312 443148
rect 468576 443096 468628 443148
rect 484676 443096 484728 443148
rect 494520 443096 494572 443148
rect 511632 443096 511684 443148
rect 36820 443028 36872 443080
rect 62304 443028 62356 443080
rect 64144 443028 64196 443080
rect 89352 443028 89404 443080
rect 90364 443028 90416 443080
rect 116308 443028 116360 443080
rect 116584 443028 116636 443080
rect 143356 443028 143408 443080
rect 144276 443028 144328 443080
rect 170312 443028 170364 443080
rect 178040 443028 178092 443080
rect 200764 443028 200816 443080
rect 251456 443028 251508 443080
rect 268660 443028 268712 443080
rect 279516 443028 279568 443080
rect 295708 443028 295760 443080
rect 313004 443028 313056 443080
rect 333336 443028 333388 443080
rect 334624 443028 334676 443080
rect 349712 443028 349764 443080
rect 359464 443028 359516 443080
rect 376668 443028 376720 443080
rect 386512 443028 386564 443080
rect 403348 443028 403400 443080
rect 421012 443028 421064 443080
rect 443644 443028 443696 443080
rect 475016 443028 475068 443080
rect 494704 443028 494756 443080
rect 522304 443028 522356 443080
rect 538680 443028 538732 443080
rect 43352 442960 43404 443012
rect 62764 442960 62816 443012
rect 144184 442960 144236 443012
rect 160652 442960 160704 443012
rect 171784 442960 171836 443012
rect 197360 442960 197412 443012
rect 199384 442960 199436 443012
rect 224316 442960 224368 443012
rect 225604 442960 225656 443012
rect 251364 442960 251416 443012
rect 253204 442960 253256 443012
rect 278320 442960 278372 443012
rect 279424 442960 279476 443012
rect 305368 442960 305420 443012
rect 307024 442960 307076 443012
rect 332324 442960 332376 443012
rect 333244 442960 333296 443012
rect 359372 442960 359424 443012
rect 359556 442960 359608 443012
rect 386328 442960 386380 443012
rect 387064 442960 387116 443012
rect 412916 442960 412968 443012
rect 414664 442960 414716 443012
rect 440332 442960 440384 443012
rect 442264 442960 442316 443012
rect 467012 442960 467064 443012
rect 468484 442960 468536 443012
rect 494336 442960 494388 443012
rect 496084 442960 496136 443012
rect 521292 442960 521344 443012
rect 522396 442960 522448 443012
rect 548340 442960 548392 443012
rect 37924 440852 37976 440904
rect 526444 440852 526496 440904
rect 68928 440376 68980 440428
rect 118700 440376 118752 440428
rect 311808 440376 311860 440428
rect 361580 440376 361632 440428
rect 41328 440308 41380 440360
rect 91100 440308 91152 440360
rect 122748 440308 122800 440360
rect 172520 440308 172572 440360
rect 176568 440308 176620 440360
rect 226340 440308 226392 440360
rect 230388 440308 230440 440360
rect 280160 440308 280212 440360
rect 284208 440308 284260 440360
rect 335360 440308 335412 440360
rect 338028 440308 338080 440360
rect 13728 440240 13780 440292
rect 64880 440240 64932 440292
rect 95148 440240 95200 440292
rect 146300 440240 146352 440292
rect 148968 440240 149020 440292
rect 200120 440240 200172 440292
rect 202788 440240 202840 440292
rect 253940 440240 253992 440292
rect 256608 440240 256660 440292
rect 307760 440240 307812 440292
rect 339592 440240 339644 440292
rect 340144 440240 340196 440292
rect 365628 440308 365680 440360
rect 415400 440308 415452 440360
rect 419448 440308 419500 440360
rect 469220 440308 469272 440360
rect 473268 440308 473320 440360
rect 523040 440308 523092 440360
rect 389180 440240 389232 440292
rect 391848 440240 391900 440292
rect 443000 440240 443052 440292
rect 445668 440240 445720 440292
rect 496820 440240 496872 440292
rect 500868 440240 500920 440292
rect 550640 440240 550692 440292
rect 89720 423784 89772 423836
rect 90456 423784 90508 423836
rect 522488 423036 522540 423088
rect 528652 423036 528704 423088
rect 333336 422900 333388 422952
rect 339868 422900 339920 422952
rect 35624 422220 35676 422272
rect 36728 422220 36780 422272
rect 278688 421676 278740 421728
rect 279516 421676 279568 421728
rect 332508 421676 332560 421728
rect 334624 421676 334676 421728
rect 467656 421676 467708 421728
rect 468576 421676 468628 421728
rect 170220 421608 170272 421660
rect 170496 421608 170548 421660
rect 53104 419432 53156 419484
rect 64144 419432 64196 419484
rect 69112 419432 69164 419484
rect 15200 419364 15252 419416
rect 42800 419364 42852 419416
rect 62764 419364 62816 419416
rect 69756 419364 69808 419416
rect 96712 419432 96764 419484
rect 96804 419364 96856 419416
rect 200764 419432 200816 419484
rect 204628 419432 204680 419484
rect 251824 419432 251876 419484
rect 258724 419432 258776 419484
rect 443644 419432 443696 419484
rect 447692 419432 447744 419484
rect 494704 419432 494756 419484
rect 501604 419432 501656 419484
rect 123668 419364 123720 419416
rect 149704 419364 149756 419416
rect 547972 419364 548024 419416
rect 26056 419296 26108 419348
rect 36820 419296 36872 419348
rect 79968 419296 80020 419348
rect 90364 419296 90416 419348
rect 106556 419296 106608 419348
rect 116584 419296 116636 419348
rect 133788 419296 133840 419348
rect 144276 419296 144328 419348
rect 150532 419296 150584 419348
rect 178132 419296 178184 419348
rect 187976 419296 188028 419348
rect 199384 419296 199436 419348
rect 204352 419296 204404 419348
rect 231860 419296 231912 419348
rect 242072 419296 242124 419348
rect 253204 419296 253256 419348
rect 258172 419296 258224 419348
rect 122932 419228 122984 419280
rect 150716 419228 150768 419280
rect 160560 419228 160612 419280
rect 171784 419228 171836 419280
rect 215024 419228 215076 419280
rect 225604 419228 225656 419280
rect 268936 419228 268988 419280
rect 279424 419228 279476 419280
rect 285772 419296 285824 419348
rect 312636 419296 312688 419348
rect 322848 419296 322900 419348
rect 333244 419296 333296 419348
rect 339592 419296 339644 419348
rect 286140 419228 286192 419280
rect 295984 419228 296036 419280
rect 307024 419228 307076 419280
rect 350080 419228 350132 419280
rect 359556 419228 359608 419280
rect 365812 419296 365864 419348
rect 393596 419296 393648 419348
rect 366732 419228 366784 419280
rect 376576 419228 376628 419280
rect 387064 419228 387116 419280
rect 393412 419228 393464 419280
rect 420920 419296 420972 419348
rect 431040 419296 431092 419348
rect 442264 419296 442316 419348
rect 447232 419296 447284 419348
rect 474740 419296 474792 419348
rect 484952 419296 485004 419348
rect 496084 419296 496136 419348
rect 511908 419296 511960 419348
rect 522396 419296 522448 419348
rect 403992 419228 404044 419280
rect 414664 419228 414716 419280
rect 458088 419228 458140 419280
rect 468484 419228 468536 419280
rect 36636 419160 36688 419212
rect 538404 419160 538456 419212
rect 16304 416032 16356 416084
rect 528744 416032 528796 416084
rect 25964 415692 26016 415744
rect 149704 415692 149756 415744
rect 36728 415624 36780 415676
rect 52460 415624 52512 415676
rect 475384 415624 475436 415676
rect 494704 415624 494756 415676
rect 43352 415556 43404 415608
rect 62764 415556 62816 415608
rect 90456 415556 90508 415608
rect 106372 415556 106424 415608
rect 116492 415556 116544 415608
rect 133420 415556 133472 415608
rect 144276 415556 144328 415608
rect 160284 415556 160336 415608
rect 170496 415556 170548 415608
rect 187792 415556 187844 415608
rect 197544 415556 197596 415608
rect 214380 415556 214432 415608
rect 224500 415556 224552 415608
rect 241520 415556 241572 415608
rect 251456 415556 251508 415608
rect 268292 415556 268344 415608
rect 413468 415556 413520 415608
rect 430580 415556 430632 415608
rect 440516 415556 440568 415608
rect 457260 415556 457312 415608
rect 468576 415556 468628 415608
rect 484400 415556 484452 415608
rect 36820 415488 36872 415540
rect 62120 415488 62172 415540
rect 64144 415488 64196 415540
rect 89076 415488 89128 415540
rect 90364 415488 90416 415540
rect 115940 415488 115992 415540
rect 116584 415488 116636 415540
rect 142988 415488 143040 415540
rect 144184 415488 144236 415540
rect 170036 415488 170088 415540
rect 178408 415488 178460 415540
rect 200764 415488 200816 415540
rect 232320 415488 232372 415540
rect 251824 415488 251876 415540
rect 279516 415488 279568 415540
rect 295800 415488 295852 415540
rect 305644 415488 305696 415540
rect 322388 415488 322440 415540
rect 336004 415488 336056 415540
rect 349804 415488 349856 415540
rect 359648 415488 359700 415540
rect 376300 415488 376352 415540
rect 386512 415488 386564 415540
rect 403348 415488 403400 415540
rect 421288 415488 421340 415540
rect 445024 415488 445076 415540
rect 494520 415488 494572 415540
rect 511356 415488 511408 415540
rect 522304 415488 522356 415540
rect 538404 415488 538456 415540
rect 62488 415420 62540 415472
rect 79324 415420 79376 415472
rect 171784 415420 171836 415472
rect 197452 415420 197504 415472
rect 199384 415420 199436 415472
rect 223948 415420 224000 415472
rect 225604 415420 225656 415472
rect 251180 415420 251232 415472
rect 253204 415420 253256 415472
rect 278044 415420 278096 415472
rect 279424 415420 279476 415472
rect 305552 415420 305604 415472
rect 307024 415420 307076 415472
rect 331956 415420 332008 415472
rect 333244 415420 333296 415472
rect 359464 415420 359516 415472
rect 359740 415420 359792 415472
rect 386052 415420 386104 415472
rect 387064 415420 387116 415472
rect 412916 415420 412968 415472
rect 414664 415420 414716 415472
rect 440240 415420 440292 415472
rect 442264 415420 442316 415472
rect 467012 415420 467064 415472
rect 468484 415420 468536 415472
rect 494060 415420 494112 415472
rect 496084 415420 496136 415472
rect 520924 415420 520976 415472
rect 522396 415420 522448 415472
rect 548064 415420 548116 415472
rect 37924 414672 37976 414724
rect 526444 414672 526496 414724
rect 339592 413312 339644 413364
rect 340144 413312 340196 413364
rect 35624 412632 35676 412684
rect 36636 412632 36688 412684
rect 13728 394612 13780 394664
rect 64880 394612 64932 394664
rect 89720 394612 89772 394664
rect 90456 394612 90508 394664
rect 95148 394612 95200 394664
rect 143632 394612 143684 394664
rect 144276 394612 144328 394664
rect 445024 394680 445076 394732
rect 447692 394680 447744 394732
rect 146300 394612 146352 394664
rect 148968 394612 149020 394664
rect 200120 394612 200172 394664
rect 202788 394612 202840 394664
rect 253940 394612 253992 394664
rect 278688 394612 278740 394664
rect 279516 394612 279568 394664
rect 284208 394612 284260 394664
rect 335360 394612 335412 394664
rect 338028 394612 338080 394664
rect 389180 394612 389232 394664
rect 391848 394612 391900 394664
rect 443000 394612 443052 394664
rect 445668 394612 445720 394664
rect 496820 394612 496872 394664
rect 500868 394612 500920 394664
rect 550640 394612 550692 394664
rect 35624 394544 35676 394596
rect 36728 394544 36780 394596
rect 41328 394544 41380 394596
rect 91100 394544 91152 394596
rect 122748 394544 122800 394596
rect 172520 394544 172572 394596
rect 176568 394544 176620 394596
rect 226340 394544 226392 394596
rect 256608 394544 256660 394596
rect 307760 394544 307812 394596
rect 311808 394544 311860 394596
rect 361580 394544 361632 394596
rect 365628 394544 365680 394596
rect 415400 394544 415452 394596
rect 419448 394544 419500 394596
rect 68928 394476 68980 394528
rect 118700 394476 118752 394528
rect 230388 394476 230440 394528
rect 280160 394476 280212 394528
rect 332600 394476 332652 394528
rect 336004 394476 336056 394528
rect 467656 394544 467708 394596
rect 468576 394544 468628 394596
rect 473268 394544 473320 394596
rect 523040 394544 523092 394596
rect 469220 394476 469272 394528
rect 52736 391892 52788 391944
rect 64144 391892 64196 391944
rect 69112 391892 69164 391944
rect 15200 391824 15252 391876
rect 42984 391824 43036 391876
rect 62764 391824 62816 391876
rect 70032 391824 70084 391876
rect 96712 391892 96764 391944
rect 96988 391824 97040 391876
rect 200764 391892 200816 391944
rect 204996 391892 205048 391944
rect 251824 391892 251876 391944
rect 259000 391892 259052 391944
rect 494704 391892 494756 391944
rect 501972 391892 502024 391944
rect 124036 391824 124088 391876
rect 133696 391824 133748 391876
rect 144184 391824 144236 391876
rect 146944 391824 146996 391876
rect 548340 391824 548392 391876
rect 25688 391756 25740 391808
rect 36820 391756 36872 391808
rect 79692 391756 79744 391808
rect 90364 391756 90416 391808
rect 106648 391756 106700 391808
rect 116584 391756 116636 391808
rect 122932 391756 122984 391808
rect 150532 391756 150584 391808
rect 178040 391756 178092 391808
rect 187700 391756 187752 391808
rect 199384 391756 199436 391808
rect 204352 391756 204404 391808
rect 232044 391756 232096 391808
rect 241704 391756 241756 391808
rect 253204 391756 253256 391808
rect 258172 391756 258224 391808
rect 150992 391688 151044 391740
rect 160652 391688 160704 391740
rect 171784 391688 171836 391740
rect 214656 391688 214708 391740
rect 225604 391688 225656 391740
rect 268660 391688 268712 391740
rect 279424 391688 279476 391740
rect 285772 391756 285824 391808
rect 313004 391756 313056 391808
rect 286048 391688 286100 391740
rect 295708 391688 295760 391740
rect 307024 391688 307076 391740
rect 311992 391688 312044 391740
rect 340052 391756 340104 391808
rect 322664 391688 322716 391740
rect 333244 391688 333296 391740
rect 339592 391688 339644 391740
rect 366732 391756 366784 391808
rect 349712 391688 349764 391740
rect 359556 391688 359608 391740
rect 365812 391688 365864 391740
rect 393964 391756 394016 391808
rect 376668 391688 376720 391740
rect 387064 391688 387116 391740
rect 393412 391688 393464 391740
rect 421012 391756 421064 391808
rect 430672 391756 430724 391808
rect 442264 391756 442316 391808
rect 447232 391756 447284 391808
rect 475016 391756 475068 391808
rect 484676 391756 484728 391808
rect 496084 391756 496136 391808
rect 501052 391756 501104 391808
rect 529020 391756 529072 391808
rect 403716 391688 403768 391740
rect 414664 391688 414716 391740
rect 457720 391688 457772 391740
rect 468484 391688 468536 391740
rect 511724 391688 511776 391740
rect 522396 391688 522448 391740
rect 36544 391620 36596 391672
rect 538680 391620 538732 391672
rect 16028 389784 16080 389836
rect 528744 389784 528796 389836
rect 25964 389444 26016 389496
rect 146944 389444 146996 389496
rect 36820 389376 36872 389428
rect 52460 389376 52512 389428
rect 232320 389376 232372 389428
rect 251824 389376 251876 389428
rect 475384 389376 475436 389428
rect 494704 389376 494756 389428
rect 43352 389308 43404 389360
rect 62764 389308 62816 389360
rect 90456 389308 90508 389360
rect 106372 389308 106424 389360
rect 116492 389308 116544 389360
rect 133420 389308 133472 389360
rect 170496 389308 170548 389360
rect 187792 389308 187844 389360
rect 197544 389308 197596 389360
rect 214380 389308 214432 389360
rect 224500 389308 224552 389360
rect 241520 389308 241572 389360
rect 413468 389308 413520 389360
rect 430580 389308 430632 389360
rect 440516 389308 440568 389360
rect 457260 389308 457312 389360
rect 468576 389308 468628 389360
rect 484400 389308 484452 389360
rect 36728 389240 36780 389292
rect 62120 389240 62172 389292
rect 64144 389240 64196 389292
rect 89076 389240 89128 389292
rect 90364 389240 90416 389292
rect 115940 389240 115992 389292
rect 116584 389240 116636 389292
rect 142988 389240 143040 389292
rect 144276 389240 144328 389292
rect 170036 389240 170088 389292
rect 178408 389240 178460 389292
rect 200764 389240 200816 389292
rect 251456 389240 251508 389292
rect 268292 389240 268344 389292
rect 279424 389240 279476 389292
rect 295800 389240 295852 389292
rect 305644 389240 305696 389292
rect 322388 389240 322440 389292
rect 336004 389240 336056 389292
rect 349804 389240 349856 389292
rect 359556 389240 359608 389292
rect 376300 389240 376352 389292
rect 386512 389240 386564 389292
rect 403348 389240 403400 389292
rect 421288 389240 421340 389292
rect 446404 389240 446456 389292
rect 494520 389240 494572 389292
rect 511356 389240 511408 389292
rect 522304 389240 522356 389292
rect 538404 389240 538456 389292
rect 62488 389172 62540 389224
rect 79324 389172 79376 389224
rect 144184 389172 144236 389224
rect 160284 389172 160336 389224
rect 171784 389172 171836 389224
rect 197452 389172 197504 389224
rect 199384 389172 199436 389224
rect 223948 389172 224000 389224
rect 225604 389172 225656 389224
rect 251180 389172 251232 389224
rect 253204 389172 253256 389224
rect 278044 389172 278096 389224
rect 279516 389172 279568 389224
rect 305552 389172 305604 389224
rect 307024 389172 307076 389224
rect 331956 389172 332008 389224
rect 333244 389172 333296 389224
rect 359464 389172 359516 389224
rect 359740 389172 359792 389224
rect 386052 389172 386104 389224
rect 387064 389172 387116 389224
rect 412916 389172 412968 389224
rect 414664 389172 414716 389224
rect 440240 389172 440292 389224
rect 442264 389172 442316 389224
rect 467012 389172 467064 389224
rect 468484 389172 468536 389224
rect 494060 389172 494112 389224
rect 496084 389172 496136 389224
rect 520924 389172 520976 389224
rect 522396 389172 522448 389224
rect 548064 389172 548116 389224
rect 37924 387064 37976 387116
rect 526444 387064 526496 387116
rect 285772 386248 285824 386300
rect 286140 386248 286192 386300
rect 339592 386248 339644 386300
rect 340144 386248 340196 386300
rect 89720 370540 89772 370592
rect 90456 370540 90508 370592
rect 13728 368432 13780 368484
rect 64880 368432 64932 368484
rect 95148 368432 95200 368484
rect 144828 368432 144880 368484
rect 148968 368432 149020 368484
rect 200120 368432 200172 368484
rect 202788 368432 202840 368484
rect 253940 368432 253992 368484
rect 284208 368432 284260 368484
rect 335360 368432 335412 368484
rect 338028 368432 338080 368484
rect 389180 368432 389232 368484
rect 391848 368432 391900 368484
rect 443000 368432 443052 368484
rect 446404 368432 446456 368484
rect 447692 368432 447744 368484
rect 41328 368364 41380 368416
rect 91100 368364 91152 368416
rect 122748 368364 122800 368416
rect 172520 368364 172572 368416
rect 176568 368364 176620 368416
rect 226340 368364 226392 368416
rect 256608 368364 256660 368416
rect 307760 368364 307812 368416
rect 311808 368364 311860 368416
rect 361580 368364 361632 368416
rect 365628 368364 365680 368416
rect 415400 368364 415452 368416
rect 419448 368364 419500 368416
rect 68928 368296 68980 368348
rect 118700 368296 118752 368348
rect 230388 368296 230440 368348
rect 280160 368296 280212 368348
rect 445668 368296 445720 368348
rect 496820 368432 496872 368484
rect 500868 368432 500920 368484
rect 550640 368432 550692 368484
rect 469220 368364 469272 368416
rect 473268 368364 473320 368416
rect 523040 368364 523092 368416
rect 467656 368296 467708 368348
rect 468576 368296 468628 368348
rect 170220 367616 170272 367668
rect 170496 367616 170548 367668
rect 35624 367004 35676 367056
rect 36820 367004 36872 367056
rect 53104 365644 53156 365696
rect 64144 365644 64196 365696
rect 69112 365644 69164 365696
rect 15200 365576 15252 365628
rect 42800 365576 42852 365628
rect 62764 365576 62816 365628
rect 69756 365576 69808 365628
rect 96712 365644 96764 365696
rect 96804 365576 96856 365628
rect 200764 365644 200816 365696
rect 204628 365644 204680 365696
rect 251824 365644 251876 365696
rect 258724 365644 258776 365696
rect 332508 365644 332560 365696
rect 336004 365644 336056 365696
rect 494704 365644 494756 365696
rect 501604 365644 501656 365696
rect 123668 365576 123720 365628
rect 149704 365576 149756 365628
rect 548064 365576 548116 365628
rect 26056 365508 26108 365560
rect 36728 365508 36780 365560
rect 79968 365508 80020 365560
rect 90364 365508 90416 365560
rect 106556 365508 106608 365560
rect 116584 365508 116636 365560
rect 133788 365508 133840 365560
rect 144276 365508 144328 365560
rect 150532 365508 150584 365560
rect 178132 365508 178184 365560
rect 187976 365508 188028 365560
rect 199384 365508 199436 365560
rect 204352 365508 204404 365560
rect 231860 365508 231912 365560
rect 242072 365508 242124 365560
rect 253204 365508 253256 365560
rect 258172 365508 258224 365560
rect 286140 365508 286192 365560
rect 122932 365440 122984 365492
rect 150716 365440 150768 365492
rect 160560 365440 160612 365492
rect 171784 365440 171836 365492
rect 215024 365440 215076 365492
rect 225604 365440 225656 365492
rect 268936 365440 268988 365492
rect 279516 365440 279568 365492
rect 285772 365440 285824 365492
rect 312636 365508 312688 365560
rect 295984 365440 296036 365492
rect 307024 365440 307076 365492
rect 311992 365440 312044 365492
rect 340144 365508 340196 365560
rect 322848 365440 322900 365492
rect 333244 365440 333296 365492
rect 339592 365440 339644 365492
rect 366732 365508 366784 365560
rect 350080 365440 350132 365492
rect 359556 365440 359608 365492
rect 365812 365440 365864 365492
rect 393596 365508 393648 365560
rect 376576 365440 376628 365492
rect 387064 365440 387116 365492
rect 393412 365440 393464 365492
rect 420920 365508 420972 365560
rect 431040 365508 431092 365560
rect 442264 365508 442316 365560
rect 447232 365508 447284 365560
rect 474740 365508 474792 365560
rect 484952 365508 485004 365560
rect 496084 365508 496136 365560
rect 501052 365508 501104 365560
rect 528652 365508 528704 365560
rect 403992 365440 404044 365492
rect 414664 365440 414716 365492
rect 458088 365440 458140 365492
rect 468484 365440 468536 365492
rect 511908 365440 511960 365492
rect 522396 365440 522448 365492
rect 36636 365372 36688 365424
rect 538404 365372 538456 365424
rect 16120 362176 16172 362228
rect 529020 362176 529072 362228
rect 25688 361836 25740 361888
rect 149704 361836 149756 361888
rect 36820 361768 36872 361820
rect 52644 361768 52696 361820
rect 232044 361768 232096 361820
rect 251824 361768 251876 361820
rect 475016 361768 475068 361820
rect 494704 361768 494756 361820
rect 62488 361700 62540 361752
rect 79692 361700 79744 361752
rect 90364 361700 90416 361752
rect 106648 361700 106700 361752
rect 116492 361700 116544 361752
rect 133696 361700 133748 361752
rect 144276 361700 144328 361752
rect 160652 361700 160704 361752
rect 170496 361700 170548 361752
rect 187700 361700 187752 361752
rect 197452 361700 197504 361752
rect 214656 361700 214708 361752
rect 224500 361700 224552 361752
rect 241704 361700 241756 361752
rect 413468 361700 413520 361752
rect 430672 361700 430724 361752
rect 440516 361700 440568 361752
rect 457628 361700 457680 361752
rect 468576 361700 468628 361752
rect 484676 361700 484728 361752
rect 36636 361632 36688 361684
rect 62304 361632 62356 361684
rect 64144 361632 64196 361684
rect 89352 361632 89404 361684
rect 90456 361632 90508 361684
rect 116308 361632 116360 361684
rect 116584 361632 116636 361684
rect 143356 361632 143408 361684
rect 144184 361632 144236 361684
rect 170312 361632 170364 361684
rect 178040 361632 178092 361684
rect 200764 361632 200816 361684
rect 251456 361632 251508 361684
rect 268660 361632 268712 361684
rect 279516 361632 279568 361684
rect 295708 361632 295760 361684
rect 305460 361632 305512 361684
rect 322664 361632 322716 361684
rect 334624 361632 334676 361684
rect 349712 361632 349764 361684
rect 359464 361632 359516 361684
rect 376668 361632 376720 361684
rect 386512 361632 386564 361684
rect 403624 361632 403676 361684
rect 421012 361632 421064 361684
rect 443644 361632 443696 361684
rect 494520 361632 494572 361684
rect 511632 361632 511684 361684
rect 522304 361632 522356 361684
rect 538680 361632 538732 361684
rect 43076 361564 43128 361616
rect 62764 361564 62816 361616
rect 171784 361564 171836 361616
rect 197360 361564 197412 361616
rect 199384 361564 199436 361616
rect 224316 361564 224368 361616
rect 225604 361564 225656 361616
rect 251364 361564 251416 361616
rect 253204 361564 253256 361616
rect 278320 361564 278372 361616
rect 279424 361564 279476 361616
rect 305368 361564 305420 361616
rect 307024 361564 307076 361616
rect 332324 361564 332376 361616
rect 333244 361564 333296 361616
rect 359372 361564 359424 361616
rect 359556 361564 359608 361616
rect 386328 361564 386380 361616
rect 387064 361564 387116 361616
rect 413284 361564 413336 361616
rect 414664 361564 414716 361616
rect 440332 361564 440384 361616
rect 442264 361564 442316 361616
rect 467288 361564 467340 361616
rect 468484 361564 468536 361616
rect 494336 361564 494388 361616
rect 496084 361564 496136 361616
rect 521292 361564 521344 361616
rect 522396 361564 522448 361616
rect 548340 361564 548392 361616
rect 37924 359456 37976 359508
rect 526444 359456 526496 359508
rect 35624 358776 35676 358828
rect 36728 358776 36780 358828
rect 143632 342524 143684 342576
rect 144276 342524 144328 342576
rect 443644 340892 443696 340944
rect 447692 340892 447744 340944
rect 13728 340824 13780 340876
rect 64880 340824 64932 340876
rect 95148 340824 95200 340876
rect 146300 340824 146352 340876
rect 148968 340824 149020 340876
rect 200120 340824 200172 340876
rect 202788 340824 202840 340876
rect 253940 340824 253992 340876
rect 256608 340824 256660 340876
rect 307760 340824 307812 340876
rect 332508 340824 332560 340876
rect 334624 340824 334676 340876
rect 338028 340824 338080 340876
rect 389180 340824 389232 340876
rect 391848 340824 391900 340876
rect 443000 340824 443052 340876
rect 445668 340824 445720 340876
rect 496820 340824 496872 340876
rect 500868 340824 500920 340876
rect 550640 340824 550692 340876
rect 35624 340756 35676 340808
rect 36820 340756 36872 340808
rect 41328 340756 41380 340808
rect 91100 340756 91152 340808
rect 122748 340756 122800 340808
rect 172520 340756 172572 340808
rect 176568 340756 176620 340808
rect 226340 340756 226392 340808
rect 230388 340756 230440 340808
rect 280160 340756 280212 340808
rect 284208 340756 284260 340808
rect 335360 340756 335412 340808
rect 365628 340756 365680 340808
rect 415400 340756 415452 340808
rect 419448 340756 419500 340808
rect 469220 340756 469272 340808
rect 473268 340756 473320 340808
rect 523040 340756 523092 340808
rect 68928 340688 68980 340740
rect 118700 340688 118752 340740
rect 200764 340688 200816 340740
rect 204628 340688 204680 340740
rect 278688 340688 278740 340740
rect 279516 340688 279568 340740
rect 311808 340688 311860 340740
rect 361580 340688 361632 340740
rect 467656 340688 467708 340740
rect 468576 340688 468628 340740
rect 25688 338036 25740 338088
rect 36636 338036 36688 338088
rect 52736 338036 52788 338088
rect 64144 338036 64196 338088
rect 69112 338036 69164 338088
rect 15200 337968 15252 338020
rect 42984 337968 43036 338020
rect 62764 337968 62816 338020
rect 70032 337968 70084 338020
rect 96712 338036 96764 338088
rect 96988 337968 97040 338020
rect 146944 338036 146996 338088
rect 124036 337968 124088 338020
rect 133696 337968 133748 338020
rect 144184 337968 144236 338020
rect 150532 337968 150584 338020
rect 251824 338036 251876 338088
rect 259000 338036 259052 338088
rect 494704 338036 494756 338088
rect 501972 338036 502024 338088
rect 79692 337900 79744 337952
rect 90456 337900 90508 337952
rect 106648 337900 106700 337952
rect 116584 337900 116636 337952
rect 122932 337900 122984 337952
rect 150992 337900 151044 337952
rect 548340 337968 548392 338020
rect 178040 337900 178092 337952
rect 187700 337900 187752 337952
rect 199384 337900 199436 337952
rect 204352 337900 204404 337952
rect 232044 337900 232096 337952
rect 241704 337900 241756 337952
rect 253204 337900 253256 337952
rect 258172 337900 258224 337952
rect 286048 337900 286100 337952
rect 160652 337832 160704 337884
rect 171784 337832 171836 337884
rect 214656 337832 214708 337884
rect 225604 337832 225656 337884
rect 268660 337832 268712 337884
rect 279424 337832 279476 337884
rect 285772 337832 285824 337884
rect 313004 337900 313056 337952
rect 295708 337832 295760 337884
rect 307024 337832 307076 337884
rect 311992 337832 312044 337884
rect 340052 337900 340104 337952
rect 322664 337832 322716 337884
rect 333244 337832 333296 337884
rect 339592 337832 339644 337884
rect 367008 337900 367060 337952
rect 349712 337832 349764 337884
rect 359556 337832 359608 337884
rect 365812 337832 365864 337884
rect 393964 337900 394016 337952
rect 376668 337832 376720 337884
rect 387064 337832 387116 337884
rect 393412 337832 393464 337884
rect 421012 337900 421064 337952
rect 430672 337900 430724 337952
rect 442264 337900 442316 337952
rect 447232 337900 447284 337952
rect 475016 337900 475068 337952
rect 484676 337900 484728 337952
rect 496084 337900 496136 337952
rect 501052 337900 501104 337952
rect 529020 337900 529072 337952
rect 403716 337832 403768 337884
rect 414664 337832 414716 337884
rect 457720 337832 457772 337884
rect 468484 337832 468536 337884
rect 511724 337832 511776 337884
rect 522396 337832 522448 337884
rect 36544 337764 36596 337816
rect 538680 337764 538732 337816
rect 16028 335996 16080 336048
rect 528652 335996 528704 336048
rect 26056 335588 26108 335640
rect 146944 335588 146996 335640
rect 36544 335520 36596 335572
rect 52460 335520 52512 335572
rect 232320 335520 232372 335572
rect 251824 335520 251876 335572
rect 475384 335520 475436 335572
rect 494704 335520 494756 335572
rect 62488 335452 62540 335504
rect 79324 335452 79376 335504
rect 90456 335452 90508 335504
rect 106464 335452 106516 335504
rect 116492 335452 116544 335504
rect 133420 335452 133472 335504
rect 170496 335452 170548 335504
rect 187792 335452 187844 335504
rect 197544 335452 197596 335504
rect 214380 335452 214432 335504
rect 224500 335452 224552 335504
rect 241612 335452 241664 335504
rect 413468 335452 413520 335504
rect 430580 335452 430632 335504
rect 440516 335452 440568 335504
rect 457260 335452 457312 335504
rect 468484 335452 468536 335504
rect 484400 335452 484452 335504
rect 36820 335384 36872 335436
rect 62120 335384 62172 335436
rect 64144 335384 64196 335436
rect 89076 335384 89128 335436
rect 90364 335384 90416 335436
rect 116124 335384 116176 335436
rect 116584 335384 116636 335436
rect 142988 335384 143040 335436
rect 144276 335384 144328 335436
rect 170036 335384 170088 335436
rect 178408 335384 178460 335436
rect 200764 335384 200816 335436
rect 251456 335384 251508 335436
rect 268292 335384 268344 335436
rect 279516 335384 279568 335436
rect 295800 335384 295852 335436
rect 305552 335384 305604 335436
rect 322388 335384 322440 335436
rect 336004 335384 336056 335436
rect 349804 335384 349856 335436
rect 359648 335384 359700 335436
rect 376300 335384 376352 335436
rect 386512 335384 386564 335436
rect 403348 335384 403400 335436
rect 421288 335384 421340 335436
rect 446404 335384 446456 335436
rect 494520 335384 494572 335436
rect 511356 335384 511408 335436
rect 522304 335384 522356 335436
rect 538404 335384 538456 335436
rect 43352 335316 43404 335368
rect 62764 335316 62816 335368
rect 144184 335316 144236 335368
rect 160284 335316 160336 335368
rect 171784 335316 171836 335368
rect 197452 335316 197504 335368
rect 199384 335316 199436 335368
rect 223948 335316 224000 335368
rect 225604 335316 225656 335368
rect 251272 335316 251324 335368
rect 253204 335316 253256 335368
rect 278044 335316 278096 335368
rect 279424 335316 279476 335368
rect 305460 335316 305512 335368
rect 307024 335316 307076 335368
rect 331956 335316 332008 335368
rect 333244 335316 333296 335368
rect 359464 335316 359516 335368
rect 359556 335316 359608 335368
rect 386052 335316 386104 335368
rect 387064 335316 387116 335368
rect 412916 335316 412968 335368
rect 414664 335316 414716 335368
rect 440240 335316 440292 335368
rect 442264 335316 442316 335368
rect 467012 335316 467064 335368
rect 468576 335316 468628 335368
rect 494060 335316 494112 335368
rect 496084 335316 496136 335368
rect 520924 335316 520976 335368
rect 522396 335316 522448 335368
rect 547972 335316 548024 335368
rect 37924 333208 37976 333260
rect 526444 333208 526496 333260
rect 35624 332528 35676 332580
rect 36636 332528 36688 332580
rect 285772 332256 285824 332308
rect 286140 332256 286192 332308
rect 339592 332256 339644 332308
rect 340144 332256 340196 332308
rect 359556 330624 359608 330676
rect 359556 330420 359608 330472
rect 445668 314644 445720 314696
rect 13728 314576 13780 314628
rect 64880 314576 64932 314628
rect 89720 314576 89772 314628
rect 90456 314576 90508 314628
rect 95148 314576 95200 314628
rect 146300 314576 146352 314628
rect 148968 314576 149020 314628
rect 200120 314576 200172 314628
rect 202788 314576 202840 314628
rect 253940 314576 253992 314628
rect 256608 314576 256660 314628
rect 307760 314576 307812 314628
rect 338028 314576 338080 314628
rect 389180 314576 389232 314628
rect 391848 314576 391900 314628
rect 443000 314576 443052 314628
rect 446404 314576 446456 314628
rect 447692 314576 447744 314628
rect 496820 314576 496872 314628
rect 500868 314576 500920 314628
rect 550640 314576 550692 314628
rect 41328 314508 41380 314560
rect 91100 314508 91152 314560
rect 122748 314508 122800 314560
rect 172520 314508 172572 314560
rect 176568 314508 176620 314560
rect 226340 314508 226392 314560
rect 230388 314508 230440 314560
rect 280160 314508 280212 314560
rect 284208 314508 284260 314560
rect 335360 314508 335412 314560
rect 365628 314508 365680 314560
rect 415400 314508 415452 314560
rect 419448 314508 419500 314560
rect 68928 314440 68980 314492
rect 118700 314440 118752 314492
rect 278688 314440 278740 314492
rect 279516 314440 279568 314492
rect 311808 314440 311860 314492
rect 361580 314440 361632 314492
rect 469220 314508 469272 314560
rect 473268 314508 473320 314560
rect 523040 314508 523092 314560
rect 170220 313624 170272 313676
rect 170496 313624 170548 313676
rect 62764 311788 62816 311840
rect 69756 311788 69808 311840
rect 96712 311788 96764 311840
rect 15200 311720 15252 311772
rect 42800 311720 42852 311772
rect 53104 311720 53156 311772
rect 64144 311720 64196 311772
rect 69112 311720 69164 311772
rect 96804 311720 96856 311772
rect 200764 311788 200816 311840
rect 204628 311788 204680 311840
rect 251824 311788 251876 311840
rect 258724 311788 258776 311840
rect 332508 311788 332560 311840
rect 336004 311788 336056 311840
rect 494704 311788 494756 311840
rect 501604 311788 501656 311840
rect 123668 311720 123720 311772
rect 149704 311720 149756 311772
rect 548064 311720 548116 311772
rect 25964 311652 26016 311704
rect 36820 311652 36872 311704
rect 79968 311652 80020 311704
rect 90364 311652 90416 311704
rect 106556 311652 106608 311704
rect 116584 311652 116636 311704
rect 133788 311652 133840 311704
rect 144276 311652 144328 311704
rect 150532 311652 150584 311704
rect 178132 311652 178184 311704
rect 187976 311652 188028 311704
rect 199384 311652 199436 311704
rect 204352 311652 204404 311704
rect 231860 311652 231912 311704
rect 242072 311652 242124 311704
rect 253204 311652 253256 311704
rect 258172 311652 258224 311704
rect 286140 311652 286192 311704
rect 122932 311584 122984 311636
rect 150716 311584 150768 311636
rect 160560 311584 160612 311636
rect 171784 311584 171836 311636
rect 215024 311584 215076 311636
rect 225604 311584 225656 311636
rect 268936 311584 268988 311636
rect 279424 311584 279476 311636
rect 285772 311584 285824 311636
rect 312636 311652 312688 311704
rect 295984 311584 296036 311636
rect 307024 311584 307076 311636
rect 311992 311584 312044 311636
rect 340144 311652 340196 311704
rect 322848 311584 322900 311636
rect 333244 311584 333296 311636
rect 339592 311584 339644 311636
rect 366732 311652 366784 311704
rect 350080 311584 350132 311636
rect 359556 311584 359608 311636
rect 365812 311584 365864 311636
rect 393596 311652 393648 311704
rect 376576 311584 376628 311636
rect 387064 311584 387116 311636
rect 393412 311584 393464 311636
rect 420920 311652 420972 311704
rect 431040 311652 431092 311704
rect 442264 311652 442316 311704
rect 447232 311652 447284 311704
rect 474740 311652 474792 311704
rect 484952 311652 485004 311704
rect 496084 311652 496136 311704
rect 501052 311652 501104 311704
rect 528744 311652 528796 311704
rect 403992 311584 404044 311636
rect 414664 311584 414716 311636
rect 458088 311584 458140 311636
rect 468576 311584 468628 311636
rect 511908 311584 511960 311636
rect 522396 311584 522448 311636
rect 36728 311516 36780 311568
rect 538404 311516 538456 311568
rect 16304 308388 16356 308440
rect 529020 308388 529072 308440
rect 25688 308048 25740 308100
rect 149704 308048 149756 308100
rect 36820 307980 36872 308032
rect 52644 307980 52696 308032
rect 232044 307980 232096 308032
rect 251824 307980 251876 308032
rect 475016 307980 475068 308032
rect 494704 307980 494756 308032
rect 62488 307912 62540 307964
rect 79692 307912 79744 307964
rect 90364 307912 90416 307964
rect 106648 307912 106700 307964
rect 116492 307912 116544 307964
rect 133696 307912 133748 307964
rect 144184 307912 144236 307964
rect 160652 307912 160704 307964
rect 170496 307912 170548 307964
rect 187700 307912 187752 307964
rect 197452 307912 197504 307964
rect 214656 307912 214708 307964
rect 224500 307912 224552 307964
rect 241704 307912 241756 307964
rect 413468 307912 413520 307964
rect 430672 307912 430724 307964
rect 440516 307912 440568 307964
rect 457628 307912 457680 307964
rect 468576 307912 468628 307964
rect 484676 307912 484728 307964
rect 36728 307844 36780 307896
rect 62304 307844 62356 307896
rect 64144 307844 64196 307896
rect 89352 307844 89404 307896
rect 90456 307844 90508 307896
rect 116308 307844 116360 307896
rect 116584 307844 116636 307896
rect 143356 307844 143408 307896
rect 144276 307844 144328 307896
rect 170312 307844 170364 307896
rect 178040 307844 178092 307896
rect 200764 307844 200816 307896
rect 251456 307844 251508 307896
rect 268660 307844 268712 307896
rect 279516 307844 279568 307896
rect 295708 307844 295760 307896
rect 305460 307844 305512 307896
rect 322664 307844 322716 307896
rect 334624 307844 334676 307896
rect 349712 307844 349764 307896
rect 359464 307844 359516 307896
rect 376668 307844 376720 307896
rect 386512 307844 386564 307896
rect 403624 307844 403676 307896
rect 421012 307844 421064 307896
rect 443644 307844 443696 307896
rect 494520 307844 494572 307896
rect 511632 307844 511684 307896
rect 522304 307844 522356 307896
rect 538680 307844 538732 307896
rect 43076 307776 43128 307828
rect 62764 307776 62816 307828
rect 171784 307776 171836 307828
rect 197360 307776 197412 307828
rect 199384 307776 199436 307828
rect 224316 307776 224368 307828
rect 225604 307776 225656 307828
rect 251364 307776 251416 307828
rect 253204 307776 253256 307828
rect 278320 307776 278372 307828
rect 279424 307776 279476 307828
rect 305368 307776 305420 307828
rect 307024 307776 307076 307828
rect 332324 307776 332376 307828
rect 333244 307776 333296 307828
rect 359372 307776 359424 307828
rect 359556 307776 359608 307828
rect 386328 307776 386380 307828
rect 387064 307776 387116 307828
rect 413284 307776 413336 307828
rect 414664 307776 414716 307828
rect 440332 307776 440384 307828
rect 442264 307776 442316 307828
rect 467288 307776 467340 307828
rect 468484 307776 468536 307828
rect 494336 307776 494388 307828
rect 496084 307776 496136 307828
rect 521292 307776 521344 307828
rect 522396 307776 522448 307828
rect 548340 307776 548392 307828
rect 37924 305600 37976 305652
rect 526444 305600 526496 305652
rect 13728 286968 13780 287020
rect 64880 286968 64932 287020
rect 95148 286968 95200 287020
rect 146300 286968 146352 287020
rect 148968 286968 149020 287020
rect 200120 286968 200172 287020
rect 202788 286968 202840 287020
rect 253940 286968 253992 287020
rect 256608 286968 256660 287020
rect 307760 286968 307812 287020
rect 338028 286968 338080 287020
rect 389180 286968 389232 287020
rect 391848 286968 391900 287020
rect 443000 286968 443052 287020
rect 445668 286968 445720 287020
rect 496820 286968 496872 287020
rect 500868 286968 500920 287020
rect 550640 286968 550692 287020
rect 35624 286900 35676 286952
rect 36820 286900 36872 286952
rect 41328 286900 41380 286952
rect 91100 286900 91152 286952
rect 122748 286900 122800 286952
rect 172520 286900 172572 286952
rect 176568 286900 176620 286952
rect 226340 286900 226392 286952
rect 230388 286900 230440 286952
rect 280160 286900 280212 286952
rect 284208 286900 284260 286952
rect 335360 286900 335412 286952
rect 365628 286900 365680 286952
rect 415400 286900 415452 286952
rect 419448 286900 419500 286952
rect 469220 286900 469272 286952
rect 473268 286900 473320 286952
rect 523040 286900 523092 286952
rect 68928 286832 68980 286884
rect 118700 286832 118752 286884
rect 311808 286832 311860 286884
rect 361580 286832 361632 286884
rect 200764 286764 200816 286816
rect 204628 286764 204680 286816
rect 278688 286764 278740 286816
rect 279516 286764 279568 286816
rect 332508 286764 332560 286816
rect 334624 286764 334676 286816
rect 467656 286764 467708 286816
rect 468576 286764 468628 286816
rect 62764 284248 62816 284300
rect 70032 284248 70084 284300
rect 96712 284248 96764 284300
rect 15200 284180 15252 284232
rect 42984 284180 43036 284232
rect 52736 284180 52788 284232
rect 64144 284180 64196 284232
rect 69112 284180 69164 284232
rect 96988 284180 97040 284232
rect 146944 284248 146996 284300
rect 124036 284180 124088 284232
rect 133696 284180 133748 284232
rect 144276 284180 144328 284232
rect 150532 284180 150584 284232
rect 251824 284248 251876 284300
rect 259000 284248 259052 284300
rect 443644 284248 443696 284300
rect 447968 284248 448020 284300
rect 494704 284248 494756 284300
rect 501972 284248 502024 284300
rect 25688 284112 25740 284164
rect 36728 284112 36780 284164
rect 79692 284112 79744 284164
rect 90456 284112 90508 284164
rect 106648 284112 106700 284164
rect 116584 284112 116636 284164
rect 122932 284112 122984 284164
rect 150992 284112 151044 284164
rect 548340 284180 548392 284232
rect 178040 284112 178092 284164
rect 187700 284112 187752 284164
rect 199384 284112 199436 284164
rect 204352 284112 204404 284164
rect 232044 284112 232096 284164
rect 241704 284112 241756 284164
rect 253204 284112 253256 284164
rect 258172 284112 258224 284164
rect 286048 284112 286100 284164
rect 160652 284044 160704 284096
rect 171784 284044 171836 284096
rect 214656 284044 214708 284096
rect 225604 284044 225656 284096
rect 268660 284044 268712 284096
rect 279424 284044 279476 284096
rect 285772 284044 285824 284096
rect 313004 284112 313056 284164
rect 295708 284044 295760 284096
rect 307024 284044 307076 284096
rect 311992 284044 312044 284096
rect 340052 284112 340104 284164
rect 322664 284044 322716 284096
rect 333244 284044 333296 284096
rect 339592 284044 339644 284096
rect 367008 284112 367060 284164
rect 349712 284044 349764 284096
rect 359556 284044 359608 284096
rect 365812 284044 365864 284096
rect 393964 284112 394016 284164
rect 376668 284044 376720 284096
rect 387064 284044 387116 284096
rect 393412 284044 393464 284096
rect 421012 284112 421064 284164
rect 430672 284112 430724 284164
rect 442264 284112 442316 284164
rect 447232 284112 447284 284164
rect 475016 284112 475068 284164
rect 484676 284112 484728 284164
rect 496084 284112 496136 284164
rect 501052 284112 501104 284164
rect 529020 284112 529072 284164
rect 403716 284044 403768 284096
rect 414664 284044 414716 284096
rect 457720 284044 457772 284096
rect 468484 284044 468536 284096
rect 511724 284044 511776 284096
rect 522396 284044 522448 284096
rect 36636 283976 36688 284028
rect 538680 283976 538732 284028
rect 16028 280780 16080 280832
rect 528744 280780 528796 280832
rect 25964 280440 26016 280492
rect 146944 280440 146996 280492
rect 36820 280372 36872 280424
rect 52460 280372 52512 280424
rect 232320 280372 232372 280424
rect 251824 280372 251876 280424
rect 475384 280372 475436 280424
rect 494704 280372 494756 280424
rect 62488 280304 62540 280356
rect 79324 280304 79376 280356
rect 90364 280304 90416 280356
rect 106372 280304 106424 280356
rect 116492 280304 116544 280356
rect 133420 280304 133472 280356
rect 170496 280304 170548 280356
rect 187792 280304 187844 280356
rect 197544 280304 197596 280356
rect 214380 280304 214432 280356
rect 224500 280304 224552 280356
rect 241520 280304 241572 280356
rect 413468 280304 413520 280356
rect 430580 280304 430632 280356
rect 440516 280304 440568 280356
rect 457260 280304 457312 280356
rect 468576 280304 468628 280356
rect 484400 280304 484452 280356
rect 36728 280236 36780 280288
rect 62120 280236 62172 280288
rect 64144 280236 64196 280288
rect 89076 280236 89128 280288
rect 90456 280236 90508 280288
rect 115940 280236 115992 280288
rect 116584 280236 116636 280288
rect 142988 280236 143040 280288
rect 144276 280236 144328 280288
rect 170036 280236 170088 280288
rect 178408 280236 178460 280288
rect 200764 280236 200816 280288
rect 251456 280236 251508 280288
rect 268292 280236 268344 280288
rect 279516 280236 279568 280288
rect 295800 280236 295852 280288
rect 305552 280236 305604 280288
rect 322388 280236 322440 280288
rect 336004 280236 336056 280288
rect 349804 280236 349856 280288
rect 359648 280236 359700 280288
rect 376300 280236 376352 280288
rect 386512 280236 386564 280288
rect 403348 280236 403400 280288
rect 421288 280236 421340 280288
rect 446404 280236 446456 280288
rect 494520 280236 494572 280288
rect 511356 280236 511408 280288
rect 522304 280236 522356 280288
rect 538404 280236 538456 280288
rect 43352 280168 43404 280220
rect 62764 280168 62816 280220
rect 144184 280168 144236 280220
rect 160284 280168 160336 280220
rect 171784 280168 171836 280220
rect 197452 280168 197504 280220
rect 199384 280168 199436 280220
rect 223948 280168 224000 280220
rect 225604 280168 225656 280220
rect 251180 280168 251232 280220
rect 253204 280168 253256 280220
rect 278044 280168 278096 280220
rect 279424 280168 279476 280220
rect 305460 280168 305512 280220
rect 307024 280168 307076 280220
rect 331956 280168 332008 280220
rect 333244 280168 333296 280220
rect 359464 280168 359516 280220
rect 359740 280168 359792 280220
rect 386052 280168 386104 280220
rect 387064 280168 387116 280220
rect 412916 280168 412968 280220
rect 414664 280168 414716 280220
rect 440240 280168 440292 280220
rect 442264 280168 442316 280220
rect 467012 280168 467064 280220
rect 468484 280168 468536 280220
rect 494060 280168 494112 280220
rect 496084 280168 496136 280220
rect 520924 280168 520976 280220
rect 522396 280168 522448 280220
rect 548064 280168 548116 280220
rect 37924 279420 37976 279472
rect 526444 279420 526496 279472
rect 285772 278264 285824 278316
rect 286140 278264 286192 278316
rect 339592 278264 339644 278316
rect 340144 278264 340196 278316
rect 68928 277516 68980 277568
rect 118700 277516 118752 277568
rect 311808 277516 311860 277568
rect 361580 277516 361632 277568
rect 35624 277448 35676 277500
rect 36636 277448 36688 277500
rect 41328 277448 41380 277500
rect 91100 277448 91152 277500
rect 122748 277448 122800 277500
rect 172520 277448 172572 277500
rect 176568 277448 176620 277500
rect 226340 277448 226392 277500
rect 230388 277448 230440 277500
rect 280160 277448 280212 277500
rect 284208 277448 284260 277500
rect 335360 277448 335412 277500
rect 365628 277448 365680 277500
rect 415400 277448 415452 277500
rect 419448 277448 419500 277500
rect 469220 277448 469272 277500
rect 473268 277448 473320 277500
rect 523040 277448 523092 277500
rect 13728 277380 13780 277432
rect 64880 277380 64932 277432
rect 95148 277380 95200 277432
rect 146300 277380 146352 277432
rect 148968 277380 149020 277432
rect 200120 277380 200172 277432
rect 202788 277380 202840 277432
rect 253940 277380 253992 277432
rect 256608 277380 256660 277432
rect 307760 277380 307812 277432
rect 338028 277380 338080 277432
rect 389180 277380 389232 277432
rect 391848 277380 391900 277432
rect 443000 277380 443052 277432
rect 445668 277380 445720 277432
rect 496820 277380 496872 277432
rect 500868 277380 500920 277432
rect 550640 277380 550692 277432
rect 170220 259632 170272 259684
rect 170496 259632 170548 259684
rect 446404 259428 446456 259480
rect 447692 259428 447744 259480
rect 35624 259360 35676 259412
rect 36820 259360 36872 259412
rect 278688 259360 278740 259412
rect 279516 259360 279568 259412
rect 332600 259360 332652 259412
rect 336004 259360 336056 259412
rect 467656 259360 467708 259412
rect 468576 259360 468628 259412
rect 26056 256640 26108 256692
rect 36728 256640 36780 256692
rect 62764 256640 62816 256692
rect 69756 256640 69808 256692
rect 96620 256640 96672 256692
rect 15200 256572 15252 256624
rect 42800 256572 42852 256624
rect 53104 256572 53156 256624
rect 64144 256572 64196 256624
rect 69112 256572 69164 256624
rect 96712 256572 96764 256624
rect 200764 256640 200816 256692
rect 204628 256640 204680 256692
rect 251824 256640 251876 256692
rect 258724 256640 258776 256692
rect 494704 256640 494756 256692
rect 501604 256640 501656 256692
rect 123668 256572 123720 256624
rect 149704 256572 149756 256624
rect 547972 256572 548024 256624
rect 79968 256504 80020 256556
rect 90456 256504 90508 256556
rect 106556 256504 106608 256556
rect 116584 256504 116636 256556
rect 133788 256504 133840 256556
rect 144276 256504 144328 256556
rect 150532 256504 150584 256556
rect 178132 256504 178184 256556
rect 187976 256504 188028 256556
rect 199384 256504 199436 256556
rect 204352 256504 204404 256556
rect 231952 256504 232004 256556
rect 242072 256504 242124 256556
rect 253204 256504 253256 256556
rect 258172 256504 258224 256556
rect 122932 256436 122984 256488
rect 150716 256436 150768 256488
rect 160560 256436 160612 256488
rect 171784 256436 171836 256488
rect 215024 256436 215076 256488
rect 225604 256436 225656 256488
rect 268936 256436 268988 256488
rect 279424 256436 279476 256488
rect 285772 256504 285824 256556
rect 312636 256504 312688 256556
rect 286140 256436 286192 256488
rect 295984 256436 296036 256488
rect 307024 256436 307076 256488
rect 311992 256436 312044 256488
rect 340144 256504 340196 256556
rect 322848 256436 322900 256488
rect 333244 256436 333296 256488
rect 339592 256436 339644 256488
rect 350080 256436 350132 256488
rect 359556 256436 359608 256488
rect 365812 256504 365864 256556
rect 393596 256504 393648 256556
rect 366732 256436 366784 256488
rect 376576 256436 376628 256488
rect 387064 256436 387116 256488
rect 393412 256436 393464 256488
rect 420920 256504 420972 256556
rect 431040 256504 431092 256556
rect 442264 256504 442316 256556
rect 447232 256504 447284 256556
rect 474740 256504 474792 256556
rect 484952 256504 485004 256556
rect 496084 256504 496136 256556
rect 501052 256504 501104 256556
rect 528652 256504 528704 256556
rect 403992 256436 404044 256488
rect 414664 256436 414716 256488
rect 458088 256436 458140 256488
rect 468484 256436 468536 256488
rect 511816 256436 511868 256488
rect 522396 256436 522448 256488
rect 36544 256368 36596 256420
rect 538404 256368 538456 256420
rect 16304 254532 16356 254584
rect 529020 254532 529072 254584
rect 25688 254192 25740 254244
rect 148324 254192 148376 254244
rect 36820 254124 36872 254176
rect 52644 254124 52696 254176
rect 232044 254124 232096 254176
rect 251824 254124 251876 254176
rect 475016 254124 475068 254176
rect 494704 254124 494756 254176
rect 62488 254056 62540 254108
rect 79692 254056 79744 254108
rect 90364 254056 90416 254108
rect 106648 254056 106700 254108
rect 116492 254056 116544 254108
rect 133696 254056 133748 254108
rect 170496 254056 170548 254108
rect 187700 254056 187752 254108
rect 197452 254056 197504 254108
rect 214656 254056 214708 254108
rect 224500 254056 224552 254108
rect 241704 254056 241756 254108
rect 413468 254056 413520 254108
rect 430672 254056 430724 254108
rect 440516 254056 440568 254108
rect 457628 254056 457680 254108
rect 468576 254056 468628 254108
rect 484676 254056 484728 254108
rect 36728 253988 36780 254040
rect 62304 253988 62356 254040
rect 64144 253988 64196 254040
rect 89352 253988 89404 254040
rect 90456 253988 90508 254040
rect 116308 253988 116360 254040
rect 116584 253988 116636 254040
rect 143356 253988 143408 254040
rect 144276 253988 144328 254040
rect 170312 253988 170364 254040
rect 178040 253988 178092 254040
rect 200764 253988 200816 254040
rect 251456 253988 251508 254040
rect 268660 253988 268712 254040
rect 279424 253988 279476 254040
rect 295708 253988 295760 254040
rect 305460 253988 305512 254040
rect 322664 253988 322716 254040
rect 334624 253988 334676 254040
rect 349712 253988 349764 254040
rect 359464 253988 359516 254040
rect 376668 253988 376720 254040
rect 386512 253988 386564 254040
rect 403624 253988 403676 254040
rect 421012 253988 421064 254040
rect 443644 253988 443696 254040
rect 494520 253988 494572 254040
rect 511632 253988 511684 254040
rect 522396 253988 522448 254040
rect 538680 253988 538732 254040
rect 43076 253920 43128 253972
rect 62764 253920 62816 253972
rect 144184 253920 144236 253972
rect 160652 253920 160704 253972
rect 171784 253920 171836 253972
rect 197360 253920 197412 253972
rect 199384 253920 199436 253972
rect 224316 253920 224368 253972
rect 225604 253920 225656 253972
rect 251364 253920 251416 253972
rect 253204 253920 253256 253972
rect 278320 253920 278372 253972
rect 279516 253920 279568 253972
rect 305368 253920 305420 253972
rect 307024 253920 307076 253972
rect 332324 253920 332376 253972
rect 333244 253920 333296 253972
rect 359372 253920 359424 253972
rect 359556 253920 359608 253972
rect 386328 253920 386380 253972
rect 387064 253920 387116 253972
rect 413284 253920 413336 253972
rect 414664 253920 414716 253972
rect 440332 253920 440384 253972
rect 442264 253920 442316 253972
rect 467288 253920 467340 253972
rect 468484 253920 468536 253972
rect 494336 253920 494388 253972
rect 496084 253920 496136 253972
rect 521292 253920 521344 253972
rect 522304 253920 522356 253972
rect 548340 253920 548392 253972
rect 37924 251812 37976 251864
rect 526444 251812 526496 251864
rect 68928 251268 68980 251320
rect 118700 251268 118752 251320
rect 122748 251268 122800 251320
rect 172520 251268 172572 251320
rect 230388 251268 230440 251320
rect 280160 251268 280212 251320
rect 311808 251268 311860 251320
rect 361580 251268 361632 251320
rect 500868 251268 500920 251320
rect 550640 251268 550692 251320
rect 41328 251200 41380 251252
rect 91100 251200 91152 251252
rect 148968 251200 149020 251252
rect 200120 251200 200172 251252
rect 202788 251200 202840 251252
rect 253940 251200 253992 251252
rect 284208 251200 284260 251252
rect 335360 251200 335412 251252
rect 365628 251200 365680 251252
rect 415400 251200 415452 251252
rect 419448 251200 419500 251252
rect 469220 251200 469272 251252
rect 473268 251200 473320 251252
rect 523040 251200 523092 251252
rect 521752 235356 521804 235408
rect 522396 235356 522448 235408
rect 13728 233180 13780 233232
rect 64880 233180 64932 233232
rect 95148 233180 95200 233232
rect 146300 233180 146352 233232
rect 176568 233180 176620 233232
rect 226340 233180 226392 233232
rect 256608 233180 256660 233232
rect 307760 233180 307812 233232
rect 332508 233180 332560 233232
rect 334624 233180 334676 233232
rect 338028 233180 338080 233232
rect 389180 233180 389232 233232
rect 391848 233180 391900 233232
rect 443000 233180 443052 233232
rect 445668 233180 445720 233232
rect 496820 233180 496872 233232
rect 467656 233112 467708 233164
rect 468576 233112 468628 233164
rect 35624 232704 35676 232756
rect 36820 232704 36872 232756
rect 257988 231820 258040 231872
rect 258724 231820 258776 231872
rect 494704 231820 494756 231872
rect 501604 231820 501656 231872
rect 26056 230392 26108 230444
rect 36728 230392 36780 230444
rect 62764 230392 62816 230444
rect 69756 230392 69808 230444
rect 96712 230392 96764 230444
rect 15200 230324 15252 230376
rect 42800 230324 42852 230376
rect 53104 230324 53156 230376
rect 64144 230324 64196 230376
rect 69112 230324 69164 230376
rect 96804 230324 96856 230376
rect 146944 230392 146996 230444
rect 123668 230324 123720 230376
rect 133788 230324 133840 230376
rect 144276 230324 144328 230376
rect 79968 230256 80020 230308
rect 90456 230256 90508 230308
rect 106556 230256 106608 230308
rect 116584 230256 116636 230308
rect 122932 230256 122984 230308
rect 150716 230324 150768 230376
rect 200764 230392 200816 230444
rect 204628 230392 204680 230444
rect 251824 230392 251876 230444
rect 257988 230392 258040 230444
rect 443644 230392 443696 230444
rect 447692 230392 447744 230444
rect 547972 230324 548024 230376
rect 150532 230256 150584 230308
rect 178132 230256 178184 230308
rect 187976 230256 188028 230308
rect 199384 230256 199436 230308
rect 204352 230256 204404 230308
rect 231860 230256 231912 230308
rect 242072 230256 242124 230308
rect 253204 230256 253256 230308
rect 258172 230256 258224 230308
rect 286140 230256 286192 230308
rect 160560 230188 160612 230240
rect 171784 230188 171836 230240
rect 215024 230188 215076 230240
rect 225604 230188 225656 230240
rect 268936 230188 268988 230240
rect 279516 230188 279568 230240
rect 285772 230188 285824 230240
rect 312636 230256 312688 230308
rect 295984 230188 296036 230240
rect 307024 230188 307076 230240
rect 311992 230188 312044 230240
rect 340144 230256 340196 230308
rect 322848 230188 322900 230240
rect 333244 230188 333296 230240
rect 339592 230188 339644 230240
rect 366732 230256 366784 230308
rect 350080 230188 350132 230240
rect 359556 230188 359608 230240
rect 365812 230188 365864 230240
rect 393596 230256 393648 230308
rect 376576 230188 376628 230240
rect 387064 230188 387116 230240
rect 393412 230188 393464 230240
rect 420920 230256 420972 230308
rect 431040 230256 431092 230308
rect 442264 230256 442316 230308
rect 447232 230256 447284 230308
rect 474740 230256 474792 230308
rect 484952 230256 485004 230308
rect 496084 230256 496136 230308
rect 501052 230256 501104 230308
rect 528652 230256 528704 230308
rect 403992 230188 404044 230240
rect 414664 230188 414716 230240
rect 458088 230188 458140 230240
rect 468484 230188 468536 230240
rect 511908 230188 511960 230240
rect 522304 230188 522356 230240
rect 36636 230120 36688 230172
rect 538404 230120 538456 230172
rect 15292 226992 15344 227044
rect 528744 226992 528796 227044
rect 25964 226584 26016 226636
rect 146944 226584 146996 226636
rect 36820 226516 36872 226568
rect 52460 226516 52512 226568
rect 62488 226516 62540 226568
rect 79324 226516 79376 226568
rect 259368 226516 259420 226568
rect 279608 226516 279660 226568
rect 448336 226516 448388 226568
rect 468668 226516 468720 226568
rect 43352 226448 43404 226500
rect 62764 226448 62816 226500
rect 90364 226448 90416 226500
rect 106372 226448 106424 226500
rect 116492 226448 116544 226500
rect 133420 226448 133472 226500
rect 170496 226448 170548 226500
rect 187792 226448 187844 226500
rect 197544 226448 197596 226500
rect 214380 226448 214432 226500
rect 224500 226448 224552 226500
rect 241520 226448 241572 226500
rect 251456 226448 251508 226500
rect 268292 226448 268344 226500
rect 413468 226448 413520 226500
rect 430580 226448 430632 226500
rect 440516 226448 440568 226500
rect 457260 226448 457312 226500
rect 36728 226380 36780 226432
rect 62120 226380 62172 226432
rect 64144 226380 64196 226432
rect 89076 226380 89128 226432
rect 90456 226380 90508 226432
rect 115940 226380 115992 226432
rect 116584 226380 116636 226432
rect 142988 226380 143040 226432
rect 144276 226380 144328 226432
rect 170036 226380 170088 226432
rect 178408 226380 178460 226432
rect 200764 226380 200816 226432
rect 232320 226380 232372 226432
rect 251824 226380 251876 226432
rect 279424 226380 279476 226432
rect 295800 226380 295852 226432
rect 305644 226380 305696 226432
rect 322388 226380 322440 226432
rect 336004 226380 336056 226432
rect 349804 226380 349856 226432
rect 359556 226380 359608 226432
rect 376300 226380 376352 226432
rect 386512 226380 386564 226432
rect 403348 226380 403400 226432
rect 421288 226380 421340 226432
rect 445024 226380 445076 226432
rect 468576 226380 468628 226432
rect 484400 226380 484452 226432
rect 494520 226380 494572 226432
rect 511356 226380 511408 226432
rect 522396 226380 522448 226432
rect 538404 226380 538456 226432
rect 70308 226312 70360 226364
rect 90548 226312 90600 226364
rect 144184 226312 144236 226364
rect 160284 226312 160336 226364
rect 171784 226312 171836 226364
rect 197452 226312 197504 226364
rect 199384 226312 199436 226364
rect 223948 226312 224000 226364
rect 225604 226312 225656 226364
rect 251180 226312 251232 226364
rect 253204 226312 253256 226364
rect 278044 226312 278096 226364
rect 279516 226312 279568 226364
rect 305552 226312 305604 226364
rect 307024 226312 307076 226364
rect 331956 226312 332008 226364
rect 333244 226312 333296 226364
rect 359464 226312 359516 226364
rect 359740 226312 359792 226364
rect 386052 226312 386104 226364
rect 387064 226312 387116 226364
rect 412916 226312 412968 226364
rect 414664 226312 414716 226364
rect 440240 226312 440292 226364
rect 442264 226312 442316 226364
rect 467012 226312 467064 226364
rect 468484 226312 468536 226364
rect 494060 226312 494112 226364
rect 496084 226312 496136 226364
rect 520924 226312 520976 226364
rect 522304 226312 522356 226364
rect 548064 226312 548116 226364
rect 37924 225564 37976 225616
rect 526444 225564 526496 225616
rect 285772 224272 285824 224324
rect 286140 224272 286192 224324
rect 339592 224272 339644 224324
rect 340144 224272 340196 224324
rect 35624 223592 35676 223644
rect 36636 223592 36688 223644
rect 90548 206252 90600 206304
rect 96804 206252 96856 206304
rect 468668 206252 468720 206304
rect 474740 206252 474792 206304
rect 474832 205708 474884 205760
rect 279608 205640 279660 205692
rect 286140 205640 286192 205692
rect 445024 205640 445076 205692
rect 447692 205640 447744 205692
rect 475200 205640 475252 205692
rect 521752 205640 521804 205692
rect 522396 205640 522448 205692
rect 13728 205572 13780 205624
rect 64880 205572 64932 205624
rect 95148 205572 95200 205624
rect 146300 205572 146352 205624
rect 148968 205572 149020 205624
rect 200120 205572 200172 205624
rect 202788 205572 202840 205624
rect 253940 205572 253992 205624
rect 256608 205572 256660 205624
rect 307760 205572 307812 205624
rect 338028 205572 338080 205624
rect 389180 205572 389232 205624
rect 391848 205572 391900 205624
rect 443000 205572 443052 205624
rect 445668 205572 445720 205624
rect 496820 205572 496872 205624
rect 500868 205572 500920 205624
rect 550640 205572 550692 205624
rect 35624 205504 35676 205556
rect 36820 205504 36872 205556
rect 41328 205504 41380 205556
rect 91100 205504 91152 205556
rect 122748 205504 122800 205556
rect 172520 205504 172572 205556
rect 176568 205504 176620 205556
rect 226340 205504 226392 205556
rect 230388 205504 230440 205556
rect 280160 205504 280212 205556
rect 284208 205504 284260 205556
rect 335360 205504 335412 205556
rect 365628 205504 365680 205556
rect 415400 205504 415452 205556
rect 419448 205504 419500 205556
rect 469220 205504 469272 205556
rect 473268 205504 473320 205556
rect 523040 205504 523092 205556
rect 68928 205436 68980 205488
rect 118700 205436 118752 205488
rect 200764 205436 200816 205488
rect 204628 205436 204680 205488
rect 311808 205436 311860 205488
rect 361580 205436 361632 205488
rect 467656 205436 467708 205488
rect 468576 205436 468628 205488
rect 53104 202784 53156 202836
rect 64144 202784 64196 202836
rect 251824 202784 251876 202836
rect 259000 202784 259052 202836
rect 332324 202784 332376 202836
rect 336004 202784 336056 202836
rect 15200 202716 15252 202768
rect 42984 202716 43036 202768
rect 62764 202716 62816 202768
rect 70032 202716 70084 202768
rect 79692 202716 79744 202768
rect 90456 202716 90508 202768
rect 96712 202716 96764 202768
rect 124036 202716 124088 202768
rect 148324 202716 148376 202768
rect 548340 202716 548392 202768
rect 25688 202648 25740 202700
rect 36728 202648 36780 202700
rect 106648 202648 106700 202700
rect 116584 202648 116636 202700
rect 133696 202648 133748 202700
rect 144276 202648 144328 202700
rect 150532 202648 150584 202700
rect 178040 202648 178092 202700
rect 187700 202648 187752 202700
rect 199384 202648 199436 202700
rect 204352 202648 204404 202700
rect 232044 202648 232096 202700
rect 241704 202648 241756 202700
rect 253204 202648 253256 202700
rect 268660 202648 268712 202700
rect 279516 202648 279568 202700
rect 285772 202648 285824 202700
rect 313004 202648 313056 202700
rect 122932 202580 122984 202632
rect 150992 202580 151044 202632
rect 160652 202580 160704 202632
rect 171784 202580 171836 202632
rect 214656 202580 214708 202632
rect 225604 202580 225656 202632
rect 295708 202580 295760 202632
rect 307024 202580 307076 202632
rect 311992 202580 312044 202632
rect 340052 202648 340104 202700
rect 322664 202580 322716 202632
rect 333244 202580 333296 202632
rect 339592 202580 339644 202632
rect 367008 202648 367060 202700
rect 349712 202580 349764 202632
rect 359556 202580 359608 202632
rect 365812 202580 365864 202632
rect 393596 202648 393648 202700
rect 376668 202580 376720 202632
rect 387064 202580 387116 202632
rect 393412 202580 393464 202632
rect 421012 202648 421064 202700
rect 430672 202648 430724 202700
rect 442264 202648 442316 202700
rect 457720 202648 457772 202700
rect 468484 202648 468536 202700
rect 475200 202648 475252 202700
rect 501972 202648 502024 202700
rect 403716 202580 403768 202632
rect 414664 202580 414716 202632
rect 484676 202580 484728 202632
rect 496084 202580 496136 202632
rect 501052 202580 501104 202632
rect 529020 202648 529072 202700
rect 511724 202580 511776 202632
rect 522304 202580 522356 202632
rect 36544 202512 36596 202564
rect 538680 202512 538732 202564
rect 16028 200744 16080 200796
rect 529020 200744 529072 200796
rect 25688 200404 25740 200456
rect 149704 200404 149756 200456
rect 36728 200336 36780 200388
rect 52644 200336 52696 200388
rect 232044 200336 232096 200388
rect 251824 200336 251876 200388
rect 43076 200268 43128 200320
rect 62764 200268 62816 200320
rect 90364 200268 90416 200320
rect 106648 200268 106700 200320
rect 116492 200268 116544 200320
rect 133696 200268 133748 200320
rect 144184 200268 144236 200320
rect 160652 200268 160704 200320
rect 170496 200268 170548 200320
rect 187700 200268 187752 200320
rect 197452 200268 197504 200320
rect 214656 200268 214708 200320
rect 224500 200268 224552 200320
rect 241704 200268 241756 200320
rect 413468 200268 413520 200320
rect 430672 200268 430724 200320
rect 440516 200268 440568 200320
rect 457628 200268 457680 200320
rect 468576 200268 468628 200320
rect 484676 200268 484728 200320
rect 494520 200268 494572 200320
rect 511632 200268 511684 200320
rect 36820 200200 36872 200252
rect 62304 200200 62356 200252
rect 64144 200200 64196 200252
rect 89352 200200 89404 200252
rect 90456 200200 90508 200252
rect 116308 200200 116360 200252
rect 116584 200200 116636 200252
rect 143356 200200 143408 200252
rect 144276 200200 144328 200252
rect 170312 200200 170364 200252
rect 178040 200200 178092 200252
rect 200764 200200 200816 200252
rect 251456 200200 251508 200252
rect 268660 200200 268712 200252
rect 279424 200200 279476 200252
rect 295708 200200 295760 200252
rect 305460 200200 305512 200252
rect 322664 200200 322716 200252
rect 336004 200200 336056 200252
rect 349712 200200 349764 200252
rect 359464 200200 359516 200252
rect 376668 200200 376720 200252
rect 386512 200200 386564 200252
rect 403624 200200 403676 200252
rect 421012 200200 421064 200252
rect 446404 200200 446456 200252
rect 475016 200200 475068 200252
rect 494704 200200 494756 200252
rect 522396 200200 522448 200252
rect 538680 200200 538732 200252
rect 62488 200132 62540 200184
rect 79692 200132 79744 200184
rect 171784 200132 171836 200184
rect 197360 200132 197412 200184
rect 199384 200132 199436 200184
rect 224316 200132 224368 200184
rect 225604 200132 225656 200184
rect 251364 200132 251416 200184
rect 253204 200132 253256 200184
rect 278320 200132 278372 200184
rect 279516 200132 279568 200184
rect 305368 200132 305420 200184
rect 307024 200132 307076 200184
rect 332324 200132 332376 200184
rect 333244 200132 333296 200184
rect 359372 200132 359424 200184
rect 359556 200132 359608 200184
rect 386328 200132 386380 200184
rect 387064 200132 387116 200184
rect 413284 200132 413336 200184
rect 414664 200132 414716 200184
rect 440332 200132 440384 200184
rect 442264 200132 442316 200184
rect 467288 200132 467340 200184
rect 468484 200132 468536 200184
rect 494336 200132 494388 200184
rect 496084 200132 496136 200184
rect 521292 200132 521344 200184
rect 522304 200132 522356 200184
rect 548340 200132 548392 200184
rect 37924 197956 37976 198008
rect 526444 197956 526496 198008
rect 445668 179392 445720 179444
rect 13728 179324 13780 179376
rect 64880 179324 64932 179376
rect 95148 179324 95200 179376
rect 146300 179324 146352 179376
rect 148968 179324 149020 179376
rect 200120 179324 200172 179376
rect 202788 179324 202840 179376
rect 253940 179324 253992 179376
rect 256608 179324 256660 179376
rect 307760 179324 307812 179376
rect 338028 179324 338080 179376
rect 389180 179324 389232 179376
rect 391848 179324 391900 179376
rect 443000 179324 443052 179376
rect 446404 179324 446456 179376
rect 447692 179324 447744 179376
rect 521752 179392 521804 179444
rect 522396 179392 522448 179444
rect 496820 179324 496872 179376
rect 500868 179324 500920 179376
rect 550640 179324 550692 179376
rect 35624 179256 35676 179308
rect 36728 179256 36780 179308
rect 41328 179256 41380 179308
rect 91100 179256 91152 179308
rect 122748 179256 122800 179308
rect 172520 179256 172572 179308
rect 176568 179256 176620 179308
rect 226340 179256 226392 179308
rect 230388 179256 230440 179308
rect 280160 179256 280212 179308
rect 284208 179256 284260 179308
rect 335360 179256 335412 179308
rect 365628 179256 365680 179308
rect 415400 179256 415452 179308
rect 419448 179256 419500 179308
rect 68928 179188 68980 179240
rect 118700 179188 118752 179240
rect 311808 179188 311860 179240
rect 361580 179188 361632 179240
rect 469220 179256 469272 179308
rect 473268 179256 473320 179308
rect 523040 179256 523092 179308
rect 467656 179188 467708 179240
rect 468576 179188 468628 179240
rect 62764 176604 62816 176656
rect 69756 176604 69808 176656
rect 96712 176604 96764 176656
rect 15200 176536 15252 176588
rect 42800 176536 42852 176588
rect 53104 176536 53156 176588
rect 64144 176536 64196 176588
rect 69112 176536 69164 176588
rect 96804 176536 96856 176588
rect 146944 176604 146996 176656
rect 123668 176536 123720 176588
rect 133788 176536 133840 176588
rect 144276 176536 144328 176588
rect 150532 176536 150584 176588
rect 200764 176604 200816 176656
rect 204628 176604 204680 176656
rect 251824 176604 251876 176656
rect 258724 176604 258776 176656
rect 332508 176604 332560 176656
rect 336004 176604 336056 176656
rect 494704 176604 494756 176656
rect 501604 176604 501656 176656
rect 26056 176468 26108 176520
rect 36820 176468 36872 176520
rect 79968 176468 80020 176520
rect 90456 176468 90508 176520
rect 106556 176468 106608 176520
rect 116584 176468 116636 176520
rect 122932 176468 122984 176520
rect 150716 176468 150768 176520
rect 547972 176536 548024 176588
rect 178132 176468 178184 176520
rect 187976 176468 188028 176520
rect 199384 176468 199436 176520
rect 204352 176468 204404 176520
rect 231860 176468 231912 176520
rect 242072 176468 242124 176520
rect 253204 176468 253256 176520
rect 258172 176468 258224 176520
rect 286140 176468 286192 176520
rect 160560 176400 160612 176452
rect 171784 176400 171836 176452
rect 215024 176400 215076 176452
rect 225604 176400 225656 176452
rect 268936 176400 268988 176452
rect 279516 176400 279568 176452
rect 285772 176400 285824 176452
rect 312636 176468 312688 176520
rect 295984 176400 296036 176452
rect 307024 176400 307076 176452
rect 311992 176400 312044 176452
rect 340144 176468 340196 176520
rect 322848 176400 322900 176452
rect 333244 176400 333296 176452
rect 339592 176400 339644 176452
rect 366732 176468 366784 176520
rect 350080 176400 350132 176452
rect 359556 176400 359608 176452
rect 365812 176400 365864 176452
rect 393596 176468 393648 176520
rect 376576 176400 376628 176452
rect 387064 176400 387116 176452
rect 393412 176400 393464 176452
rect 420920 176468 420972 176520
rect 431040 176468 431092 176520
rect 442264 176468 442316 176520
rect 447232 176468 447284 176520
rect 474740 176468 474792 176520
rect 484952 176468 485004 176520
rect 496084 176468 496136 176520
rect 501052 176468 501104 176520
rect 528652 176468 528704 176520
rect 403992 176400 404044 176452
rect 414664 176400 414716 176452
rect 458088 176400 458140 176452
rect 468484 176400 468536 176452
rect 511908 176400 511960 176452
rect 522304 176400 522356 176452
rect 36636 176332 36688 176384
rect 538404 176332 538456 176384
rect 16304 173136 16356 173188
rect 528652 173136 528704 173188
rect 26056 172796 26108 172848
rect 146944 172796 146996 172848
rect 36728 172728 36780 172780
rect 52460 172728 52512 172780
rect 232320 172728 232372 172780
rect 251824 172728 251876 172780
rect 475384 172728 475436 172780
rect 494704 172728 494756 172780
rect 62488 172660 62540 172712
rect 79324 172660 79376 172712
rect 90456 172660 90508 172712
rect 106464 172660 106516 172712
rect 116492 172660 116544 172712
rect 133420 172660 133472 172712
rect 170496 172660 170548 172712
rect 187792 172660 187844 172712
rect 197544 172660 197596 172712
rect 214380 172660 214432 172712
rect 224500 172660 224552 172712
rect 241612 172660 241664 172712
rect 413468 172660 413520 172712
rect 430580 172660 430632 172712
rect 440516 172660 440568 172712
rect 457260 172660 457312 172712
rect 468484 172660 468536 172712
rect 484400 172660 484452 172712
rect 36820 172592 36872 172644
rect 62120 172592 62172 172644
rect 64144 172592 64196 172644
rect 89076 172592 89128 172644
rect 90364 172592 90416 172644
rect 116124 172592 116176 172644
rect 116584 172592 116636 172644
rect 142988 172592 143040 172644
rect 144184 172592 144236 172644
rect 170036 172592 170088 172644
rect 178408 172592 178460 172644
rect 200764 172592 200816 172644
rect 251456 172592 251508 172644
rect 268292 172592 268344 172644
rect 279424 172592 279476 172644
rect 295800 172592 295852 172644
rect 305552 172592 305604 172644
rect 322388 172592 322440 172644
rect 334624 172592 334676 172644
rect 349804 172592 349856 172644
rect 359648 172592 359700 172644
rect 376300 172592 376352 172644
rect 386512 172592 386564 172644
rect 403348 172592 403400 172644
rect 421288 172592 421340 172644
rect 443644 172592 443696 172644
rect 494520 172592 494572 172644
rect 511356 172592 511408 172644
rect 522304 172592 522356 172644
rect 538404 172592 538456 172644
rect 43352 172524 43404 172576
rect 62764 172524 62816 172576
rect 144276 172524 144328 172576
rect 160284 172524 160336 172576
rect 171784 172524 171836 172576
rect 197452 172524 197504 172576
rect 199384 172524 199436 172576
rect 223948 172524 224000 172576
rect 225604 172524 225656 172576
rect 251272 172524 251324 172576
rect 253204 172524 253256 172576
rect 278044 172524 278096 172576
rect 279516 172524 279568 172576
rect 305460 172524 305512 172576
rect 307024 172524 307076 172576
rect 331956 172524 332008 172576
rect 333244 172524 333296 172576
rect 359464 172524 359516 172576
rect 359556 172524 359608 172576
rect 386052 172524 386104 172576
rect 387064 172524 387116 172576
rect 412916 172524 412968 172576
rect 414664 172524 414716 172576
rect 440240 172524 440292 172576
rect 442264 172524 442316 172576
rect 467012 172524 467064 172576
rect 468576 172524 468628 172576
rect 494060 172524 494112 172576
rect 496084 172524 496136 172576
rect 520924 172524 520976 172576
rect 522396 172524 522448 172576
rect 547972 172524 548024 172576
rect 37924 170348 37976 170400
rect 526444 170348 526496 170400
rect 285772 170280 285824 170332
rect 286140 170280 286192 170332
rect 339592 170280 339644 170332
rect 340144 170280 340196 170332
rect 35624 169736 35676 169788
rect 36636 169736 36688 169788
rect 359556 166336 359608 166388
rect 359556 166132 359608 166184
rect 89720 156612 89772 156664
rect 90456 156612 90508 156664
rect 143632 154300 143684 154352
rect 144276 154300 144328 154352
rect 13728 151716 13780 151768
rect 64880 151716 64932 151768
rect 95148 151716 95200 151768
rect 146300 151716 146352 151768
rect 148968 151716 149020 151768
rect 200120 151716 200172 151768
rect 202788 151716 202840 151768
rect 253940 151716 253992 151768
rect 256608 151716 256660 151768
rect 307760 151716 307812 151768
rect 332508 151716 332560 151768
rect 334624 151716 334676 151768
rect 338028 151716 338080 151768
rect 389180 151716 389232 151768
rect 391848 151716 391900 151768
rect 443000 151716 443052 151768
rect 445668 151716 445720 151768
rect 496820 151716 496872 151768
rect 500868 151716 500920 151768
rect 550640 151716 550692 151768
rect 35624 151648 35676 151700
rect 36728 151648 36780 151700
rect 41328 151648 41380 151700
rect 91100 151648 91152 151700
rect 122748 151648 122800 151700
rect 172520 151648 172572 151700
rect 176568 151648 176620 151700
rect 226340 151648 226392 151700
rect 230388 151648 230440 151700
rect 280160 151648 280212 151700
rect 284208 151648 284260 151700
rect 335360 151648 335412 151700
rect 365628 151648 365680 151700
rect 415400 151648 415452 151700
rect 419448 151648 419500 151700
rect 469220 151648 469272 151700
rect 473268 151648 473320 151700
rect 523040 151648 523092 151700
rect 68928 151580 68980 151632
rect 118700 151580 118752 151632
rect 200764 151580 200816 151632
rect 204628 151580 204680 151632
rect 311808 151580 311860 151632
rect 361580 151580 361632 151632
rect 443644 151580 443696 151632
rect 447692 151580 447744 151632
rect 52736 148996 52788 149048
rect 64144 148996 64196 149048
rect 69112 148996 69164 149048
rect 15200 148928 15252 148980
rect 42984 148928 43036 148980
rect 62764 148928 62816 148980
rect 70032 148928 70084 148980
rect 96712 148996 96764 149048
rect 96988 148928 97040 148980
rect 251824 148996 251876 149048
rect 259000 148996 259052 149048
rect 494704 148996 494756 149048
rect 501972 148996 502024 149048
rect 124036 148928 124088 148980
rect 149704 148928 149756 148980
rect 548340 148928 548392 148980
rect 25688 148860 25740 148912
rect 36820 148860 36872 148912
rect 79692 148860 79744 148912
rect 90364 148860 90416 148912
rect 106648 148860 106700 148912
rect 116584 148860 116636 148912
rect 133696 148860 133748 148912
rect 144184 148860 144236 148912
rect 150532 148860 150584 148912
rect 178040 148860 178092 148912
rect 187700 148860 187752 148912
rect 199384 148860 199436 148912
rect 204352 148860 204404 148912
rect 232044 148860 232096 148912
rect 241704 148860 241756 148912
rect 253204 148860 253256 148912
rect 258172 148860 258224 148912
rect 286048 148860 286100 148912
rect 122932 148792 122984 148844
rect 150992 148792 151044 148844
rect 160652 148792 160704 148844
rect 171784 148792 171836 148844
rect 214656 148792 214708 148844
rect 225604 148792 225656 148844
rect 268660 148792 268712 148844
rect 279516 148792 279568 148844
rect 285772 148792 285824 148844
rect 313004 148860 313056 148912
rect 295708 148792 295760 148844
rect 307024 148792 307076 148844
rect 311992 148792 312044 148844
rect 340052 148860 340104 148912
rect 322664 148792 322716 148844
rect 333244 148792 333296 148844
rect 339592 148792 339644 148844
rect 367008 148860 367060 148912
rect 349712 148792 349764 148844
rect 359556 148792 359608 148844
rect 365812 148792 365864 148844
rect 393964 148860 394016 148912
rect 376668 148792 376720 148844
rect 387064 148792 387116 148844
rect 393412 148792 393464 148844
rect 421012 148860 421064 148912
rect 430672 148860 430724 148912
rect 442264 148860 442316 148912
rect 447232 148860 447284 148912
rect 475016 148860 475068 148912
rect 484676 148860 484728 148912
rect 496084 148860 496136 148912
rect 501052 148860 501104 148912
rect 529020 148860 529072 148912
rect 403716 148792 403768 148844
rect 414664 148792 414716 148844
rect 457720 148792 457772 148844
rect 468576 148792 468628 148844
rect 511724 148792 511776 148844
rect 522396 148792 522448 148844
rect 36544 148724 36596 148776
rect 538680 148724 538732 148776
rect 16028 146888 16080 146940
rect 529020 146888 529072 146940
rect 25688 146548 25740 146600
rect 149704 146548 149756 146600
rect 36728 146480 36780 146532
rect 52644 146480 52696 146532
rect 232044 146480 232096 146532
rect 251824 146480 251876 146532
rect 475016 146480 475068 146532
rect 494704 146480 494756 146532
rect 62488 146412 62540 146464
rect 79692 146412 79744 146464
rect 90456 146412 90508 146464
rect 106648 146412 106700 146464
rect 116492 146412 116544 146464
rect 133696 146412 133748 146464
rect 144184 146412 144236 146464
rect 160652 146412 160704 146464
rect 170496 146412 170548 146464
rect 187700 146412 187752 146464
rect 197452 146412 197504 146464
rect 214656 146412 214708 146464
rect 224500 146412 224552 146464
rect 241704 146412 241756 146464
rect 413468 146412 413520 146464
rect 430672 146412 430724 146464
rect 440516 146412 440568 146464
rect 457628 146412 457680 146464
rect 468484 146412 468536 146464
rect 484676 146412 484728 146464
rect 36820 146344 36872 146396
rect 62304 146344 62356 146396
rect 64144 146344 64196 146396
rect 89352 146344 89404 146396
rect 90364 146344 90416 146396
rect 116308 146344 116360 146396
rect 116584 146344 116636 146396
rect 143356 146344 143408 146396
rect 144276 146344 144328 146396
rect 170312 146344 170364 146396
rect 178040 146344 178092 146396
rect 200764 146344 200816 146396
rect 251456 146344 251508 146396
rect 268660 146344 268712 146396
rect 279516 146344 279568 146396
rect 295708 146344 295760 146396
rect 305460 146344 305512 146396
rect 322664 146344 322716 146396
rect 336004 146344 336056 146396
rect 349712 146344 349764 146396
rect 359464 146344 359516 146396
rect 376668 146344 376720 146396
rect 386512 146344 386564 146396
rect 403624 146344 403676 146396
rect 421012 146344 421064 146396
rect 445024 146344 445076 146396
rect 494520 146344 494572 146396
rect 511632 146344 511684 146396
rect 522396 146344 522448 146396
rect 538680 146344 538732 146396
rect 43076 146276 43128 146328
rect 62764 146276 62816 146328
rect 171784 146276 171836 146328
rect 197360 146276 197412 146328
rect 199384 146276 199436 146328
rect 224316 146276 224368 146328
rect 225604 146276 225656 146328
rect 251364 146276 251416 146328
rect 253204 146276 253256 146328
rect 278320 146276 278372 146328
rect 279424 146276 279476 146328
rect 305368 146276 305420 146328
rect 307024 146276 307076 146328
rect 332324 146276 332376 146328
rect 333244 146276 333296 146328
rect 359372 146276 359424 146328
rect 359556 146276 359608 146328
rect 386328 146276 386380 146328
rect 387064 146276 387116 146328
rect 413284 146276 413336 146328
rect 414664 146276 414716 146328
rect 440332 146276 440384 146328
rect 442264 146276 442316 146328
rect 467288 146276 467340 146328
rect 468576 146276 468628 146328
rect 494336 146276 494388 146328
rect 496084 146276 496136 146328
rect 521292 146276 521344 146328
rect 522304 146276 522356 146328
rect 548340 146276 548392 146328
rect 37924 144168 37976 144220
rect 526444 144168 526496 144220
rect 89720 128256 89772 128308
rect 90456 128256 90508 128308
rect 13728 125536 13780 125588
rect 64880 125536 64932 125588
rect 95148 125536 95200 125588
rect 146300 125536 146352 125588
rect 148968 125536 149020 125588
rect 200120 125536 200172 125588
rect 202788 125536 202840 125588
rect 253940 125536 253992 125588
rect 256608 125536 256660 125588
rect 307760 125536 307812 125588
rect 338028 125536 338080 125588
rect 389180 125536 389232 125588
rect 391848 125536 391900 125588
rect 443000 125536 443052 125588
rect 445668 125536 445720 125588
rect 496820 125536 496872 125588
rect 500868 125536 500920 125588
rect 550640 125536 550692 125588
rect 41328 125468 41380 125520
rect 91100 125468 91152 125520
rect 122748 125468 122800 125520
rect 172520 125468 172572 125520
rect 176568 125468 176620 125520
rect 226340 125468 226392 125520
rect 230388 125468 230440 125520
rect 68928 125400 68980 125452
rect 118700 125400 118752 125452
rect 278688 125468 278740 125520
rect 279516 125468 279568 125520
rect 284208 125468 284260 125520
rect 335360 125468 335412 125520
rect 365628 125468 365680 125520
rect 415400 125468 415452 125520
rect 419448 125468 419500 125520
rect 469220 125468 469272 125520
rect 473268 125468 473320 125520
rect 523040 125468 523092 125520
rect 280160 125400 280212 125452
rect 311808 125400 311860 125452
rect 361580 125400 361632 125452
rect 445024 125400 445076 125452
rect 447692 125400 447744 125452
rect 35624 124788 35676 124840
rect 36728 124788 36780 124840
rect 116216 124584 116268 124636
rect 116492 124584 116544 124636
rect 170220 124584 170272 124636
rect 170496 124584 170548 124636
rect 62764 122748 62816 122800
rect 69756 122748 69808 122800
rect 96620 122748 96672 122800
rect 15200 122680 15252 122732
rect 42800 122680 42852 122732
rect 53104 122680 53156 122732
rect 64144 122680 64196 122732
rect 69112 122680 69164 122732
rect 96712 122680 96764 122732
rect 200764 122748 200816 122800
rect 204628 122748 204680 122800
rect 251824 122748 251876 122800
rect 258724 122748 258776 122800
rect 332508 122748 332560 122800
rect 336004 122748 336056 122800
rect 494704 122748 494756 122800
rect 501604 122748 501656 122800
rect 521476 122748 521528 122800
rect 522396 122748 522448 122800
rect 123668 122680 123720 122732
rect 133788 122680 133840 122732
rect 144276 122680 144328 122732
rect 146944 122680 146996 122732
rect 547972 122680 548024 122732
rect 26056 122612 26108 122664
rect 36820 122612 36872 122664
rect 79968 122612 80020 122664
rect 90364 122612 90416 122664
rect 106556 122612 106608 122664
rect 116584 122612 116636 122664
rect 122932 122612 122984 122664
rect 150532 122612 150584 122664
rect 178132 122612 178184 122664
rect 187976 122612 188028 122664
rect 199384 122612 199436 122664
rect 204352 122612 204404 122664
rect 231952 122612 232004 122664
rect 242072 122612 242124 122664
rect 253204 122612 253256 122664
rect 258172 122612 258224 122664
rect 150716 122544 150768 122596
rect 160560 122544 160612 122596
rect 171784 122544 171836 122596
rect 215024 122544 215076 122596
rect 225604 122544 225656 122596
rect 268936 122544 268988 122596
rect 279424 122544 279476 122596
rect 285772 122612 285824 122664
rect 312636 122612 312688 122664
rect 286140 122544 286192 122596
rect 295984 122544 296036 122596
rect 307024 122544 307076 122596
rect 311992 122544 312044 122596
rect 322848 122544 322900 122596
rect 333244 122544 333296 122596
rect 339592 122612 339644 122664
rect 366732 122612 366784 122664
rect 340144 122544 340196 122596
rect 350080 122544 350132 122596
rect 359556 122544 359608 122596
rect 365812 122544 365864 122596
rect 393596 122612 393648 122664
rect 376576 122544 376628 122596
rect 387064 122544 387116 122596
rect 393412 122544 393464 122596
rect 420920 122612 420972 122664
rect 431040 122612 431092 122664
rect 442264 122612 442316 122664
rect 447232 122612 447284 122664
rect 474740 122612 474792 122664
rect 484952 122612 485004 122664
rect 496084 122612 496136 122664
rect 501052 122612 501104 122664
rect 528652 122612 528704 122664
rect 403992 122544 404044 122596
rect 414664 122544 414716 122596
rect 458088 122544 458140 122596
rect 468576 122544 468628 122596
rect 511816 122544 511868 122596
rect 522304 122544 522356 122596
rect 36636 122476 36688 122528
rect 538404 122476 538456 122528
rect 16304 119348 16356 119400
rect 528744 119348 528796 119400
rect 25964 118940 26016 118992
rect 146944 118940 146996 118992
rect 36820 118872 36872 118924
rect 52460 118872 52512 118924
rect 232320 118872 232372 118924
rect 251824 118872 251876 118924
rect 62488 118804 62540 118856
rect 79324 118804 79376 118856
rect 90456 118804 90508 118856
rect 106372 118804 106424 118856
rect 116492 118804 116544 118856
rect 133420 118804 133472 118856
rect 170496 118804 170548 118856
rect 187792 118804 187844 118856
rect 197544 118804 197596 118856
rect 214380 118804 214432 118856
rect 224500 118804 224552 118856
rect 241520 118804 241572 118856
rect 413468 118804 413520 118856
rect 430580 118804 430632 118856
rect 440516 118804 440568 118856
rect 457260 118804 457312 118856
rect 468576 118804 468628 118856
rect 484400 118804 484452 118856
rect 494520 118804 494572 118856
rect 511356 118804 511408 118856
rect 36636 118736 36688 118788
rect 62120 118736 62172 118788
rect 64144 118736 64196 118788
rect 89076 118736 89128 118788
rect 90364 118736 90416 118788
rect 115940 118736 115992 118788
rect 116584 118736 116636 118788
rect 142988 118736 143040 118788
rect 144184 118736 144236 118788
rect 170036 118736 170088 118788
rect 178408 118736 178460 118788
rect 200764 118736 200816 118788
rect 251456 118736 251508 118788
rect 268292 118736 268344 118788
rect 279424 118736 279476 118788
rect 295800 118736 295852 118788
rect 305644 118736 305696 118788
rect 322388 118736 322440 118788
rect 334624 118736 334676 118788
rect 349804 118736 349856 118788
rect 359556 118736 359608 118788
rect 376300 118736 376352 118788
rect 386512 118736 386564 118788
rect 403348 118736 403400 118788
rect 421288 118736 421340 118788
rect 443644 118736 443696 118788
rect 475384 118736 475436 118788
rect 494704 118736 494756 118788
rect 522396 118736 522448 118788
rect 538404 118736 538456 118788
rect 43352 118668 43404 118720
rect 62764 118668 62816 118720
rect 144276 118668 144328 118720
rect 160284 118668 160336 118720
rect 171784 118668 171836 118720
rect 197452 118668 197504 118720
rect 199384 118668 199436 118720
rect 223948 118668 224000 118720
rect 225604 118668 225656 118720
rect 251180 118668 251232 118720
rect 253204 118668 253256 118720
rect 278044 118668 278096 118720
rect 279516 118668 279568 118720
rect 305552 118668 305604 118720
rect 307024 118668 307076 118720
rect 331956 118668 332008 118720
rect 333244 118668 333296 118720
rect 359464 118668 359516 118720
rect 359740 118668 359792 118720
rect 386052 118668 386104 118720
rect 387064 118668 387116 118720
rect 412916 118668 412968 118720
rect 414664 118668 414716 118720
rect 440240 118668 440292 118720
rect 442264 118668 442316 118720
rect 467012 118668 467064 118720
rect 468484 118668 468536 118720
rect 494060 118668 494112 118720
rect 496084 118668 496136 118720
rect 520924 118668 520976 118720
rect 522304 118668 522356 118720
rect 548064 118668 548116 118720
rect 37924 116560 37976 116612
rect 526444 116560 526496 116612
rect 285772 116356 285824 116408
rect 286140 116356 286192 116408
rect 339592 116288 339644 116340
rect 340144 116288 340196 116340
rect 35624 116084 35676 116136
rect 36728 116084 36780 116136
rect 89720 100240 89772 100292
rect 90456 100240 90508 100292
rect 143632 100240 143684 100292
rect 144276 100240 144328 100292
rect 521752 100240 521804 100292
rect 522396 100240 522448 100292
rect 13728 97928 13780 97980
rect 64880 97928 64932 97980
rect 95148 97928 95200 97980
rect 146300 97928 146352 97980
rect 148968 97928 149020 97980
rect 200120 97928 200172 97980
rect 202788 97928 202840 97980
rect 253940 97928 253992 97980
rect 284208 97928 284260 97980
rect 335360 97928 335412 97980
rect 338028 97928 338080 97980
rect 389180 97928 389232 97980
rect 391848 97928 391900 97980
rect 443000 97928 443052 97980
rect 445668 97928 445720 97980
rect 496820 97928 496872 97980
rect 500868 97928 500920 97980
rect 550640 97928 550692 97980
rect 41328 97860 41380 97912
rect 91100 97860 91152 97912
rect 122748 97860 122800 97912
rect 172520 97860 172572 97912
rect 176568 97860 176620 97912
rect 226340 97860 226392 97912
rect 256608 97860 256660 97912
rect 307760 97860 307812 97912
rect 311808 97860 311860 97912
rect 361580 97860 361632 97912
rect 365628 97860 365680 97912
rect 415400 97860 415452 97912
rect 419448 97860 419500 97912
rect 469220 97860 469272 97912
rect 473268 97860 473320 97912
rect 523040 97860 523092 97912
rect 68928 97792 68980 97844
rect 118700 97792 118752 97844
rect 200764 97792 200816 97844
rect 204628 97792 204680 97844
rect 230388 97792 230440 97844
rect 280160 97792 280212 97844
rect 332508 97792 332560 97844
rect 334624 97792 334676 97844
rect 443644 97792 443696 97844
rect 447692 97792 447744 97844
rect 467656 97792 467708 97844
rect 468576 97792 468628 97844
rect 35624 97656 35676 97708
rect 36820 97656 36872 97708
rect 257988 96636 258040 96688
rect 258724 96636 258776 96688
rect 494704 96636 494756 96688
rect 501604 96636 501656 96688
rect 62764 95140 62816 95192
rect 70032 95140 70084 95192
rect 96712 95140 96764 95192
rect 15200 95072 15252 95124
rect 42984 95072 43036 95124
rect 52736 95072 52788 95124
rect 64144 95072 64196 95124
rect 69112 95072 69164 95124
rect 96988 95072 97040 95124
rect 251824 95140 251876 95192
rect 257988 95140 258040 95192
rect 124036 95072 124088 95124
rect 149704 95072 149756 95124
rect 548340 95072 548392 95124
rect 25688 95004 25740 95056
rect 36636 95004 36688 95056
rect 79692 95004 79744 95056
rect 90364 95004 90416 95056
rect 106648 95004 106700 95056
rect 116584 95004 116636 95056
rect 133696 95004 133748 95056
rect 144184 95004 144236 95056
rect 150532 95004 150584 95056
rect 178040 95004 178092 95056
rect 187700 95004 187752 95056
rect 199384 95004 199436 95056
rect 204352 95004 204404 95056
rect 232044 95004 232096 95056
rect 241704 95004 241756 95056
rect 253204 95004 253256 95056
rect 258172 95004 258224 95056
rect 286048 95004 286100 95056
rect 122932 94936 122984 94988
rect 150992 94936 151044 94988
rect 160652 94936 160704 94988
rect 171784 94936 171836 94988
rect 214656 94936 214708 94988
rect 225604 94936 225656 94988
rect 268660 94936 268712 94988
rect 279516 94936 279568 94988
rect 285772 94936 285824 94988
rect 313004 95004 313056 95056
rect 295708 94936 295760 94988
rect 307024 94936 307076 94988
rect 311992 94936 312044 94988
rect 340052 95004 340104 95056
rect 322664 94936 322716 94988
rect 333244 94936 333296 94988
rect 339592 94936 339644 94988
rect 367008 95004 367060 95056
rect 349712 94936 349764 94988
rect 359556 94936 359608 94988
rect 365812 94936 365864 94988
rect 393964 95004 394016 95056
rect 376668 94936 376720 94988
rect 387064 94936 387116 94988
rect 393412 94936 393464 94988
rect 421012 95004 421064 95056
rect 430672 95004 430724 95056
rect 442264 95004 442316 95056
rect 447232 95004 447284 95056
rect 475016 95004 475068 95056
rect 484676 95004 484728 95056
rect 496084 95004 496136 95056
rect 501052 95004 501104 95056
rect 529020 95004 529072 95056
rect 403716 94936 403768 94988
rect 414664 94936 414716 94988
rect 457720 94936 457772 94988
rect 468484 94936 468536 94988
rect 511724 94936 511776 94988
rect 522304 94936 522356 94988
rect 36544 94868 36596 94920
rect 538680 94868 538732 94920
rect 15292 91740 15344 91792
rect 529020 91740 529072 91792
rect 25688 91332 25740 91384
rect 149704 91332 149756 91384
rect 36544 91264 36596 91316
rect 52644 91264 52696 91316
rect 475016 91264 475068 91316
rect 494704 91264 494756 91316
rect 43076 91196 43128 91248
rect 62764 91196 62816 91248
rect 90456 91196 90508 91248
rect 106648 91196 106700 91248
rect 116492 91196 116544 91248
rect 133696 91196 133748 91248
rect 144276 91196 144328 91248
rect 160652 91196 160704 91248
rect 170496 91196 170548 91248
rect 187700 91196 187752 91248
rect 197452 91196 197504 91248
rect 214656 91196 214708 91248
rect 224500 91196 224552 91248
rect 241704 91196 241756 91248
rect 251456 91196 251508 91248
rect 268660 91196 268712 91248
rect 413468 91196 413520 91248
rect 430672 91196 430724 91248
rect 440516 91196 440568 91248
rect 457628 91196 457680 91248
rect 468484 91196 468536 91248
rect 484676 91196 484728 91248
rect 36820 91128 36872 91180
rect 62304 91128 62356 91180
rect 64144 91128 64196 91180
rect 89352 91128 89404 91180
rect 90364 91128 90416 91180
rect 116308 91128 116360 91180
rect 116584 91128 116636 91180
rect 143356 91128 143408 91180
rect 144184 91128 144236 91180
rect 170312 91128 170364 91180
rect 178040 91128 178092 91180
rect 200764 91128 200816 91180
rect 232044 91128 232096 91180
rect 251824 91128 251876 91180
rect 279424 91128 279476 91180
rect 295708 91128 295760 91180
rect 305460 91128 305512 91180
rect 322664 91128 322716 91180
rect 334624 91128 334676 91180
rect 349712 91128 349764 91180
rect 359464 91128 359516 91180
rect 376668 91128 376720 91180
rect 386512 91128 386564 91180
rect 403624 91128 403676 91180
rect 421012 91128 421064 91180
rect 443644 91128 443696 91180
rect 494520 91128 494572 91180
rect 511632 91128 511684 91180
rect 522304 91128 522356 91180
rect 538680 91128 538732 91180
rect 62488 91060 62540 91112
rect 79692 91060 79744 91112
rect 171784 91060 171836 91112
rect 197360 91060 197412 91112
rect 199384 91060 199436 91112
rect 224316 91060 224368 91112
rect 225604 91060 225656 91112
rect 251364 91060 251416 91112
rect 253204 91060 253256 91112
rect 278320 91060 278372 91112
rect 279516 91060 279568 91112
rect 305368 91060 305420 91112
rect 307024 91060 307076 91112
rect 332324 91060 332376 91112
rect 333244 91060 333296 91112
rect 359372 91060 359424 91112
rect 359556 91060 359608 91112
rect 386328 91060 386380 91112
rect 387064 91060 387116 91112
rect 413284 91060 413336 91112
rect 414664 91060 414716 91112
rect 440332 91060 440384 91112
rect 442264 91060 442316 91112
rect 467288 91060 467340 91112
rect 468576 91060 468628 91112
rect 494336 91060 494388 91112
rect 496084 91060 496136 91112
rect 521292 91060 521344 91112
rect 522396 91060 522448 91112
rect 548340 91060 548392 91112
rect 37924 90312 37976 90364
rect 526444 90312 526496 90364
rect 68928 88476 68980 88528
rect 118700 88476 118752 88528
rect 230388 88476 230440 88528
rect 280160 88476 280212 88528
rect 35624 88408 35676 88460
rect 36636 88408 36688 88460
rect 41328 88408 41380 88460
rect 91100 88408 91152 88460
rect 122748 88408 122800 88460
rect 172520 88408 172572 88460
rect 176568 88408 176620 88460
rect 226340 88408 226392 88460
rect 256608 88408 256660 88460
rect 307760 88408 307812 88460
rect 311808 88408 311860 88460
rect 361580 88408 361632 88460
rect 365628 88408 365680 88460
rect 415400 88408 415452 88460
rect 419448 88408 419500 88460
rect 469220 88408 469272 88460
rect 473268 88408 473320 88460
rect 523040 88408 523092 88460
rect 13728 88340 13780 88392
rect 64880 88340 64932 88392
rect 95148 88340 95200 88392
rect 146300 88340 146352 88392
rect 148968 88340 149020 88392
rect 200120 88340 200172 88392
rect 202788 88340 202840 88392
rect 253940 88340 253992 88392
rect 284208 88340 284260 88392
rect 335360 88340 335412 88392
rect 338028 88340 338080 88392
rect 389180 88340 389232 88392
rect 391848 88340 391900 88392
rect 443000 88340 443052 88392
rect 445668 88340 445720 88392
rect 496820 88340 496872 88392
rect 500868 88340 500920 88392
rect 550640 88340 550692 88392
rect 89720 72292 89772 72344
rect 90456 72292 90508 72344
rect 143632 72292 143684 72344
rect 144276 72292 144328 72344
rect 332508 71680 332560 71732
rect 334624 71680 334676 71732
rect 116216 70592 116268 70644
rect 116492 70592 116544 70644
rect 170220 70592 170272 70644
rect 170496 70592 170548 70644
rect 53104 68960 53156 69012
rect 64144 68960 64196 69012
rect 69112 68960 69164 69012
rect 15200 68892 15252 68944
rect 42800 68892 42852 68944
rect 62764 68892 62816 68944
rect 69756 68892 69808 68944
rect 96712 68960 96764 69012
rect 96804 68892 96856 68944
rect 146944 68960 146996 69012
rect 123668 68892 123720 68944
rect 133788 68892 133840 68944
rect 144184 68892 144236 68944
rect 25964 68824 26016 68876
rect 36820 68824 36872 68876
rect 79968 68824 80020 68876
rect 90364 68824 90416 68876
rect 106556 68824 106608 68876
rect 116584 68824 116636 68876
rect 122932 68824 122984 68876
rect 150716 68892 150768 68944
rect 200764 68960 200816 69012
rect 204628 68960 204680 69012
rect 251824 68960 251876 69012
rect 258724 68960 258776 69012
rect 443644 68960 443696 69012
rect 447692 68960 447744 69012
rect 494704 68960 494756 69012
rect 501604 68960 501656 69012
rect 548064 68892 548116 68944
rect 150532 68824 150584 68876
rect 178132 68824 178184 68876
rect 187976 68824 188028 68876
rect 199384 68824 199436 68876
rect 204352 68824 204404 68876
rect 231860 68824 231912 68876
rect 242072 68824 242124 68876
rect 253204 68824 253256 68876
rect 258172 68824 258224 68876
rect 160560 68756 160612 68808
rect 171784 68756 171836 68808
rect 215024 68756 215076 68808
rect 225604 68756 225656 68808
rect 268936 68756 268988 68808
rect 279516 68756 279568 68808
rect 285772 68824 285824 68876
rect 312636 68824 312688 68876
rect 286140 68756 286192 68808
rect 295984 68756 296036 68808
rect 307024 68756 307076 68808
rect 311992 68756 312044 68808
rect 340144 68824 340196 68876
rect 322848 68756 322900 68808
rect 333244 68756 333296 68808
rect 339592 68756 339644 68808
rect 350080 68756 350132 68808
rect 359556 68756 359608 68808
rect 365812 68824 365864 68876
rect 393596 68824 393648 68876
rect 366732 68756 366784 68808
rect 376576 68756 376628 68808
rect 387064 68756 387116 68808
rect 393412 68756 393464 68808
rect 420920 68824 420972 68876
rect 431040 68824 431092 68876
rect 442264 68824 442316 68876
rect 447232 68824 447284 68876
rect 474740 68824 474792 68876
rect 484952 68824 485004 68876
rect 496084 68824 496136 68876
rect 501052 68824 501104 68876
rect 528744 68824 528796 68876
rect 403992 68756 404044 68808
rect 414664 68756 414716 68808
rect 458088 68756 458140 68808
rect 468576 68756 468628 68808
rect 511908 68756 511960 68808
rect 522396 68756 522448 68808
rect 36728 68688 36780 68740
rect 538404 68688 538456 68740
rect 16304 65492 16356 65544
rect 528652 65492 528704 65544
rect 26056 65152 26108 65204
rect 146944 65152 146996 65204
rect 36728 65084 36780 65136
rect 52460 65084 52512 65136
rect 232320 65084 232372 65136
rect 251824 65084 251876 65136
rect 475384 65084 475436 65136
rect 494704 65084 494756 65136
rect 43352 65016 43404 65068
rect 62764 65016 62816 65068
rect 90456 65016 90508 65068
rect 106464 65016 106516 65068
rect 116492 65016 116544 65068
rect 133420 65016 133472 65068
rect 170496 65016 170548 65068
rect 187792 65016 187844 65068
rect 197544 65016 197596 65068
rect 214380 65016 214432 65068
rect 224500 65016 224552 65068
rect 241612 65016 241664 65068
rect 413468 65016 413520 65068
rect 430580 65016 430632 65068
rect 440516 65016 440568 65068
rect 457260 65016 457312 65068
rect 468576 65016 468628 65068
rect 484400 65016 484452 65068
rect 36820 64948 36872 65000
rect 62120 64948 62172 65000
rect 64144 64948 64196 65000
rect 89076 64948 89128 65000
rect 90364 64948 90416 65000
rect 116124 64948 116176 65000
rect 116584 64948 116636 65000
rect 142988 64948 143040 65000
rect 144276 64948 144328 65000
rect 170036 64948 170088 65000
rect 178408 64948 178460 65000
rect 200764 64948 200816 65000
rect 251456 64948 251508 65000
rect 268292 64948 268344 65000
rect 279424 64948 279476 65000
rect 295800 64948 295852 65000
rect 305552 64948 305604 65000
rect 322388 64948 322440 65000
rect 334624 64948 334676 65000
rect 349804 64948 349856 65000
rect 359648 64948 359700 65000
rect 376300 64948 376352 65000
rect 386512 64948 386564 65000
rect 403348 64948 403400 65000
rect 421288 64948 421340 65000
rect 443644 64948 443696 65000
rect 494520 64948 494572 65000
rect 511356 64948 511408 65000
rect 522304 64948 522356 65000
rect 538404 64948 538456 65000
rect 62488 64880 62540 64932
rect 79324 64880 79376 64932
rect 144184 64880 144236 64932
rect 160284 64880 160336 64932
rect 171784 64880 171836 64932
rect 197452 64880 197504 64932
rect 199384 64880 199436 64932
rect 223948 64880 224000 64932
rect 225604 64880 225656 64932
rect 251272 64880 251324 64932
rect 253204 64880 253256 64932
rect 278044 64880 278096 64932
rect 279516 64880 279568 64932
rect 305460 64880 305512 64932
rect 307024 64880 307076 64932
rect 331956 64880 332008 64932
rect 333244 64880 333296 64932
rect 359464 64880 359516 64932
rect 359556 64880 359608 64932
rect 386052 64880 386104 64932
rect 387064 64880 387116 64932
rect 412916 64880 412968 64932
rect 414664 64880 414716 64932
rect 440240 64880 440292 64932
rect 442264 64880 442316 64932
rect 467012 64880 467064 64932
rect 468484 64880 468536 64932
rect 494060 64880 494112 64932
rect 496084 64880 496136 64932
rect 520924 64880 520976 64932
rect 522396 64880 522448 64932
rect 547972 64880 548024 64932
rect 37924 62772 37976 62824
rect 526444 62772 526496 62824
rect 285772 62364 285824 62416
rect 286140 62364 286192 62416
rect 339592 62296 339644 62348
rect 340144 62296 340196 62348
rect 68928 62160 68980 62212
rect 118700 62160 118752 62212
rect 122748 62160 122800 62212
rect 172520 62160 172572 62212
rect 230388 62160 230440 62212
rect 280160 62160 280212 62212
rect 311808 62160 311860 62212
rect 361580 62160 361632 62212
rect 473268 62160 473320 62212
rect 523040 62160 523092 62212
rect 41328 62092 41380 62144
rect 91100 62092 91152 62144
rect 148968 62092 149020 62144
rect 200120 62092 200172 62144
rect 202788 62092 202840 62144
rect 253940 62092 253992 62144
rect 284208 62092 284260 62144
rect 335360 62092 335412 62144
rect 365628 62092 365680 62144
rect 415400 62092 415452 62144
rect 419448 62092 419500 62144
rect 469220 62092 469272 62144
rect 500868 62092 500920 62144
rect 550640 62092 550692 62144
rect 359556 60120 359608 60172
rect 359556 59916 359608 59968
rect 89720 50328 89772 50380
rect 90456 50328 90508 50380
rect 13728 44072 13780 44124
rect 64880 44072 64932 44124
rect 95148 44072 95200 44124
rect 146300 44072 146352 44124
rect 176568 44072 176620 44124
rect 226340 44072 226392 44124
rect 256608 44072 256660 44124
rect 307760 44072 307812 44124
rect 332508 44072 332560 44124
rect 334624 44072 334676 44124
rect 338028 44072 338080 44124
rect 389180 44072 389232 44124
rect 391848 44072 391900 44124
rect 443000 44072 443052 44124
rect 445668 44072 445720 44124
rect 496820 44072 496872 44124
rect 35624 44004 35676 44056
rect 36728 44004 36780 44056
rect 467656 44004 467708 44056
rect 468576 44004 468628 44056
rect 62764 41352 62816 41404
rect 70032 41352 70084 41404
rect 96712 41352 96764 41404
rect 15200 41284 15252 41336
rect 42984 41284 43036 41336
rect 52736 41284 52788 41336
rect 64144 41284 64196 41336
rect 69112 41284 69164 41336
rect 96988 41284 97040 41336
rect 200764 41352 200816 41404
rect 204996 41352 205048 41404
rect 251824 41352 251876 41404
rect 259000 41352 259052 41404
rect 443644 41352 443696 41404
rect 447968 41352 448020 41404
rect 494704 41352 494756 41404
rect 501972 41352 502024 41404
rect 124036 41284 124088 41336
rect 149704 41284 149756 41336
rect 548340 41284 548392 41336
rect 25688 41216 25740 41268
rect 36820 41216 36872 41268
rect 79692 41216 79744 41268
rect 90364 41216 90416 41268
rect 106648 41216 106700 41268
rect 116584 41216 116636 41268
rect 133696 41216 133748 41268
rect 144276 41216 144328 41268
rect 150532 41216 150584 41268
rect 178040 41216 178092 41268
rect 187700 41216 187752 41268
rect 199384 41216 199436 41268
rect 204352 41216 204404 41268
rect 232044 41216 232096 41268
rect 241704 41216 241756 41268
rect 253204 41216 253256 41268
rect 258172 41216 258224 41268
rect 286048 41216 286100 41268
rect 122932 41148 122984 41200
rect 150992 41148 151044 41200
rect 160652 41148 160704 41200
rect 171784 41148 171836 41200
rect 214656 41148 214708 41200
rect 225604 41148 225656 41200
rect 268660 41148 268712 41200
rect 279516 41148 279568 41200
rect 285772 41148 285824 41200
rect 313004 41216 313056 41268
rect 295708 41148 295760 41200
rect 307024 41148 307076 41200
rect 311992 41148 312044 41200
rect 340052 41216 340104 41268
rect 322664 41148 322716 41200
rect 333244 41148 333296 41200
rect 339592 41148 339644 41200
rect 367008 41216 367060 41268
rect 349712 41148 349764 41200
rect 359556 41148 359608 41200
rect 365812 41148 365864 41200
rect 393964 41216 394016 41268
rect 376668 41148 376720 41200
rect 387064 41148 387116 41200
rect 393412 41148 393464 41200
rect 421012 41216 421064 41268
rect 430672 41216 430724 41268
rect 442264 41216 442316 41268
rect 447232 41216 447284 41268
rect 475016 41216 475068 41268
rect 484676 41216 484728 41268
rect 496084 41216 496136 41268
rect 501052 41216 501104 41268
rect 529020 41216 529072 41268
rect 403716 41148 403768 41200
rect 414664 41148 414716 41200
rect 457720 41148 457772 41200
rect 468484 41148 468536 41200
rect 511724 41148 511776 41200
rect 522396 41148 522448 41200
rect 36636 41080 36688 41132
rect 538680 41080 538732 41132
rect 16028 38020 16080 38072
rect 529020 38020 529072 38072
rect 35348 37952 35400 38004
rect 580540 37952 580592 38004
rect 25688 37884 25740 37936
rect 580356 37884 580408 37936
rect 43076 37476 43128 37528
rect 62764 37476 62816 37528
rect 232044 37476 232096 37528
rect 251824 37476 251876 37528
rect 36636 37408 36688 37460
rect 52644 37408 52696 37460
rect 170496 37408 170548 37460
rect 187700 37408 187752 37460
rect 197452 37408 197504 37460
rect 214656 37408 214708 37460
rect 224500 37408 224552 37460
rect 241704 37408 241756 37460
rect 413468 37408 413520 37460
rect 430672 37408 430724 37460
rect 440516 37408 440568 37460
rect 457628 37408 457680 37460
rect 468484 37408 468536 37460
rect 484676 37408 484728 37460
rect 494520 37408 494572 37460
rect 511632 37408 511684 37460
rect 62488 37340 62540 37392
rect 79692 37340 79744 37392
rect 90364 37340 90416 37392
rect 106648 37340 106700 37392
rect 116492 37340 116544 37392
rect 133696 37340 133748 37392
rect 144184 37340 144236 37392
rect 160652 37340 160704 37392
rect 178040 37340 178092 37392
rect 200764 37340 200816 37392
rect 251456 37340 251508 37392
rect 268660 37340 268712 37392
rect 279424 37340 279476 37392
rect 295708 37340 295760 37392
rect 305460 37340 305512 37392
rect 322664 37340 322716 37392
rect 336004 37340 336056 37392
rect 349712 37340 349764 37392
rect 359464 37340 359516 37392
rect 376668 37340 376720 37392
rect 386512 37340 386564 37392
rect 403624 37340 403676 37392
rect 421012 37340 421064 37392
rect 446404 37340 446456 37392
rect 475016 37340 475068 37392
rect 494704 37340 494756 37392
rect 522396 37340 522448 37392
rect 538680 37340 538732 37392
rect 36728 37272 36780 37324
rect 62304 37272 62356 37324
rect 64144 37272 64196 37324
rect 89352 37272 89404 37324
rect 90456 37272 90508 37324
rect 116308 37272 116360 37324
rect 116584 37272 116636 37324
rect 143356 37272 143408 37324
rect 144276 37272 144328 37324
rect 170312 37272 170364 37324
rect 171784 37272 171836 37324
rect 197360 37272 197412 37324
rect 199384 37272 199436 37324
rect 224316 37272 224368 37324
rect 225604 37272 225656 37324
rect 251364 37272 251416 37324
rect 253204 37272 253256 37324
rect 278320 37272 278372 37324
rect 279516 37272 279568 37324
rect 305368 37272 305420 37324
rect 307024 37272 307076 37324
rect 332324 37272 332376 37324
rect 333244 37272 333296 37324
rect 359372 37272 359424 37324
rect 359556 37272 359608 37324
rect 386328 37272 386380 37324
rect 387064 37272 387116 37324
rect 413284 37272 413336 37324
rect 414664 37272 414716 37324
rect 440332 37272 440384 37324
rect 442264 37272 442316 37324
rect 467288 37272 467340 37324
rect 468576 37272 468628 37324
rect 494336 37272 494388 37324
rect 496084 37272 496136 37324
rect 521292 37272 521344 37324
rect 522304 37272 522356 37324
rect 548340 37272 548392 37324
rect 37924 36592 37976 36644
rect 526444 36592 526496 36644
rect 38016 36524 38068 36576
rect 580448 36524 580500 36576
rect 68928 34620 68980 34672
rect 118700 34620 118752 34672
rect 311808 34620 311860 34672
rect 361580 34620 361632 34672
rect 41328 34552 41380 34604
rect 91100 34552 91152 34604
rect 122748 34552 122800 34604
rect 172520 34552 172572 34604
rect 176568 34552 176620 34604
rect 226340 34552 226392 34604
rect 230388 34552 230440 34604
rect 280160 34552 280212 34604
rect 284208 34552 284260 34604
rect 335360 34552 335412 34604
rect 365628 34552 365680 34604
rect 415400 34552 415452 34604
rect 419448 34552 419500 34604
rect 469220 34552 469272 34604
rect 473268 34552 473320 34604
rect 523040 34552 523092 34604
rect 13728 34484 13780 34536
rect 64880 34484 64932 34536
rect 95148 34484 95200 34536
rect 146300 34484 146352 34536
rect 148968 34484 149020 34536
rect 200120 34484 200172 34536
rect 202788 34484 202840 34536
rect 253940 34484 253992 34536
rect 256608 34484 256660 34536
rect 307760 34484 307812 34536
rect 338028 34484 338080 34536
rect 389180 34484 389232 34536
rect 391848 34484 391900 34536
rect 443000 34484 443052 34536
rect 445668 34484 445720 34536
rect 496820 34484 496872 34536
rect 500868 34484 500920 34536
rect 550640 34484 550692 34536
rect 35624 16532 35676 16584
rect 36636 16532 36688 16584
rect 200764 16532 200816 16584
rect 204628 16532 204680 16584
rect 332508 16532 332560 16584
rect 336004 16532 336056 16584
rect 446404 16532 446456 16584
rect 447692 16532 447744 16584
rect 521752 16532 521804 16584
rect 522396 16532 522448 16584
rect 62764 13744 62816 13796
rect 69756 13744 69808 13796
rect 36544 13676 36596 13728
rect 146944 13676 146996 13728
rect 251824 13744 251876 13796
rect 258724 13744 258776 13796
rect 350080 13744 350132 13796
rect 359556 13744 359608 13796
rect 494704 13744 494756 13796
rect 501604 13744 501656 13796
rect 15200 13608 15252 13660
rect 42800 13608 42852 13660
rect 53104 13608 53156 13660
rect 64144 13608 64196 13660
rect 69112 13608 69164 13660
rect 96804 13608 96856 13660
rect 25964 13540 26016 13592
rect 36728 13540 36780 13592
rect 79968 13540 80020 13592
rect 90456 13540 90508 13592
rect 96712 13540 96764 13592
rect 123668 13608 123720 13660
rect 133788 13608 133840 13660
rect 144276 13608 144328 13660
rect 106556 13540 106608 13592
rect 116584 13540 116636 13592
rect 122932 13540 122984 13592
rect 150716 13608 150768 13660
rect 538404 13676 538456 13728
rect 548064 13608 548116 13660
rect 150532 13540 150584 13592
rect 178132 13540 178184 13592
rect 187976 13540 188028 13592
rect 199384 13540 199436 13592
rect 204352 13540 204404 13592
rect 231860 13540 231912 13592
rect 242072 13540 242124 13592
rect 253204 13540 253256 13592
rect 258172 13540 258224 13592
rect 160560 13472 160612 13524
rect 171784 13472 171836 13524
rect 215024 13472 215076 13524
rect 225604 13472 225656 13524
rect 268936 13472 268988 13524
rect 279516 13472 279568 13524
rect 285772 13540 285824 13592
rect 312636 13540 312688 13592
rect 286140 13472 286192 13524
rect 295984 13472 296036 13524
rect 307024 13472 307076 13524
rect 311992 13472 312044 13524
rect 340144 13540 340196 13592
rect 322848 13472 322900 13524
rect 333244 13472 333296 13524
rect 339592 13472 339644 13524
rect 365812 13540 365864 13592
rect 393596 13540 393648 13592
rect 366732 13472 366784 13524
rect 376576 13472 376628 13524
rect 387064 13472 387116 13524
rect 393412 13472 393464 13524
rect 420920 13540 420972 13592
rect 431040 13540 431092 13592
rect 442264 13540 442316 13592
rect 447232 13540 447284 13592
rect 474740 13540 474792 13592
rect 484952 13540 485004 13592
rect 496084 13540 496136 13592
rect 501052 13540 501104 13592
rect 528744 13540 528796 13592
rect 403992 13472 404044 13524
rect 414664 13472 414716 13524
rect 458088 13472 458140 13524
rect 468576 13472 468628 13524
rect 511908 13472 511960 13524
rect 522304 13472 522356 13524
rect 16304 13404 16356 13456
rect 580264 13404 580316 13456
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 25964 686180 26016 686186
rect 25964 686122 26016 686128
rect 149704 686180 149756 686186
rect 149704 686122 149756 686128
rect 25976 683890 26004 686122
rect 36636 686112 36688 686118
rect 36636 686054 36688 686060
rect 52460 686112 52512 686118
rect 52460 686054 52512 686060
rect 25714 683862 26004 683890
rect 15212 683318 16054 683346
rect 35374 683318 35848 683346
rect 13726 674248 13782 674257
rect 13726 674183 13782 674192
rect 13740 665174 13768 674183
rect 13728 665168 13780 665174
rect 13728 665110 13780 665116
rect 15212 662250 15240 683318
rect 35820 683210 35848 683318
rect 35820 683182 35940 683210
rect 35912 683114 35940 683182
rect 35912 683086 36584 683114
rect 35624 665100 35676 665106
rect 35624 665042 35676 665048
rect 35636 664714 35664 665042
rect 35374 664686 35664 664714
rect 15200 662244 15252 662250
rect 15200 662186 15252 662192
rect 16040 658986 16068 664020
rect 25700 662318 25728 664020
rect 25688 662312 25740 662318
rect 25688 662254 25740 662260
rect 16028 658980 16080 658986
rect 16028 658922 16080 658928
rect 25688 658572 25740 658578
rect 25688 658514 25740 658520
rect 25700 656948 25728 658514
rect 35374 656946 35664 656962
rect 35374 656940 35676 656946
rect 35374 656934 35624 656940
rect 35624 656882 35676 656888
rect 15212 656254 16054 656282
rect 13728 655580 13780 655586
rect 13728 655522 13780 655528
rect 13740 647329 13768 655522
rect 13726 647320 13782 647329
rect 13726 647255 13782 647264
rect 15212 634710 15240 656254
rect 35624 637560 35676 637566
rect 35374 637508 35624 637514
rect 35374 637502 35676 637508
rect 35374 637486 35664 637502
rect 16054 637078 16344 637106
rect 25714 637078 26096 637106
rect 15200 634704 15252 634710
rect 15200 634646 15252 634652
rect 16316 632738 16344 637078
rect 26068 634642 26096 637078
rect 26056 634636 26108 634642
rect 26056 634578 26108 634584
rect 36556 634506 36584 683086
rect 36648 665106 36676 686054
rect 36728 685976 36780 685982
rect 36728 685918 36780 685924
rect 36636 665100 36688 665106
rect 36636 665042 36688 665048
rect 36740 662318 36768 685918
rect 43352 685908 43404 685914
rect 43352 685850 43404 685856
rect 43364 683890 43392 685850
rect 43102 683862 43392 683890
rect 52472 683890 52500 686054
rect 62488 686044 62540 686050
rect 62488 685986 62540 685992
rect 79324 686044 79376 686050
rect 79324 685986 79376 685992
rect 90364 686044 90416 686050
rect 90364 685986 90416 685992
rect 106372 686044 106424 686050
rect 106372 685986 106424 685992
rect 116492 686044 116544 686050
rect 116492 685986 116544 685992
rect 133420 686044 133472 686050
rect 133420 685986 133472 685992
rect 144276 686044 144328 686050
rect 144276 685986 144328 685992
rect 62120 685976 62172 685982
rect 62120 685918 62172 685924
rect 62132 683890 62160 685918
rect 52472 683862 52670 683890
rect 62132 683862 62330 683890
rect 41328 683188 41380 683194
rect 41328 683130 41380 683136
rect 41340 674393 41368 683130
rect 41326 674384 41382 674393
rect 41326 674319 41382 674328
rect 37922 673840 37978 673849
rect 37922 673775 37978 673784
rect 36728 662312 36780 662318
rect 36728 662254 36780 662260
rect 36728 658504 36780 658510
rect 36728 658446 36780 658452
rect 36636 656940 36688 656946
rect 36636 656882 36688 656888
rect 36544 634500 36596 634506
rect 36544 634442 36596 634448
rect 16304 632732 16356 632738
rect 16304 632674 16356 632680
rect 25964 632392 26016 632398
rect 25964 632334 26016 632340
rect 25976 629898 26004 632334
rect 25714 629870 26004 629898
rect 15212 629326 16054 629354
rect 35374 629326 35940 629354
rect 13726 620256 13782 620265
rect 13726 620191 13782 620200
rect 13740 611318 13768 620191
rect 13728 611312 13780 611318
rect 13728 611254 13780 611260
rect 15212 608530 15240 629326
rect 35912 625154 35940 629326
rect 35912 625126 36584 625154
rect 35624 611244 35676 611250
rect 35624 611186 35676 611192
rect 35636 610722 35664 611186
rect 35374 610694 35664 610722
rect 15304 610014 16054 610042
rect 15200 608524 15252 608530
rect 15200 608466 15252 608472
rect 15304 605130 15332 610014
rect 25700 608462 25728 610028
rect 25688 608456 25740 608462
rect 25688 608398 25740 608404
rect 15292 605124 15344 605130
rect 15292 605066 15344 605072
rect 25688 604784 25740 604790
rect 25688 604726 25740 604732
rect 25700 602956 25728 604726
rect 15212 602262 16054 602290
rect 35374 602262 35664 602290
rect 13726 593192 13782 593201
rect 13726 593127 13782 593136
rect 13740 583710 13768 593127
rect 13728 583704 13780 583710
rect 13728 583646 13780 583652
rect 15212 580922 15240 602262
rect 35636 601730 35664 602262
rect 35624 601724 35676 601730
rect 35624 601666 35676 601672
rect 35374 583642 35664 583658
rect 35374 583636 35676 583642
rect 35374 583630 35624 583636
rect 35624 583578 35676 583584
rect 16054 583086 16344 583114
rect 25714 583086 26004 583114
rect 15200 580916 15252 580922
rect 15200 580858 15252 580864
rect 16316 578950 16344 583086
rect 25976 580854 26004 583086
rect 25964 580848 26016 580854
rect 25964 580790 26016 580796
rect 36556 580718 36584 625126
rect 36648 608326 36676 656882
rect 36740 637566 36768 658446
rect 36820 658368 36872 658374
rect 36820 658310 36872 658316
rect 36728 637560 36780 637566
rect 36728 637502 36780 637508
rect 36832 634642 36860 658310
rect 37936 657558 37964 673775
rect 62500 664714 62528 685986
rect 64144 685976 64196 685982
rect 64144 685918 64196 685924
rect 62764 685908 62816 685914
rect 62764 685850 62816 685856
rect 62422 664686 62528 664714
rect 42996 662250 43024 664020
rect 52762 664006 53144 664034
rect 53116 662318 53144 664006
rect 62776 662386 62804 685850
rect 62764 662380 62816 662386
rect 62764 662322 62816 662328
rect 64156 662318 64184 685918
rect 79336 683890 79364 685986
rect 89076 685976 89128 685982
rect 89076 685918 89128 685924
rect 89088 683890 89116 685918
rect 79336 683862 79718 683890
rect 89088 683862 89378 683890
rect 69124 683318 70058 683346
rect 68928 683256 68980 683262
rect 68928 683198 68980 683204
rect 68940 674801 68968 683198
rect 68926 674792 68982 674801
rect 68926 674727 68982 674736
rect 64878 673568 64934 673577
rect 64878 673503 64934 673512
rect 64892 665174 64920 673503
rect 64880 665168 64932 665174
rect 64880 665110 64932 665116
rect 53104 662312 53156 662318
rect 53104 662254 53156 662260
rect 64144 662312 64196 662318
rect 64144 662254 64196 662260
rect 69124 662250 69152 683318
rect 90376 673454 90404 685986
rect 90456 685976 90508 685982
rect 90456 685918 90508 685924
rect 89824 673426 90404 673454
rect 89824 664714 89852 673426
rect 89378 664686 89852 664714
rect 70044 662386 70072 664020
rect 70032 662380 70084 662386
rect 70032 662322 70084 662328
rect 79704 662318 79732 664020
rect 90468 662318 90496 685918
rect 106384 683890 106412 685986
rect 115940 685976 115992 685982
rect 115940 685918 115992 685924
rect 115952 683890 115980 685918
rect 106384 683862 106674 683890
rect 115952 683862 116334 683890
rect 96724 683318 97014 683346
rect 91100 683188 91152 683194
rect 91100 683130 91152 683136
rect 91112 673713 91140 683130
rect 95146 674248 95202 674257
rect 95146 674183 95202 674192
rect 91098 673704 91154 673713
rect 91098 673639 91154 673648
rect 95160 665174 95188 674183
rect 95148 665168 95200 665174
rect 95148 665110 95200 665116
rect 96724 662386 96752 683318
rect 96712 662380 96764 662386
rect 96712 662322 96764 662328
rect 79692 662312 79744 662318
rect 79692 662254 79744 662260
rect 90456 662312 90508 662318
rect 90456 662254 90508 662260
rect 97000 662250 97028 664020
rect 106660 662318 106688 664020
rect 116320 663898 116348 664020
rect 116504 663898 116532 685986
rect 116584 685976 116636 685982
rect 116584 685918 116636 685924
rect 116320 663870 116532 663898
rect 116596 662318 116624 685918
rect 133432 683890 133460 685986
rect 142988 685976 143040 685982
rect 142988 685918 143040 685924
rect 144184 685976 144236 685982
rect 144184 685918 144236 685924
rect 143000 683890 143028 685918
rect 133432 683862 133722 683890
rect 143000 683862 143382 683890
rect 122944 683318 124062 683346
rect 118700 683256 118752 683262
rect 118700 683198 118752 683204
rect 122748 683256 122800 683262
rect 122748 683198 122800 683204
rect 118712 673713 118740 683198
rect 122760 674393 122788 683198
rect 122746 674384 122802 674393
rect 122746 674319 122802 674328
rect 118698 673704 118754 673713
rect 118698 673639 118754 673648
rect 106648 662312 106700 662318
rect 106648 662254 106700 662260
rect 116584 662312 116636 662318
rect 116584 662254 116636 662260
rect 122944 662250 122972 683318
rect 143632 666188 143684 666194
rect 143632 666130 143684 666136
rect 143644 664714 143672 666130
rect 143382 664686 143672 664714
rect 124048 662386 124076 664020
rect 124036 662380 124088 662386
rect 124036 662322 124088 662328
rect 133708 662318 133736 664020
rect 144196 662318 144224 685918
rect 144288 666194 144316 685986
rect 148968 683188 149020 683194
rect 148968 683130 149020 683136
rect 148980 674393 149008 683130
rect 148966 674384 149022 674393
rect 148966 674319 149022 674328
rect 146298 673568 146354 673577
rect 146298 673503 146354 673512
rect 144276 666188 144328 666194
rect 144276 666130 144328 666136
rect 146312 665174 146340 673503
rect 146300 665168 146352 665174
rect 146300 665110 146352 665116
rect 133696 662312 133748 662318
rect 133696 662254 133748 662260
rect 144184 662312 144236 662318
rect 144184 662254 144236 662260
rect 42984 662244 43036 662250
rect 42984 662186 43036 662192
rect 69112 662244 69164 662250
rect 69112 662186 69164 662192
rect 96988 662244 97040 662250
rect 96988 662186 97040 662192
rect 122932 662244 122984 662250
rect 122932 662186 122984 662192
rect 146944 658572 146996 658578
rect 146944 658514 146996 658520
rect 52644 658504 52696 658510
rect 52644 658446 52696 658452
rect 43076 658300 43128 658306
rect 43076 658242 43128 658248
rect 37924 657552 37976 657558
rect 37924 657494 37976 657500
rect 43088 656948 43116 658242
rect 52656 656948 52684 658446
rect 62488 658436 62540 658442
rect 62488 658378 62540 658384
rect 79692 658436 79744 658442
rect 79692 658378 79744 658384
rect 90456 658436 90508 658442
rect 90456 658378 90508 658384
rect 106648 658436 106700 658442
rect 106648 658378 106700 658384
rect 116492 658436 116544 658442
rect 116492 658378 116544 658384
rect 133696 658436 133748 658442
rect 133696 658378 133748 658384
rect 62304 658368 62356 658374
rect 62304 658310 62356 658316
rect 62316 656948 62344 658310
rect 41328 655648 41380 655654
rect 41328 655590 41380 655596
rect 41340 647329 41368 655590
rect 41326 647320 41382 647329
rect 41326 647255 41382 647264
rect 37922 645960 37978 645969
rect 37922 645895 37978 645904
rect 36820 634636 36872 634642
rect 36820 634578 36872 634584
rect 36728 632324 36780 632330
rect 36728 632266 36780 632272
rect 36740 611250 36768 632266
rect 36820 632188 36872 632194
rect 36820 632130 36872 632136
rect 36728 611244 36780 611250
rect 36728 611186 36780 611192
rect 36832 608462 36860 632130
rect 37936 629950 37964 645895
rect 62500 637786 62528 658378
rect 64144 658368 64196 658374
rect 64144 658310 64196 658316
rect 62764 658300 62816 658306
rect 62764 658242 62816 658248
rect 62422 637758 62528 637786
rect 42812 637078 43010 637106
rect 52762 637078 53144 637106
rect 42812 634710 42840 637078
rect 53116 634710 53144 637078
rect 62776 634778 62804 658242
rect 62764 634772 62816 634778
rect 62764 634714 62816 634720
rect 64156 634710 64184 658310
rect 79704 656948 79732 658378
rect 89352 658368 89404 658374
rect 89352 658310 89404 658316
rect 90364 658368 90416 658374
rect 90364 658310 90416 658316
rect 89364 656948 89392 658310
rect 69124 656254 70058 656282
rect 68928 655716 68980 655722
rect 68928 655658 68980 655664
rect 64880 655580 64932 655586
rect 64880 655522 64932 655528
rect 64892 646649 64920 655522
rect 68940 647873 68968 655658
rect 68926 647864 68982 647873
rect 68926 647799 68982 647808
rect 64878 646640 64934 646649
rect 64878 646575 64934 646584
rect 69124 634710 69152 656254
rect 89720 637560 89772 637566
rect 89378 637508 89720 637514
rect 89378 637502 89772 637508
rect 89378 637486 89760 637502
rect 69768 637078 70058 637106
rect 79718 637078 80008 637106
rect 69768 634778 69796 637078
rect 69756 634772 69808 634778
rect 69756 634714 69808 634720
rect 42800 634704 42852 634710
rect 42800 634646 42852 634652
rect 53104 634704 53156 634710
rect 53104 634646 53156 634652
rect 64144 634704 64196 634710
rect 64144 634646 64196 634652
rect 69112 634704 69164 634710
rect 69112 634646 69164 634652
rect 79980 634642 80008 637078
rect 90376 634642 90404 658310
rect 90468 637566 90496 658378
rect 106660 656948 106688 658378
rect 116308 658368 116360 658374
rect 116308 658310 116360 658316
rect 116320 656948 116348 658310
rect 96724 656254 97014 656282
rect 91100 655648 91152 655654
rect 91100 655590 91152 655596
rect 91112 646649 91140 655590
rect 96620 655580 96672 655586
rect 96620 655522 96672 655528
rect 96632 654090 96660 655522
rect 95148 654084 95200 654090
rect 95148 654026 95200 654032
rect 96620 654084 96672 654090
rect 96620 654026 96672 654032
rect 95160 647329 95188 654026
rect 95146 647320 95202 647329
rect 95146 647255 95202 647264
rect 91098 646640 91154 646649
rect 91098 646575 91154 646584
rect 90456 637560 90508 637566
rect 90456 637502 90508 637508
rect 96724 634778 96752 656254
rect 96816 637078 97014 637106
rect 106568 637078 106674 637106
rect 116228 637078 116334 637106
rect 96712 634772 96764 634778
rect 96712 634714 96764 634720
rect 96816 634710 96844 637078
rect 96804 634704 96856 634710
rect 96804 634646 96856 634652
rect 106568 634642 106596 637078
rect 116228 636970 116256 637078
rect 116504 636970 116532 658378
rect 116584 658368 116636 658374
rect 116584 658310 116636 658316
rect 116228 636942 116532 636970
rect 116596 634642 116624 658310
rect 133708 656948 133736 658378
rect 143356 658368 143408 658374
rect 143356 658310 143408 658316
rect 144276 658368 144328 658374
rect 144276 658310 144328 658316
rect 143368 656948 143396 658310
rect 144184 658300 144236 658306
rect 144184 658242 144236 658248
rect 122944 656254 124062 656282
rect 118700 655716 118752 655722
rect 118700 655658 118752 655664
rect 118712 646649 118740 655658
rect 122748 655648 122800 655654
rect 122748 655590 122800 655596
rect 122760 647329 122788 655590
rect 122746 647320 122802 647329
rect 122746 647255 122802 647264
rect 118698 646640 118754 646649
rect 118698 646575 118754 646584
rect 79968 634636 80020 634642
rect 79968 634578 80020 634584
rect 90364 634636 90416 634642
rect 90364 634578 90416 634584
rect 106556 634636 106608 634642
rect 106556 634578 106608 634584
rect 116584 634636 116636 634642
rect 116584 634578 116636 634584
rect 122944 634574 122972 656254
rect 144196 644474 144224 658242
rect 143736 644446 144224 644474
rect 143736 637786 143764 644446
rect 143382 637758 143764 637786
rect 123680 637078 124062 637106
rect 133722 637078 133828 637106
rect 123680 634710 123708 637078
rect 123668 634704 123720 634710
rect 123668 634646 123720 634652
rect 133800 634642 133828 637078
rect 144288 634642 144316 658310
rect 146300 655580 146352 655586
rect 146300 655522 146352 655528
rect 146312 647193 146340 655522
rect 146298 647184 146354 647193
rect 146298 647119 146354 647128
rect 133788 634636 133840 634642
rect 133788 634578 133840 634584
rect 144276 634636 144328 634642
rect 144276 634578 144328 634584
rect 122932 634568 122984 634574
rect 122932 634510 122984 634516
rect 52460 632324 52512 632330
rect 52460 632266 52512 632272
rect 43352 632120 43404 632126
rect 43352 632062 43404 632068
rect 37924 629944 37976 629950
rect 43364 629898 43392 632062
rect 37924 629886 37976 629892
rect 43102 629870 43392 629898
rect 52472 629898 52500 632266
rect 62488 632256 62540 632262
rect 62488 632198 62540 632204
rect 79324 632256 79376 632262
rect 79324 632198 79376 632204
rect 90364 632256 90416 632262
rect 90364 632198 90416 632204
rect 106372 632256 106424 632262
rect 106372 632198 106424 632204
rect 116492 632256 116544 632262
rect 116492 632198 116544 632204
rect 133420 632256 133472 632262
rect 133420 632198 133472 632204
rect 62120 632188 62172 632194
rect 62120 632130 62172 632136
rect 62132 629898 62160 632130
rect 52472 629870 52670 629898
rect 62132 629870 62330 629898
rect 41326 620256 41382 620265
rect 41326 620191 41382 620200
rect 37922 619032 37978 619041
rect 37922 618967 37978 618976
rect 36820 608456 36872 608462
rect 36820 608398 36872 608404
rect 36636 608320 36688 608326
rect 36636 608262 36688 608268
rect 36728 604716 36780 604722
rect 36728 604658 36780 604664
rect 36636 601724 36688 601730
rect 36636 601666 36688 601672
rect 36544 580712 36596 580718
rect 36544 580654 36596 580660
rect 16304 578944 16356 578950
rect 16304 578886 16356 578892
rect 26056 578536 26108 578542
rect 26056 578478 26108 578484
rect 26068 575906 26096 578478
rect 25714 575878 26096 575906
rect 35374 575470 35940 575498
rect 15212 575334 16054 575362
rect 13726 566264 13782 566273
rect 13726 566199 13782 566208
rect 13740 557530 13768 566199
rect 13728 557524 13780 557530
rect 13728 557466 13780 557472
rect 15212 554674 15240 575334
rect 35912 567194 35940 575470
rect 35912 567166 36584 567194
rect 35624 557456 35676 557462
rect 35624 557398 35676 557404
rect 35636 556730 35664 557398
rect 35374 556702 35664 556730
rect 15200 554668 15252 554674
rect 15200 554610 15252 554616
rect 16040 551342 16068 556036
rect 25700 554606 25728 556036
rect 25688 554600 25740 554606
rect 25688 554542 25740 554548
rect 16028 551336 16080 551342
rect 16028 551278 16080 551284
rect 25688 550928 25740 550934
rect 25688 550870 25740 550876
rect 25700 548964 25728 550870
rect 15212 548270 16054 548298
rect 35374 548270 35664 548298
rect 13726 539200 13782 539209
rect 13726 539135 13782 539144
rect 13740 529922 13768 539135
rect 13728 529916 13780 529922
rect 13728 529858 13780 529864
rect 15212 527066 15240 548270
rect 35636 547942 35664 548270
rect 35624 547936 35676 547942
rect 35624 547878 35676 547884
rect 35624 529848 35676 529854
rect 35624 529790 35676 529796
rect 35636 529666 35664 529790
rect 35374 529638 35664 529666
rect 16054 529094 16344 529122
rect 25714 529094 26096 529122
rect 15200 527060 15252 527066
rect 15200 527002 15252 527008
rect 16316 523734 16344 529094
rect 26068 526998 26096 529094
rect 26056 526992 26108 526998
rect 26056 526934 26108 526940
rect 36556 526862 36584 567166
rect 36648 554470 36676 601666
rect 36740 583642 36768 604658
rect 36820 604580 36872 604586
rect 36820 604522 36872 604528
rect 36728 583636 36780 583642
rect 36728 583578 36780 583584
rect 36832 580854 36860 604522
rect 37936 602410 37964 618967
rect 41340 611250 41368 620191
rect 41328 611244 41380 611250
rect 41328 611186 41380 611192
rect 62500 610722 62528 632198
rect 64144 632188 64196 632194
rect 64144 632130 64196 632136
rect 62764 632120 62816 632126
rect 62764 632062 62816 632068
rect 62422 610694 62528 610722
rect 42996 608530 43024 610028
rect 52748 608598 52776 610028
rect 52736 608592 52788 608598
rect 52736 608534 52788 608540
rect 62776 608530 62804 632062
rect 64156 608598 64184 632130
rect 79336 629898 79364 632198
rect 89076 632188 89128 632194
rect 89076 632130 89128 632136
rect 89088 629898 89116 632130
rect 79336 629870 79718 629898
rect 89088 629870 89378 629898
rect 69124 629326 70058 629354
rect 68926 619712 68982 619721
rect 68926 619647 68982 619656
rect 64878 619576 64934 619585
rect 64878 619511 64934 619520
rect 64892 611318 64920 619511
rect 64880 611312 64932 611318
rect 64880 611254 64932 611260
rect 68940 611182 68968 619647
rect 68928 611176 68980 611182
rect 68928 611118 68980 611124
rect 69124 608598 69152 629326
rect 90376 615494 90404 632198
rect 90456 632188 90508 632194
rect 90456 632130 90508 632136
rect 89824 615466 90404 615494
rect 89824 610722 89852 615466
rect 89378 610694 89852 610722
rect 64144 608592 64196 608598
rect 64144 608534 64196 608540
rect 69112 608592 69164 608598
rect 69112 608534 69164 608540
rect 70044 608530 70072 610028
rect 42984 608524 43036 608530
rect 42984 608466 43036 608472
rect 62764 608524 62816 608530
rect 62764 608466 62816 608472
rect 70032 608524 70084 608530
rect 70032 608466 70084 608472
rect 79704 608462 79732 610028
rect 90468 608462 90496 632130
rect 106384 629898 106412 632198
rect 115940 632188 115992 632194
rect 115940 632130 115992 632136
rect 115952 629898 115980 632130
rect 106384 629870 106674 629898
rect 115952 629870 116334 629898
rect 96724 629326 97014 629354
rect 95146 620256 95202 620265
rect 95146 620191 95202 620200
rect 91098 619576 91154 619585
rect 91098 619511 91154 619520
rect 91112 611250 91140 619511
rect 95160 611318 95188 620191
rect 95148 611312 95200 611318
rect 95148 611254 95200 611260
rect 91100 611244 91152 611250
rect 91100 611186 91152 611192
rect 96724 608598 96752 629326
rect 96712 608592 96764 608598
rect 96712 608534 96764 608540
rect 97000 608530 97028 610028
rect 96988 608524 97040 608530
rect 96988 608466 97040 608472
rect 106660 608462 106688 610028
rect 116320 609906 116348 610028
rect 116504 609906 116532 632198
rect 116584 632188 116636 632194
rect 116584 632130 116636 632136
rect 116320 609878 116532 609906
rect 116596 608462 116624 632130
rect 133432 629898 133460 632198
rect 142988 632188 143040 632194
rect 142988 632130 143040 632136
rect 144276 632188 144328 632194
rect 144276 632130 144328 632136
rect 143000 629898 143028 632130
rect 144184 632120 144236 632126
rect 144184 632062 144236 632068
rect 133432 629870 133722 629898
rect 143000 629870 143382 629898
rect 122944 629326 124062 629354
rect 122746 620256 122802 620265
rect 122746 620191 122802 620200
rect 118698 619576 118754 619585
rect 118698 619511 118754 619520
rect 118712 611182 118740 619511
rect 122760 611250 122788 620191
rect 122748 611244 122800 611250
rect 122748 611186 122800 611192
rect 118700 611176 118752 611182
rect 118700 611118 118752 611124
rect 122944 608462 122972 629326
rect 144196 615494 144224 632062
rect 143736 615466 144224 615494
rect 143736 610722 143764 615466
rect 143382 610694 143764 610722
rect 124048 608530 124076 610028
rect 133708 608530 133736 610028
rect 144288 608530 144316 632130
rect 146298 619032 146354 619041
rect 146298 618967 146354 618976
rect 146312 611318 146340 618967
rect 146300 611312 146352 611318
rect 146300 611254 146352 611260
rect 146956 608598 146984 658514
rect 148968 655580 149020 655586
rect 148968 655522 149020 655528
rect 148980 647329 149008 655522
rect 148966 647320 149022 647329
rect 148966 647255 149022 647264
rect 149716 634710 149744 686122
rect 232320 686112 232372 686118
rect 232320 686054 232372 686060
rect 251824 686112 251876 686118
rect 251824 686054 251876 686060
rect 160284 686044 160336 686050
rect 160284 685986 160336 685992
rect 170496 686044 170548 686050
rect 170496 685986 170548 685992
rect 187792 686044 187844 686050
rect 187792 685986 187844 685992
rect 197544 686044 197596 686050
rect 197544 685986 197596 685992
rect 214380 686044 214432 686050
rect 214380 685986 214432 685992
rect 224500 686044 224552 686050
rect 224500 685986 224552 685992
rect 160296 683890 160324 685986
rect 170036 685976 170088 685982
rect 170036 685918 170088 685924
rect 170048 683890 170076 685918
rect 160296 683862 160678 683890
rect 170048 683862 170338 683890
rect 150544 683318 151018 683346
rect 150544 662386 150572 683318
rect 150532 662380 150584 662386
rect 150532 662322 150584 662328
rect 151004 662250 151032 664020
rect 160664 662318 160692 664020
rect 170324 663898 170352 664020
rect 170508 663898 170536 685986
rect 178408 685976 178460 685982
rect 178408 685918 178460 685924
rect 171784 685908 171836 685914
rect 171784 685850 171836 685856
rect 170324 663870 170536 663898
rect 171796 662318 171824 685850
rect 178420 683890 178448 685918
rect 187804 683890 187832 685986
rect 197452 685908 197504 685914
rect 197452 685850 197504 685856
rect 197464 683890 197492 685850
rect 178066 683862 178448 683890
rect 187726 683862 187832 683890
rect 197386 683862 197492 683890
rect 172520 683256 172572 683262
rect 172520 683198 172572 683204
rect 172532 673713 172560 683198
rect 176566 673840 176622 673849
rect 176566 673775 176622 673784
rect 172518 673704 172574 673713
rect 172518 673639 172574 673648
rect 176580 665174 176608 673775
rect 176568 665168 176620 665174
rect 176568 665110 176620 665116
rect 197556 664714 197584 685986
rect 200764 685976 200816 685982
rect 200764 685918 200816 685924
rect 199384 685908 199436 685914
rect 199384 685850 199436 685856
rect 197386 664686 197584 664714
rect 178052 662386 178080 664020
rect 187712 662386 187740 664020
rect 199396 662386 199424 685850
rect 200120 683188 200172 683194
rect 200120 683130 200172 683136
rect 200132 673713 200160 683130
rect 200118 673704 200174 673713
rect 200118 673639 200174 673648
rect 200776 662386 200804 685918
rect 214392 683890 214420 685986
rect 223948 685908 224000 685914
rect 223948 685850 224000 685856
rect 223960 683890 223988 685850
rect 214392 683862 214682 683890
rect 223960 683862 224342 683890
rect 204364 683318 205022 683346
rect 202788 683188 202840 683194
rect 202788 683130 202840 683136
rect 202800 674393 202828 683130
rect 202786 674384 202842 674393
rect 202786 674319 202842 674328
rect 178040 662380 178092 662386
rect 178040 662322 178092 662328
rect 187700 662380 187752 662386
rect 187700 662322 187752 662328
rect 199384 662380 199436 662386
rect 199384 662322 199436 662328
rect 200764 662380 200816 662386
rect 200764 662322 200816 662328
rect 204364 662318 204392 683318
rect 224512 664714 224540 685986
rect 225604 685908 225656 685914
rect 225604 685850 225656 685856
rect 224342 664686 224540 664714
rect 205008 662386 205036 664020
rect 204996 662380 205048 662386
rect 204996 662322 205048 662328
rect 214668 662318 214696 664020
rect 225616 662318 225644 685850
rect 232332 683890 232360 686054
rect 241520 686044 241572 686050
rect 241520 685986 241572 685992
rect 232070 683862 232360 683890
rect 241532 683890 241560 685986
rect 251456 685976 251508 685982
rect 251456 685918 251508 685924
rect 251180 685908 251232 685914
rect 251180 685850 251232 685856
rect 251192 683890 251220 685850
rect 241532 683862 241730 683890
rect 251192 683862 251390 683890
rect 230388 683256 230440 683262
rect 230388 683198 230440 683204
rect 230400 674393 230428 683198
rect 230386 674384 230442 674393
rect 230386 674319 230442 674328
rect 226338 673568 226394 673577
rect 226338 673503 226394 673512
rect 226352 665174 226380 673503
rect 226340 665168 226392 665174
rect 226340 665110 226392 665116
rect 251468 664714 251496 685918
rect 251390 664686 251496 664714
rect 232056 662386 232084 664020
rect 232044 662380 232096 662386
rect 232044 662322 232096 662328
rect 241716 662318 241744 664020
rect 251836 662386 251864 686054
rect 413468 686044 413520 686050
rect 413468 685986 413520 685992
rect 430580 686044 430632 686050
rect 430580 685986 430632 685992
rect 440516 686044 440568 686050
rect 440516 685986 440568 685992
rect 457260 686044 457312 686050
rect 457260 685986 457312 685992
rect 468576 686044 468628 686050
rect 468576 685986 468628 685992
rect 484400 686044 484452 686050
rect 484400 685986 484452 685992
rect 494520 686044 494572 686050
rect 494520 685986 494572 685992
rect 511356 686044 511408 686050
rect 511356 685986 511408 685992
rect 268292 685976 268344 685982
rect 268292 685918 268344 685924
rect 279424 685976 279476 685982
rect 279424 685918 279476 685924
rect 295800 685976 295852 685982
rect 295800 685918 295852 685924
rect 305552 685976 305604 685982
rect 305552 685918 305604 685924
rect 322388 685976 322440 685982
rect 322388 685918 322440 685924
rect 334624 685976 334676 685982
rect 334624 685918 334676 685924
rect 349804 685976 349856 685982
rect 349804 685918 349856 685924
rect 359648 685976 359700 685982
rect 359648 685918 359700 685924
rect 376300 685976 376352 685982
rect 376300 685918 376352 685924
rect 386512 685976 386564 685982
rect 386512 685918 386564 685924
rect 403348 685976 403400 685982
rect 403348 685918 403400 685924
rect 253204 685908 253256 685914
rect 253204 685850 253256 685856
rect 251824 662380 251876 662386
rect 251824 662322 251876 662328
rect 253216 662318 253244 685850
rect 268304 683890 268332 685918
rect 278044 685908 278096 685914
rect 278044 685850 278096 685856
rect 278056 683890 278084 685850
rect 268304 683862 268686 683890
rect 278056 683862 278346 683890
rect 258184 683318 259026 683346
rect 253940 683188 253992 683194
rect 253940 683130 253992 683136
rect 253952 674257 253980 683130
rect 253938 674248 253994 674257
rect 253938 674183 253994 674192
rect 256606 674248 256662 674257
rect 256606 674183 256662 674192
rect 256620 665174 256648 674183
rect 256608 665168 256660 665174
rect 256608 665110 256660 665116
rect 160652 662312 160704 662318
rect 160652 662254 160704 662260
rect 171784 662312 171836 662318
rect 171784 662254 171836 662260
rect 204352 662312 204404 662318
rect 204352 662254 204404 662260
rect 214656 662312 214708 662318
rect 214656 662254 214708 662260
rect 225604 662312 225656 662318
rect 225604 662254 225656 662260
rect 241704 662312 241756 662318
rect 241704 662254 241756 662260
rect 253204 662312 253256 662318
rect 253204 662254 253256 662260
rect 258184 662250 258212 683318
rect 279436 673454 279464 685918
rect 279516 685908 279568 685914
rect 279516 685850 279568 685856
rect 278792 673426 279464 673454
rect 278792 664714 278820 673426
rect 278346 664686 278820 664714
rect 259012 662386 259040 664020
rect 259000 662380 259052 662386
rect 259000 662322 259052 662328
rect 268672 662318 268700 664020
rect 279528 662318 279556 685850
rect 295812 683890 295840 685918
rect 305460 685908 305512 685914
rect 305460 685850 305512 685856
rect 305472 683890 305500 685850
rect 295734 683862 295840 683890
rect 305394 683862 305500 683890
rect 286074 683330 286180 683346
rect 285772 683324 285824 683330
rect 286074 683324 286192 683330
rect 286074 683318 286140 683324
rect 285772 683266 285824 683272
rect 286140 683266 286192 683272
rect 280160 683256 280212 683262
rect 280160 683198 280212 683204
rect 280172 673713 280200 683198
rect 284208 683188 284260 683194
rect 284208 683130 284260 683136
rect 284220 674801 284248 683130
rect 284206 674792 284262 674801
rect 284206 674727 284262 674736
rect 280158 673704 280214 673713
rect 280158 673639 280214 673648
rect 285784 662386 285812 683266
rect 305564 683114 305592 685918
rect 307024 685908 307076 685914
rect 307024 685850 307076 685856
rect 305472 683086 305592 683114
rect 305472 664714 305500 683086
rect 305394 664686 305500 664714
rect 285772 662380 285824 662386
rect 285772 662322 285824 662328
rect 268660 662312 268712 662318
rect 268660 662254 268712 662260
rect 279516 662312 279568 662318
rect 279516 662254 279568 662260
rect 286060 662250 286088 664020
rect 295720 662318 295748 664020
rect 307036 662318 307064 685850
rect 322400 683890 322428 685918
rect 331956 685908 332008 685914
rect 331956 685850 332008 685856
rect 333244 685908 333296 685914
rect 333244 685850 333296 685856
rect 331968 683890 331996 685850
rect 322400 683862 322690 683890
rect 331968 683862 332350 683890
rect 312004 683318 313030 683346
rect 311808 683256 311860 683262
rect 311808 683198 311860 683204
rect 311820 674393 311848 683198
rect 311806 674384 311862 674393
rect 311806 674319 311862 674328
rect 307758 673568 307814 673577
rect 307758 673503 307814 673512
rect 307772 665174 307800 673503
rect 307760 665168 307812 665174
rect 307760 665110 307812 665116
rect 295708 662312 295760 662318
rect 295708 662254 295760 662260
rect 307024 662312 307076 662318
rect 307024 662254 307076 662260
rect 312004 662250 312032 683318
rect 332508 665168 332560 665174
rect 332508 665110 332560 665116
rect 332520 664714 332548 665110
rect 332350 664686 332548 664714
rect 313016 662386 313044 664020
rect 313004 662380 313056 662386
rect 313004 662322 313056 662328
rect 322676 662318 322704 664020
rect 333256 662318 333284 685850
rect 334636 665174 334664 685918
rect 349816 683890 349844 685918
rect 359464 685908 359516 685914
rect 359464 685850 359516 685856
rect 359476 683890 359504 685850
rect 349738 683862 349844 683890
rect 359398 683862 359504 683890
rect 359660 683618 359688 685918
rect 359740 685908 359792 685914
rect 359740 685850 359792 685856
rect 359476 683590 359688 683618
rect 340078 683330 340184 683346
rect 339592 683324 339644 683330
rect 340078 683324 340196 683330
rect 340078 683318 340144 683324
rect 339592 683266 339644 683272
rect 340144 683266 340196 683272
rect 335360 683188 335412 683194
rect 335360 683130 335412 683136
rect 335372 673713 335400 683130
rect 338026 674248 338082 674257
rect 338026 674183 338082 674192
rect 335358 673704 335414 673713
rect 335358 673639 335414 673648
rect 338040 665174 338068 674183
rect 334624 665168 334676 665174
rect 334624 665110 334676 665116
rect 338028 665168 338080 665174
rect 338028 665110 338080 665116
rect 339604 662386 339632 683266
rect 359476 664714 359504 683590
rect 359752 683114 359780 685850
rect 376312 683890 376340 685918
rect 386052 685908 386104 685914
rect 386052 685850 386104 685856
rect 386064 683890 386092 685850
rect 376312 683862 376694 683890
rect 386064 683862 386354 683890
rect 365824 683318 367034 683346
rect 361580 683256 361632 683262
rect 361580 683198 361632 683204
rect 359398 664686 359504 664714
rect 359568 683086 359780 683114
rect 339592 662380 339644 662386
rect 339592 662322 339644 662328
rect 322664 662312 322716 662318
rect 322664 662254 322716 662260
rect 333244 662312 333296 662318
rect 333244 662254 333296 662260
rect 340064 662250 340092 664020
rect 349724 662318 349752 664020
rect 359568 662318 359596 683086
rect 361592 674257 361620 683198
rect 365628 683188 365680 683194
rect 365628 683130 365680 683136
rect 365640 674393 365668 683130
rect 365626 674384 365682 674393
rect 365626 674319 365682 674328
rect 361578 674248 361634 674257
rect 361578 674183 361634 674192
rect 365824 662318 365852 683318
rect 386524 664714 386552 685918
rect 387064 685908 387116 685914
rect 387064 685850 387116 685856
rect 386354 664686 386552 664714
rect 366744 664006 367034 664034
rect 366744 662386 366772 664006
rect 366732 662380 366784 662386
rect 366732 662322 366784 662328
rect 376680 662318 376708 664020
rect 387076 662318 387104 685850
rect 403360 683890 403388 685918
rect 412916 685908 412968 685914
rect 412916 685850 412968 685856
rect 412928 683890 412956 685850
rect 403360 683862 403650 683890
rect 412928 683862 413310 683890
rect 393424 683318 393990 683346
rect 391846 674248 391902 674257
rect 391846 674183 391902 674192
rect 389178 673568 389234 673577
rect 389178 673503 389234 673512
rect 389192 665174 389220 673503
rect 391860 665174 391888 674183
rect 389180 665168 389232 665174
rect 389180 665110 389232 665116
rect 391848 665168 391900 665174
rect 391848 665110 391900 665116
rect 393424 662318 393452 683318
rect 413480 664714 413508 685986
rect 421288 685976 421340 685982
rect 421288 685918 421340 685924
rect 414664 685908 414716 685914
rect 414664 685850 414716 685856
rect 413402 664686 413508 664714
rect 393608 664006 393990 664034
rect 393608 662386 393636 664006
rect 393596 662380 393648 662386
rect 393596 662322 393648 662328
rect 403728 662318 403756 664020
rect 414676 662318 414704 685850
rect 421300 683890 421328 685918
rect 421038 683862 421328 683890
rect 430592 683890 430620 685986
rect 440240 685908 440292 685914
rect 440240 685850 440292 685856
rect 440252 683890 440280 685850
rect 430592 683862 430698 683890
rect 440252 683862 440358 683890
rect 415400 683188 415452 683194
rect 415400 683130 415452 683136
rect 419448 683188 419500 683194
rect 419448 683130 419500 683136
rect 415412 673713 415440 683130
rect 419460 674393 419488 683130
rect 419446 674384 419502 674393
rect 419446 674319 419502 674328
rect 415398 673704 415454 673713
rect 415398 673639 415454 673648
rect 440528 664714 440556 685986
rect 443644 685976 443696 685982
rect 443644 685918 443696 685924
rect 442264 685908 442316 685914
rect 442264 685850 442316 685856
rect 440358 664686 440556 664714
rect 421024 662386 421052 664020
rect 430684 662386 430712 664020
rect 442276 662386 442304 685850
rect 442998 673568 443054 673577
rect 442998 673503 443054 673512
rect 443012 665174 443040 673503
rect 443000 665168 443052 665174
rect 443000 665110 443052 665116
rect 443656 662386 443684 685918
rect 457272 683890 457300 685986
rect 467012 685908 467064 685914
rect 467012 685850 467064 685856
rect 468484 685908 468536 685914
rect 468484 685850 468536 685856
rect 467024 683890 467052 685850
rect 457272 683862 457654 683890
rect 467024 683862 467314 683890
rect 447244 683318 447994 683346
rect 445666 674248 445722 674257
rect 445666 674183 445722 674192
rect 445680 665174 445708 674183
rect 445668 665168 445720 665174
rect 445668 665110 445720 665116
rect 421012 662380 421064 662386
rect 421012 662322 421064 662328
rect 430672 662380 430724 662386
rect 430672 662322 430724 662328
rect 442264 662380 442316 662386
rect 442264 662322 442316 662328
rect 443644 662380 443696 662386
rect 443644 662322 443696 662328
rect 349712 662312 349764 662318
rect 349712 662254 349764 662260
rect 359556 662312 359608 662318
rect 359556 662254 359608 662260
rect 365812 662312 365864 662318
rect 365812 662254 365864 662260
rect 376668 662312 376720 662318
rect 376668 662254 376720 662260
rect 387064 662312 387116 662318
rect 387064 662254 387116 662260
rect 393412 662312 393464 662318
rect 393412 662254 393464 662260
rect 403716 662312 403768 662318
rect 403716 662254 403768 662260
rect 414664 662312 414716 662318
rect 414664 662254 414716 662260
rect 447244 662250 447272 683318
rect 467656 665100 467708 665106
rect 467656 665042 467708 665048
rect 467668 664714 467696 665042
rect 467406 664686 467696 664714
rect 447704 664006 447994 664034
rect 447704 662386 447732 664006
rect 447692 662380 447744 662386
rect 447692 662322 447744 662328
rect 457732 662318 457760 664020
rect 468496 662318 468524 685850
rect 468588 665106 468616 685986
rect 475384 685976 475436 685982
rect 475384 685918 475436 685924
rect 475396 683890 475424 685918
rect 475042 683862 475424 683890
rect 484412 683890 484440 685986
rect 494060 685908 494112 685914
rect 494060 685850 494112 685856
rect 494072 683890 494100 685850
rect 484412 683862 484702 683890
rect 494072 683862 494362 683890
rect 469220 683188 469272 683194
rect 469220 683130 469272 683136
rect 473268 683188 473320 683194
rect 473268 683130 473320 683136
rect 469232 674257 469260 683130
rect 473280 674801 473308 683130
rect 473266 674792 473322 674801
rect 473266 674727 473322 674736
rect 469218 674248 469274 674257
rect 469218 674183 469274 674192
rect 468576 665100 468628 665106
rect 468576 665042 468628 665048
rect 494532 664714 494560 685986
rect 494704 685976 494756 685982
rect 494704 685918 494756 685924
rect 494362 664686 494560 664714
rect 457720 662312 457772 662318
rect 457720 662254 457772 662260
rect 468484 662312 468536 662318
rect 468484 662254 468536 662260
rect 475028 662250 475056 664020
rect 484688 662318 484716 664020
rect 494716 662386 494744 685918
rect 496084 685908 496136 685914
rect 496084 685850 496136 685856
rect 494704 662380 494756 662386
rect 494704 662322 494756 662328
rect 496096 662318 496124 685850
rect 511368 683890 511396 685986
rect 522396 685976 522448 685982
rect 522396 685918 522448 685924
rect 538404 685976 538456 685982
rect 538404 685918 538456 685924
rect 520924 685908 520976 685914
rect 520924 685850 520976 685856
rect 522304 685908 522356 685914
rect 522304 685850 522356 685856
rect 520936 683890 520964 685850
rect 511368 683862 511658 683890
rect 520936 683862 521318 683890
rect 501064 683318 501998 683346
rect 500868 683256 500920 683262
rect 500868 683198 500920 683204
rect 500880 674393 500908 683198
rect 500866 674384 500922 674393
rect 500866 674319 500922 674328
rect 496818 673568 496874 673577
rect 496818 673503 496874 673512
rect 496832 665174 496860 673503
rect 496820 665168 496872 665174
rect 496820 665110 496872 665116
rect 484676 662312 484728 662318
rect 484676 662254 484728 662260
rect 496084 662312 496136 662318
rect 496084 662254 496136 662260
rect 501064 662250 501092 683318
rect 501984 662386 502012 664020
rect 501972 662380 502024 662386
rect 501972 662322 502024 662328
rect 511736 662318 511764 664020
rect 521396 663746 521424 664020
rect 521384 663740 521436 663746
rect 521384 663682 521436 663688
rect 522316 662318 522344 685850
rect 522408 663746 522436 685918
rect 538416 683890 538444 685918
rect 548064 685908 548116 685914
rect 548064 685850 548116 685856
rect 548076 683890 548104 685850
rect 538416 683862 538706 683890
rect 548076 683862 548366 683890
rect 550640 683256 550692 683262
rect 550640 683198 550692 683204
rect 523040 683188 523092 683194
rect 523040 683130 523092 683136
rect 523052 673713 523080 683130
rect 527086 674248 527142 674257
rect 527086 674183 527142 674192
rect 523038 673704 523094 673713
rect 523038 673639 523094 673648
rect 522396 663740 522448 663746
rect 522396 663682 522448 663688
rect 511724 662312 511776 662318
rect 511724 662254 511776 662260
rect 522304 662312 522356 662318
rect 522304 662254 522356 662260
rect 150992 662244 151044 662250
rect 150992 662186 151044 662192
rect 258172 662244 258224 662250
rect 258172 662186 258224 662192
rect 286048 662244 286100 662250
rect 286048 662186 286100 662192
rect 311992 662244 312044 662250
rect 311992 662186 312044 662192
rect 340052 662244 340104 662250
rect 340052 662186 340104 662192
rect 447232 662244 447284 662250
rect 447232 662186 447284 662192
rect 475016 662244 475068 662250
rect 475016 662186 475068 662192
rect 501052 662244 501104 662250
rect 501052 662186 501104 662192
rect 232044 658504 232096 658510
rect 232044 658446 232096 658452
rect 251824 658504 251876 658510
rect 251824 658446 251876 658452
rect 475016 658504 475068 658510
rect 475016 658446 475068 658452
rect 494704 658504 494756 658510
rect 494704 658446 494756 658452
rect 170496 658436 170548 658442
rect 170496 658378 170548 658384
rect 187700 658436 187752 658442
rect 187700 658378 187752 658384
rect 197452 658436 197504 658442
rect 197452 658378 197504 658384
rect 214656 658436 214708 658442
rect 214656 658378 214708 658384
rect 224500 658436 224552 658442
rect 224500 658378 224552 658384
rect 170312 658368 170364 658374
rect 170312 658310 170364 658316
rect 160652 658300 160704 658306
rect 160652 658242 160704 658248
rect 160664 656948 160692 658242
rect 170324 656948 170352 658310
rect 150544 656254 151018 656282
rect 149704 634704 149756 634710
rect 149704 634646 149756 634652
rect 150544 634642 150572 656254
rect 150728 637078 151018 637106
rect 160572 637078 160678 637106
rect 170232 637078 170338 637106
rect 150532 634636 150584 634642
rect 150532 634578 150584 634584
rect 150728 634574 150756 637078
rect 160572 634574 160600 637078
rect 170232 636970 170260 637078
rect 170508 636970 170536 658378
rect 178040 658368 178092 658374
rect 178040 658310 178092 658316
rect 171784 658300 171836 658306
rect 171784 658242 171836 658248
rect 170232 636942 170536 636970
rect 171796 634574 171824 658242
rect 178052 656948 178080 658310
rect 187712 656948 187740 658378
rect 197360 658300 197412 658306
rect 197360 658242 197412 658248
rect 197372 656948 197400 658242
rect 172520 655648 172572 655654
rect 172520 655590 172572 655596
rect 176568 655648 176620 655654
rect 176568 655590 176620 655596
rect 172532 646649 172560 655590
rect 176580 647873 176608 655590
rect 176566 647864 176622 647873
rect 176566 647799 176622 647808
rect 172518 646640 172574 646649
rect 172518 646575 172574 646584
rect 197464 637786 197492 658378
rect 200764 658368 200816 658374
rect 200764 658310 200816 658316
rect 199384 658300 199436 658306
rect 199384 658242 199436 658248
rect 197386 637758 197492 637786
rect 178066 637078 178172 637106
rect 187726 637078 188016 637106
rect 178144 634642 178172 637078
rect 187988 634642 188016 637078
rect 199396 634642 199424 658242
rect 200120 655580 200172 655586
rect 200120 655522 200172 655528
rect 200132 646649 200160 655522
rect 200118 646640 200174 646649
rect 200118 646575 200174 646584
rect 200776 634778 200804 658310
rect 214668 656948 214696 658378
rect 224316 658300 224368 658306
rect 224316 658242 224368 658248
rect 224328 656948 224356 658242
rect 204364 656254 205022 656282
rect 202788 655580 202840 655586
rect 202788 655522 202840 655528
rect 202800 647329 202828 655522
rect 202786 647320 202842 647329
rect 202786 647255 202842 647264
rect 200764 634772 200816 634778
rect 200764 634714 200816 634720
rect 204364 634642 204392 656254
rect 224512 637786 224540 658378
rect 225604 658300 225656 658306
rect 225604 658242 225656 658248
rect 224342 637758 224540 637786
rect 204640 637078 205022 637106
rect 214682 637078 215064 637106
rect 204640 634778 204668 637078
rect 204628 634772 204680 634778
rect 204628 634714 204680 634720
rect 178132 634636 178184 634642
rect 178132 634578 178184 634584
rect 187976 634636 188028 634642
rect 187976 634578 188028 634584
rect 199384 634636 199436 634642
rect 199384 634578 199436 634584
rect 204352 634636 204404 634642
rect 204352 634578 204404 634584
rect 215036 634574 215064 637078
rect 225616 634574 225644 658242
rect 232056 656948 232084 658446
rect 241704 658436 241756 658442
rect 241704 658378 241756 658384
rect 241716 656948 241744 658378
rect 251456 658368 251508 658374
rect 251456 658310 251508 658316
rect 251364 658300 251416 658306
rect 251364 658242 251416 658248
rect 251376 656948 251404 658242
rect 226340 655648 226392 655654
rect 226340 655590 226392 655596
rect 230388 655648 230440 655654
rect 230388 655590 230440 655596
rect 226352 646649 226380 655590
rect 230400 647329 230428 655590
rect 230386 647320 230442 647329
rect 230386 647255 230442 647264
rect 226338 646640 226394 646649
rect 226338 646575 226394 646584
rect 251468 637786 251496 658310
rect 251390 637758 251496 637786
rect 231964 637078 232070 637106
rect 241730 637078 242112 637106
rect 231964 634642 231992 637078
rect 242084 634642 242112 637078
rect 251836 634778 251864 658446
rect 413468 658436 413520 658442
rect 413468 658378 413520 658384
rect 430672 658436 430724 658442
rect 430672 658378 430724 658384
rect 440516 658436 440568 658442
rect 440516 658378 440568 658384
rect 457628 658436 457680 658442
rect 457628 658378 457680 658384
rect 468484 658436 468536 658442
rect 468484 658378 468536 658384
rect 268660 658368 268712 658374
rect 268660 658310 268712 658316
rect 279424 658368 279476 658374
rect 279424 658310 279476 658316
rect 295708 658368 295760 658374
rect 295708 658310 295760 658316
rect 305460 658368 305512 658374
rect 305460 658310 305512 658316
rect 322664 658368 322716 658374
rect 322664 658310 322716 658316
rect 336004 658368 336056 658374
rect 336004 658310 336056 658316
rect 349712 658368 349764 658374
rect 349712 658310 349764 658316
rect 359464 658368 359516 658374
rect 359464 658310 359516 658316
rect 376668 658368 376720 658374
rect 376668 658310 376720 658316
rect 386512 658368 386564 658374
rect 386512 658310 386564 658316
rect 403624 658368 403676 658374
rect 403624 658310 403676 658316
rect 253204 658300 253256 658306
rect 253204 658242 253256 658248
rect 251824 634772 251876 634778
rect 251824 634714 251876 634720
rect 253216 634642 253244 658242
rect 268672 656948 268700 658310
rect 278320 658300 278372 658306
rect 278320 658242 278372 658248
rect 278332 656948 278360 658242
rect 258184 656254 259026 656282
rect 253940 655580 253992 655586
rect 253940 655522 253992 655528
rect 256608 655580 256660 655586
rect 256608 655522 256660 655528
rect 253952 647193 253980 655522
rect 256620 647329 256648 655522
rect 256606 647320 256662 647329
rect 256606 647255 256662 647264
rect 253938 647184 253994 647193
rect 253938 647119 253994 647128
rect 258184 634642 258212 656254
rect 279436 644474 279464 658310
rect 279516 658300 279568 658306
rect 279516 658242 279568 658248
rect 278792 644446 279464 644474
rect 278792 637514 278820 644446
rect 278346 637486 278820 637514
rect 258736 637078 259026 637106
rect 268686 637078 268976 637106
rect 258736 634778 258764 637078
rect 258724 634772 258776 634778
rect 258724 634714 258776 634720
rect 231952 634636 232004 634642
rect 231952 634578 232004 634584
rect 242072 634636 242124 634642
rect 242072 634578 242124 634584
rect 253204 634636 253256 634642
rect 253204 634578 253256 634584
rect 258172 634636 258224 634642
rect 258172 634578 258224 634584
rect 268948 634574 268976 637078
rect 279528 634574 279556 658242
rect 285784 657070 286088 657098
rect 280160 655648 280212 655654
rect 280160 655590 280212 655596
rect 284208 655648 284260 655654
rect 284208 655590 284260 655596
rect 280172 646649 280200 655590
rect 284220 647873 284248 655590
rect 284206 647864 284262 647873
rect 284206 647799 284262 647808
rect 280158 646640 280214 646649
rect 280158 646575 280214 646584
rect 285784 634642 285812 657070
rect 286060 656948 286088 657070
rect 295720 656948 295748 658310
rect 305368 658300 305420 658306
rect 305368 658242 305420 658248
rect 305380 656948 305408 658242
rect 305472 637786 305500 658310
rect 307024 658300 307076 658306
rect 307024 658242 307076 658248
rect 305394 637758 305500 637786
rect 286074 637078 286180 637106
rect 295734 637078 296024 637106
rect 285772 634636 285824 634642
rect 285772 634578 285824 634584
rect 286152 634574 286180 637078
rect 295996 634574 296024 637078
rect 307036 634574 307064 658242
rect 322676 656948 322704 658310
rect 332324 658300 332376 658306
rect 332324 658242 332376 658248
rect 333244 658300 333296 658306
rect 333244 658242 333296 658248
rect 332336 656948 332364 658242
rect 312004 656254 313030 656282
rect 311808 655716 311860 655722
rect 311808 655658 311860 655664
rect 307760 655580 307812 655586
rect 307760 655522 307812 655528
rect 307772 646649 307800 655522
rect 311820 647329 311848 655658
rect 311806 647320 311862 647329
rect 311806 647255 311862 647264
rect 307758 646640 307814 646649
rect 307758 646575 307814 646584
rect 312004 634574 312032 656254
rect 332600 637560 332652 637566
rect 332350 637508 332600 637514
rect 332350 637502 332652 637508
rect 332350 637486 332640 637502
rect 312648 637078 313030 637106
rect 322690 637078 322888 637106
rect 312648 634642 312676 637078
rect 312636 634636 312688 634642
rect 312636 634578 312688 634584
rect 322860 634574 322888 637078
rect 333256 634574 333284 658242
rect 335360 655648 335412 655654
rect 335360 655590 335412 655596
rect 335372 646649 335400 655590
rect 335358 646640 335414 646649
rect 335358 646575 335414 646584
rect 336016 637566 336044 658310
rect 339604 657070 340092 657098
rect 338028 655580 338080 655586
rect 338028 655522 338080 655528
rect 338040 647329 338068 655522
rect 338026 647320 338082 647329
rect 338026 647255 338082 647264
rect 336004 637560 336056 637566
rect 336004 637502 336056 637508
rect 339604 634574 339632 657070
rect 340064 656948 340092 657070
rect 349724 656948 349752 658310
rect 359372 658300 359424 658306
rect 359372 658242 359424 658248
rect 359384 656948 359412 658242
rect 359476 637786 359504 658310
rect 359556 658300 359608 658306
rect 359556 658242 359608 658248
rect 359398 637758 359504 637786
rect 340078 637078 340184 637106
rect 349738 637078 350120 637106
rect 340156 634642 340184 637078
rect 340144 634636 340196 634642
rect 340144 634578 340196 634584
rect 350092 634574 350120 637078
rect 359568 634574 359596 658242
rect 376680 656948 376708 658310
rect 386328 658300 386380 658306
rect 386328 658242 386380 658248
rect 386340 656948 386368 658242
rect 365824 656254 367034 656282
rect 361580 655716 361632 655722
rect 361580 655658 361632 655664
rect 361592 647193 361620 655658
rect 365628 655648 365680 655654
rect 365628 655590 365680 655596
rect 365640 647329 365668 655590
rect 365626 647320 365682 647329
rect 365626 647255 365682 647264
rect 361578 647184 361634 647193
rect 361578 647119 361634 647128
rect 365824 634574 365852 656254
rect 386524 637786 386552 658310
rect 387064 658300 387116 658306
rect 387064 658242 387116 658248
rect 386354 637758 386552 637786
rect 366744 637078 367034 637106
rect 376588 637078 376694 637106
rect 366744 634642 366772 637078
rect 366732 634636 366784 634642
rect 366732 634578 366784 634584
rect 376588 634574 376616 637078
rect 387076 634574 387104 658242
rect 403636 656948 403664 658310
rect 413284 658300 413336 658306
rect 413284 658242 413336 658248
rect 413296 656948 413324 658242
rect 393424 656254 393990 656282
rect 389180 655580 389232 655586
rect 389180 655522 389232 655528
rect 391848 655580 391900 655586
rect 391848 655522 391900 655528
rect 389192 646649 389220 655522
rect 391860 647329 391888 655522
rect 391846 647320 391902 647329
rect 391846 647255 391902 647264
rect 389178 646640 389234 646649
rect 389178 646575 389234 646584
rect 393424 634574 393452 656254
rect 413480 637786 413508 658378
rect 421012 658368 421064 658374
rect 421012 658310 421064 658316
rect 414664 658300 414716 658306
rect 414664 658242 414716 658248
rect 413402 637758 413508 637786
rect 393608 637078 393990 637106
rect 403742 637078 404032 637106
rect 393608 634642 393636 637078
rect 393596 634636 393648 634642
rect 393596 634578 393648 634584
rect 404004 634574 404032 637078
rect 414676 634574 414704 658242
rect 421024 656948 421052 658310
rect 430684 656948 430712 658378
rect 440332 658300 440384 658306
rect 440332 658242 440384 658248
rect 440344 656948 440372 658242
rect 415400 655648 415452 655654
rect 415400 655590 415452 655596
rect 419448 655648 419500 655654
rect 419448 655590 419500 655596
rect 415412 646649 415440 655590
rect 419460 647329 419488 655590
rect 419446 647320 419502 647329
rect 419446 647255 419502 647264
rect 415398 646640 415454 646649
rect 415398 646575 415454 646584
rect 440528 637786 440556 658378
rect 446404 658368 446456 658374
rect 446404 658310 446456 658316
rect 442264 658300 442316 658306
rect 442264 658242 442316 658248
rect 440358 637758 440556 637786
rect 420932 637078 421038 637106
rect 430698 637078 431080 637106
rect 420932 634642 420960 637078
rect 431052 634642 431080 637078
rect 442276 634642 442304 658242
rect 443000 655580 443052 655586
rect 443000 655522 443052 655528
rect 445668 655580 445720 655586
rect 445668 655522 445720 655528
rect 443012 646649 443040 655522
rect 445680 647329 445708 655522
rect 445666 647320 445722 647329
rect 445666 647255 445722 647264
rect 442998 646640 443054 646649
rect 442998 646575 443054 646584
rect 446416 637566 446444 658310
rect 457640 656948 457668 658378
rect 467288 658300 467340 658306
rect 467288 658242 467340 658248
rect 467300 656948 467328 658242
rect 447244 656254 447994 656282
rect 446404 637560 446456 637566
rect 446404 637502 446456 637508
rect 447244 634642 447272 656254
rect 468496 644474 468524 658378
rect 468576 658300 468628 658306
rect 468576 658242 468628 658248
rect 467852 644446 468524 644474
rect 447692 637560 447744 637566
rect 467852 637514 467880 644446
rect 447744 637508 447994 637514
rect 447692 637502 447994 637508
rect 447704 637486 447994 637502
rect 467406 637486 467880 637514
rect 457746 637078 458128 637106
rect 420920 634636 420972 634642
rect 420920 634578 420972 634584
rect 431040 634636 431092 634642
rect 431040 634578 431092 634584
rect 442264 634636 442316 634642
rect 442264 634578 442316 634584
rect 447232 634636 447284 634642
rect 447232 634578 447284 634584
rect 458100 634574 458128 637078
rect 468588 634574 468616 658242
rect 475028 656948 475056 658446
rect 484676 658436 484728 658442
rect 484676 658378 484728 658384
rect 484688 656948 484716 658378
rect 494520 658368 494572 658374
rect 494520 658310 494572 658316
rect 494336 658300 494388 658306
rect 494336 658242 494388 658248
rect 494348 656948 494376 658242
rect 469220 655648 469272 655654
rect 469220 655590 469272 655596
rect 473268 655648 473320 655654
rect 473268 655590 473320 655596
rect 469232 647193 469260 655590
rect 473280 647873 473308 655590
rect 473266 647864 473322 647873
rect 473266 647799 473322 647808
rect 469218 647184 469274 647193
rect 469218 647119 469274 647128
rect 494532 637786 494560 658310
rect 494362 637758 494560 637786
rect 474752 637078 475042 637106
rect 484702 637078 484992 637106
rect 474752 634642 474780 637078
rect 484964 634642 484992 637078
rect 494716 634778 494744 658446
rect 511632 658368 511684 658374
rect 511632 658310 511684 658316
rect 522304 658368 522356 658374
rect 522304 658310 522356 658316
rect 496084 658300 496136 658306
rect 496084 658242 496136 658248
rect 494704 634772 494756 634778
rect 494704 634714 494756 634720
rect 496096 634642 496124 658242
rect 511644 656948 511672 658310
rect 521292 658300 521344 658306
rect 521292 658242 521344 658248
rect 521304 656948 521332 658242
rect 501064 656254 501998 656282
rect 496820 655580 496872 655586
rect 496820 655522 496872 655528
rect 500868 655580 500920 655586
rect 500868 655522 500920 655528
rect 496832 646649 496860 655522
rect 500880 647329 500908 655522
rect 500866 647320 500922 647329
rect 500866 647255 500922 647264
rect 496818 646640 496874 646649
rect 496818 646575 496874 646584
rect 501064 634642 501092 656254
rect 501616 637078 501998 637106
rect 511750 637078 511856 637106
rect 521410 637078 521516 637106
rect 501616 634778 501644 637078
rect 501604 634772 501656 634778
rect 501604 634714 501656 634720
rect 474740 634636 474792 634642
rect 474740 634578 474792 634584
rect 484952 634636 485004 634642
rect 484952 634578 485004 634584
rect 496084 634636 496136 634642
rect 496084 634578 496136 634584
rect 501052 634636 501104 634642
rect 501052 634578 501104 634584
rect 511828 634574 511856 637078
rect 521488 634778 521516 637078
rect 522316 634778 522344 658310
rect 522396 658300 522448 658306
rect 522396 658242 522448 658248
rect 521476 634772 521528 634778
rect 521476 634714 521528 634720
rect 522304 634772 522356 634778
rect 522304 634714 522356 634720
rect 522408 634574 522436 658242
rect 526444 657552 526496 657558
rect 526444 657494 526496 657500
rect 523040 655648 523092 655654
rect 523040 655590 523092 655596
rect 523052 646649 523080 655590
rect 526456 647329 526484 657494
rect 526442 647320 526498 647329
rect 526442 647255 526498 647264
rect 523038 646640 523094 646649
rect 523038 646575 523094 646584
rect 150716 634568 150768 634574
rect 150716 634510 150768 634516
rect 160560 634568 160612 634574
rect 160560 634510 160612 634516
rect 171784 634568 171836 634574
rect 171784 634510 171836 634516
rect 215024 634568 215076 634574
rect 215024 634510 215076 634516
rect 225604 634568 225656 634574
rect 225604 634510 225656 634516
rect 268936 634568 268988 634574
rect 268936 634510 268988 634516
rect 279516 634568 279568 634574
rect 279516 634510 279568 634516
rect 286140 634568 286192 634574
rect 286140 634510 286192 634516
rect 295984 634568 296036 634574
rect 295984 634510 296036 634516
rect 307024 634568 307076 634574
rect 307024 634510 307076 634516
rect 311992 634568 312044 634574
rect 311992 634510 312044 634516
rect 322848 634568 322900 634574
rect 322848 634510 322900 634516
rect 333244 634568 333296 634574
rect 333244 634510 333296 634516
rect 339592 634568 339644 634574
rect 339592 634510 339644 634516
rect 350080 634568 350132 634574
rect 350080 634510 350132 634516
rect 359556 634568 359608 634574
rect 359556 634510 359608 634516
rect 365812 634568 365864 634574
rect 365812 634510 365864 634516
rect 376576 634568 376628 634574
rect 376576 634510 376628 634516
rect 387064 634568 387116 634574
rect 387064 634510 387116 634516
rect 393412 634568 393464 634574
rect 393412 634510 393464 634516
rect 403992 634568 404044 634574
rect 403992 634510 404044 634516
rect 414664 634568 414716 634574
rect 414664 634510 414716 634516
rect 458088 634568 458140 634574
rect 458088 634510 458140 634516
rect 468576 634568 468628 634574
rect 468576 634510 468628 634516
rect 511816 634568 511868 634574
rect 511816 634510 511868 634516
rect 522396 634568 522448 634574
rect 522396 634510 522448 634516
rect 148324 632392 148376 632398
rect 148324 632334 148376 632340
rect 146944 608592 146996 608598
rect 146944 608534 146996 608540
rect 124036 608524 124088 608530
rect 124036 608466 124088 608472
rect 133696 608524 133748 608530
rect 133696 608466 133748 608472
rect 144276 608524 144328 608530
rect 144276 608466 144328 608472
rect 79692 608456 79744 608462
rect 79692 608398 79744 608404
rect 90456 608456 90508 608462
rect 90456 608398 90508 608404
rect 106648 608456 106700 608462
rect 106648 608398 106700 608404
rect 116584 608456 116636 608462
rect 116584 608398 116636 608404
rect 122932 608456 122984 608462
rect 122932 608398 122984 608404
rect 146944 604784 146996 604790
rect 146944 604726 146996 604732
rect 52644 604716 52696 604722
rect 52644 604658 52696 604664
rect 43076 604512 43128 604518
rect 43076 604454 43128 604460
rect 43088 602956 43116 604454
rect 52656 602956 52684 604658
rect 62488 604648 62540 604654
rect 62488 604590 62540 604596
rect 79692 604648 79744 604654
rect 79692 604590 79744 604596
rect 90456 604648 90508 604654
rect 90456 604590 90508 604596
rect 106648 604648 106700 604654
rect 106648 604590 106700 604596
rect 116492 604648 116544 604654
rect 116492 604590 116544 604596
rect 133696 604648 133748 604654
rect 133696 604590 133748 604596
rect 62304 604580 62356 604586
rect 62304 604522 62356 604528
rect 62316 602956 62344 604522
rect 37924 602404 37976 602410
rect 37924 602346 37976 602352
rect 41326 593192 41382 593201
rect 41326 593127 41382 593136
rect 37922 592104 37978 592113
rect 37922 592039 37978 592048
rect 36820 580848 36872 580854
rect 36820 580790 36872 580796
rect 36728 578468 36780 578474
rect 36728 578410 36780 578416
rect 36740 557462 36768 578410
rect 36820 578332 36872 578338
rect 36820 578274 36872 578280
rect 36728 557456 36780 557462
rect 36728 557398 36780 557404
rect 36832 554606 36860 578274
rect 37936 576162 37964 592039
rect 41340 583642 41368 593127
rect 62500 583794 62528 604590
rect 64144 604580 64196 604586
rect 64144 604522 64196 604528
rect 62764 604512 62816 604518
rect 62764 604454 62816 604460
rect 62422 583766 62528 583794
rect 41328 583636 41380 583642
rect 41328 583578 41380 583584
rect 42812 583086 43010 583114
rect 52762 583086 53144 583114
rect 42812 580922 42840 583086
rect 53116 580922 53144 583086
rect 62776 580990 62804 604454
rect 62764 580984 62816 580990
rect 62764 580926 62816 580932
rect 64156 580922 64184 604522
rect 79704 602956 79732 604590
rect 89352 604580 89404 604586
rect 89352 604522 89404 604528
rect 90364 604580 90416 604586
rect 90364 604522 90416 604528
rect 89364 602956 89392 604522
rect 69124 602262 70058 602290
rect 68926 592648 68982 592657
rect 68926 592583 68982 592592
rect 64878 592512 64934 592521
rect 64878 592447 64934 592456
rect 64892 583710 64920 592447
rect 64880 583704 64932 583710
rect 64880 583646 64932 583652
rect 68940 583574 68968 592583
rect 68928 583568 68980 583574
rect 68928 583510 68980 583516
rect 69124 580922 69152 602262
rect 89720 583704 89772 583710
rect 89378 583652 89720 583658
rect 89378 583646 89772 583652
rect 89378 583630 89760 583646
rect 69768 583086 70058 583114
rect 79718 583086 80008 583114
rect 69768 580990 69796 583086
rect 69756 580984 69808 580990
rect 69756 580926 69808 580932
rect 42800 580916 42852 580922
rect 42800 580858 42852 580864
rect 53104 580916 53156 580922
rect 53104 580858 53156 580864
rect 64144 580916 64196 580922
rect 64144 580858 64196 580864
rect 69112 580916 69164 580922
rect 69112 580858 69164 580864
rect 79980 580854 80008 583086
rect 90376 580854 90404 604522
rect 90468 583710 90496 604590
rect 106660 602956 106688 604590
rect 116308 604580 116360 604586
rect 116308 604522 116360 604528
rect 116320 602956 116348 604522
rect 96724 602262 97014 602290
rect 95146 593192 95202 593201
rect 95146 593127 95202 593136
rect 91098 592512 91154 592521
rect 91098 592447 91154 592456
rect 90456 583704 90508 583710
rect 90456 583646 90508 583652
rect 91112 583642 91140 592447
rect 95160 583710 95188 593127
rect 95148 583704 95200 583710
rect 95148 583646 95200 583652
rect 91100 583636 91152 583642
rect 91100 583578 91152 583584
rect 96724 580990 96752 602262
rect 116228 583642 116334 583658
rect 116504 583642 116532 604590
rect 116584 604580 116636 604586
rect 116584 604522 116636 604528
rect 116216 583636 116334 583642
rect 116268 583630 116334 583636
rect 116492 583636 116544 583642
rect 116216 583578 116268 583584
rect 116492 583578 116544 583584
rect 96816 583086 97014 583114
rect 106568 583086 106674 583114
rect 96712 580984 96764 580990
rect 96712 580926 96764 580932
rect 96816 580922 96844 583086
rect 96804 580916 96856 580922
rect 96804 580858 96856 580864
rect 106568 580854 106596 583086
rect 116596 580854 116624 604522
rect 133708 602956 133736 604590
rect 143356 604580 143408 604586
rect 143356 604522 143408 604528
rect 144276 604580 144328 604586
rect 144276 604522 144328 604528
rect 143368 602956 143396 604522
rect 144184 604512 144236 604518
rect 144184 604454 144236 604460
rect 122944 602262 124062 602290
rect 122746 593192 122802 593201
rect 122746 593127 122802 593136
rect 118698 592512 118754 592521
rect 118698 592447 118754 592456
rect 118712 583574 118740 592447
rect 122760 583642 122788 593127
rect 122748 583636 122800 583642
rect 122748 583578 122800 583584
rect 118700 583568 118752 583574
rect 118700 583510 118752 583516
rect 79968 580848 80020 580854
rect 79968 580790 80020 580796
rect 90364 580848 90416 580854
rect 90364 580790 90416 580796
rect 106556 580848 106608 580854
rect 106556 580790 106608 580796
rect 116584 580848 116636 580854
rect 116584 580790 116636 580796
rect 122944 580786 122972 602262
rect 144196 586514 144224 604454
rect 143736 586486 144224 586514
rect 143736 583658 143764 586486
rect 143382 583630 143764 583658
rect 123680 583086 124062 583114
rect 133722 583086 133828 583114
rect 123680 580922 123708 583086
rect 123668 580916 123720 580922
rect 123668 580858 123720 580864
rect 133800 580854 133828 583086
rect 144288 580854 144316 604522
rect 146298 592104 146354 592113
rect 146298 592039 146354 592048
rect 146312 583710 146340 592039
rect 146300 583704 146352 583710
rect 146300 583646 146352 583652
rect 133788 580848 133840 580854
rect 133788 580790 133840 580796
rect 144276 580848 144328 580854
rect 144276 580790 144328 580796
rect 122932 580780 122984 580786
rect 122932 580722 122984 580728
rect 52460 578468 52512 578474
rect 52460 578410 52512 578416
rect 43352 578264 43404 578270
rect 43352 578206 43404 578212
rect 37924 576156 37976 576162
rect 37924 576098 37976 576104
rect 43364 575906 43392 578206
rect 43102 575878 43392 575906
rect 52472 575906 52500 578410
rect 62488 578400 62540 578406
rect 62488 578342 62540 578348
rect 79324 578400 79376 578406
rect 79324 578342 79376 578348
rect 90456 578400 90508 578406
rect 90456 578342 90508 578348
rect 106464 578400 106516 578406
rect 106464 578342 106516 578348
rect 116492 578400 116544 578406
rect 116492 578342 116544 578348
rect 133420 578400 133472 578406
rect 133420 578342 133472 578348
rect 144184 578400 144236 578406
rect 144184 578342 144236 578348
rect 62120 578332 62172 578338
rect 62120 578274 62172 578280
rect 62132 575906 62160 578274
rect 52472 575878 52670 575906
rect 62132 575878 62330 575906
rect 41326 566264 41382 566273
rect 41326 566199 41382 566208
rect 37922 565040 37978 565049
rect 37922 564975 37978 564984
rect 36820 554600 36872 554606
rect 36820 554542 36872 554548
rect 36636 554464 36688 554470
rect 36636 554406 36688 554412
rect 36636 550860 36688 550866
rect 36636 550802 36688 550808
rect 36648 529854 36676 550802
rect 36820 550724 36872 550730
rect 36820 550666 36872 550672
rect 36728 547936 36780 547942
rect 36728 547878 36780 547884
rect 36636 529848 36688 529854
rect 36636 529790 36688 529796
rect 36544 526856 36596 526862
rect 36544 526798 36596 526804
rect 16304 523728 16356 523734
rect 16304 523670 16356 523676
rect 25964 523320 26016 523326
rect 25964 523262 26016 523268
rect 25976 521914 26004 523262
rect 36544 523116 36596 523122
rect 36544 523058 36596 523064
rect 25714 521886 26004 521914
rect 35374 521762 35664 521778
rect 35374 521756 35676 521762
rect 35374 521750 35624 521756
rect 35624 521698 35676 521704
rect 15212 521206 16054 521234
rect 13728 520328 13780 520334
rect 13728 520270 13780 520276
rect 13740 512417 13768 520270
rect 13726 512408 13782 512417
rect 13726 512343 13782 512352
rect 15212 500886 15240 521206
rect 35374 502314 35664 502330
rect 35374 502308 35676 502314
rect 35374 502302 35624 502308
rect 35624 502250 35676 502256
rect 15200 500880 15252 500886
rect 15200 500822 15252 500828
rect 16040 497486 16068 502044
rect 25700 500818 25728 502044
rect 36556 500818 36584 523058
rect 36636 521756 36688 521762
rect 36636 521698 36688 521704
rect 25688 500812 25740 500818
rect 25688 500754 25740 500760
rect 36544 500812 36596 500818
rect 36544 500754 36596 500760
rect 16028 497480 16080 497486
rect 16028 497422 16080 497428
rect 25688 497140 25740 497146
rect 25688 497082 25740 497088
rect 25700 494972 25728 497082
rect 15212 494278 16054 494306
rect 35374 494278 36032 494306
rect 13726 485208 13782 485217
rect 13726 485143 13782 485152
rect 13740 476066 13768 485143
rect 13728 476060 13780 476066
rect 13728 476002 13780 476008
rect 15212 473278 15240 494278
rect 36004 489914 36032 494278
rect 36004 489886 36584 489914
rect 35624 475992 35676 475998
rect 35624 475934 35676 475940
rect 35636 475674 35664 475934
rect 35374 475646 35664 475674
rect 15304 475102 16054 475130
rect 25714 475102 26096 475130
rect 15200 473272 15252 473278
rect 15200 473214 15252 473220
rect 15304 469878 15332 475102
rect 26068 473210 26096 475102
rect 26056 473204 26108 473210
rect 26056 473146 26108 473152
rect 15292 469872 15344 469878
rect 15292 469814 15344 469820
rect 25964 469532 26016 469538
rect 25964 469474 26016 469480
rect 25976 467922 26004 469474
rect 35716 469464 35768 469470
rect 35716 469406 35768 469412
rect 25714 467894 26004 467922
rect 15212 467214 16054 467242
rect 35374 467214 35664 467242
rect 13728 466472 13780 466478
rect 13728 466414 13780 466420
rect 13740 458425 13768 466414
rect 13726 458416 13782 458425
rect 13726 458351 13782 458360
rect 15212 445670 15240 467214
rect 35636 466546 35664 467214
rect 35624 466540 35676 466546
rect 35624 466482 35676 466488
rect 35728 451274 35756 469406
rect 35452 451246 35756 451274
rect 35452 448746 35480 451246
rect 35374 448718 35480 448746
rect 15200 445664 15252 445670
rect 15200 445606 15252 445612
rect 16040 443698 16068 448052
rect 25700 445738 25728 448052
rect 25688 445732 25740 445738
rect 25688 445674 25740 445680
rect 36556 445466 36584 489886
rect 36648 473074 36676 521698
rect 36740 500682 36768 547878
rect 36832 526998 36860 550666
rect 37936 548554 37964 564975
rect 41340 557462 41368 566199
rect 41328 557456 41380 557462
rect 41328 557398 41380 557404
rect 62500 556730 62528 578342
rect 64144 578332 64196 578338
rect 64144 578274 64196 578280
rect 62764 578264 62816 578270
rect 62764 578206 62816 578212
rect 62422 556702 62528 556730
rect 42996 554674 43024 556036
rect 52748 554742 52776 556036
rect 52736 554736 52788 554742
rect 52736 554678 52788 554684
rect 62776 554674 62804 578206
rect 64156 554742 64184 578274
rect 79336 575906 79364 578342
rect 89076 578332 89128 578338
rect 89076 578274 89128 578280
rect 90364 578332 90416 578338
rect 90364 578274 90416 578280
rect 89088 575906 89116 578274
rect 79336 575878 79718 575906
rect 89088 575878 89378 575906
rect 69124 575334 70058 575362
rect 68926 565856 68982 565865
rect 68926 565791 68982 565800
rect 64878 565584 64934 565593
rect 64878 565519 64934 565528
rect 64892 557530 64920 565519
rect 64880 557524 64932 557530
rect 64880 557466 64932 557472
rect 68940 557394 68968 565791
rect 68928 557388 68980 557394
rect 68928 557330 68980 557336
rect 69124 554742 69152 575334
rect 89720 562352 89772 562358
rect 89720 562294 89772 562300
rect 89732 556730 89760 562294
rect 89378 556702 89760 556730
rect 64144 554736 64196 554742
rect 64144 554678 64196 554684
rect 69112 554736 69164 554742
rect 69112 554678 69164 554684
rect 70044 554674 70072 556036
rect 42984 554668 43036 554674
rect 42984 554610 43036 554616
rect 62764 554668 62816 554674
rect 62764 554610 62816 554616
rect 70032 554668 70084 554674
rect 70032 554610 70084 554616
rect 79704 554606 79732 556036
rect 90376 554606 90404 578274
rect 90468 562358 90496 578342
rect 106476 575906 106504 578342
rect 116124 578332 116176 578338
rect 116124 578274 116176 578280
rect 116136 575906 116164 578274
rect 106476 575878 106674 575906
rect 116136 575878 116334 575906
rect 96724 575334 97014 575362
rect 95146 566264 95202 566273
rect 95146 566199 95202 566208
rect 91098 565584 91154 565593
rect 91098 565519 91154 565528
rect 90456 562352 90508 562358
rect 90456 562294 90508 562300
rect 91112 557462 91140 565519
rect 95160 557530 95188 566199
rect 95148 557524 95200 557530
rect 95148 557466 95200 557472
rect 91100 557456 91152 557462
rect 91100 557398 91152 557404
rect 96724 554742 96752 575334
rect 96712 554736 96764 554742
rect 96712 554678 96764 554684
rect 97000 554674 97028 556036
rect 96988 554668 97040 554674
rect 96988 554610 97040 554616
rect 106660 554606 106688 556036
rect 116320 555914 116348 556036
rect 116504 555914 116532 578342
rect 116584 578332 116636 578338
rect 116584 578274 116636 578280
rect 116320 555886 116532 555914
rect 116596 554606 116624 578274
rect 133432 575906 133460 578342
rect 142988 578332 143040 578338
rect 142988 578274 143040 578280
rect 143000 575906 143028 578274
rect 133432 575878 133722 575906
rect 143000 575878 143382 575906
rect 122944 575334 124062 575362
rect 122746 566264 122802 566273
rect 122746 566199 122802 566208
rect 118698 565584 118754 565593
rect 118698 565519 118754 565528
rect 118712 557394 118740 565519
rect 122760 557462 122788 566199
rect 122748 557456 122800 557462
rect 122748 557398 122800 557404
rect 118700 557388 118752 557394
rect 118700 557330 118752 557336
rect 122944 554606 122972 575334
rect 144196 557534 144224 578342
rect 144276 578332 144328 578338
rect 144276 578274 144328 578280
rect 143736 557506 144224 557534
rect 143736 556730 143764 557506
rect 143382 556702 143764 556730
rect 124048 554674 124076 556036
rect 133708 554674 133736 556036
rect 144288 554674 144316 578274
rect 146298 565040 146354 565049
rect 146298 564975 146354 564984
rect 146312 557530 146340 564975
rect 146300 557524 146352 557530
rect 146300 557466 146352 557472
rect 146956 554742 146984 604726
rect 148336 580922 148364 632334
rect 232320 632324 232372 632330
rect 232320 632266 232372 632272
rect 251824 632324 251876 632330
rect 251824 632266 251876 632272
rect 475384 632324 475436 632330
rect 475384 632266 475436 632272
rect 494704 632324 494756 632330
rect 494704 632266 494756 632272
rect 170496 632256 170548 632262
rect 170496 632198 170548 632204
rect 187792 632256 187844 632262
rect 187792 632198 187844 632204
rect 197544 632256 197596 632262
rect 197544 632198 197596 632204
rect 214380 632256 214432 632262
rect 214380 632198 214432 632204
rect 224500 632256 224552 632262
rect 224500 632198 224552 632204
rect 170036 632188 170088 632194
rect 170036 632130 170088 632136
rect 160284 632120 160336 632126
rect 160284 632062 160336 632068
rect 160296 629898 160324 632062
rect 170048 629898 170076 632130
rect 160296 629870 160678 629898
rect 170048 629870 170338 629898
rect 150544 629326 151018 629354
rect 148966 620256 149022 620265
rect 148966 620191 149022 620200
rect 148980 611318 149008 620191
rect 148968 611312 149020 611318
rect 148968 611254 149020 611260
rect 150544 608530 150572 629326
rect 150532 608524 150584 608530
rect 150532 608466 150584 608472
rect 151004 608462 151032 610028
rect 150992 608456 151044 608462
rect 150992 608398 151044 608404
rect 160664 608394 160692 610028
rect 170324 609906 170352 610028
rect 170508 609906 170536 632198
rect 178408 632188 178460 632194
rect 178408 632130 178460 632136
rect 171784 632120 171836 632126
rect 171784 632062 171836 632068
rect 170324 609878 170536 609906
rect 171796 608394 171824 632062
rect 178420 629898 178448 632130
rect 187804 629898 187832 632198
rect 197452 632120 197504 632126
rect 197452 632062 197504 632068
rect 197464 629898 197492 632062
rect 178066 629870 178448 629898
rect 187726 629870 187832 629898
rect 197386 629870 197492 629898
rect 197556 625154 197584 632198
rect 200764 632188 200816 632194
rect 200764 632130 200816 632136
rect 199384 632120 199436 632126
rect 199384 632062 199436 632068
rect 197464 625126 197584 625154
rect 176566 619712 176622 619721
rect 176566 619647 176622 619656
rect 172518 619576 172574 619585
rect 172518 619511 172574 619520
rect 172532 611250 172560 619511
rect 176580 611250 176608 619647
rect 172520 611244 172572 611250
rect 172520 611186 172572 611192
rect 176568 611244 176620 611250
rect 176568 611186 176620 611192
rect 197464 610722 197492 625126
rect 197386 610694 197492 610722
rect 178052 608462 178080 610028
rect 187712 608462 187740 610028
rect 199396 608462 199424 632062
rect 200118 619576 200174 619585
rect 200118 619511 200174 619520
rect 200132 611318 200160 619511
rect 200120 611312 200172 611318
rect 200120 611254 200172 611260
rect 200776 608598 200804 632130
rect 214392 629898 214420 632198
rect 223948 632120 224000 632126
rect 223948 632062 224000 632068
rect 223960 629898 223988 632062
rect 214392 629870 214682 629898
rect 223960 629870 224342 629898
rect 204364 629326 205022 629354
rect 202786 620256 202842 620265
rect 202786 620191 202842 620200
rect 202800 611318 202828 620191
rect 202788 611312 202840 611318
rect 202788 611254 202840 611260
rect 200764 608592 200816 608598
rect 200764 608534 200816 608540
rect 204364 608462 204392 629326
rect 224512 610722 224540 632198
rect 225604 632120 225656 632126
rect 225604 632062 225656 632068
rect 224342 610694 224540 610722
rect 205008 608598 205036 610028
rect 204996 608592 205048 608598
rect 204996 608534 205048 608540
rect 178040 608456 178092 608462
rect 178040 608398 178092 608404
rect 187700 608456 187752 608462
rect 187700 608398 187752 608404
rect 199384 608456 199436 608462
rect 199384 608398 199436 608404
rect 204352 608456 204404 608462
rect 204352 608398 204404 608404
rect 214668 608394 214696 610028
rect 225616 608394 225644 632062
rect 232332 629898 232360 632266
rect 241520 632256 241572 632262
rect 241520 632198 241572 632204
rect 232070 629870 232360 629898
rect 241532 629898 241560 632198
rect 251456 632188 251508 632194
rect 251456 632130 251508 632136
rect 251180 632120 251232 632126
rect 251180 632062 251232 632068
rect 251192 629898 251220 632062
rect 241532 629870 241730 629898
rect 251192 629870 251390 629898
rect 230386 620256 230442 620265
rect 230386 620191 230442 620200
rect 226338 619576 226394 619585
rect 226338 619511 226394 619520
rect 226352 611250 226380 619511
rect 230400 611250 230428 620191
rect 226340 611244 226392 611250
rect 226340 611186 226392 611192
rect 230388 611244 230440 611250
rect 230388 611186 230440 611192
rect 251468 610722 251496 632130
rect 251390 610694 251496 610722
rect 232056 608462 232084 610028
rect 241716 608462 241744 610028
rect 251836 608598 251864 632266
rect 413468 632256 413520 632262
rect 413468 632198 413520 632204
rect 430580 632256 430632 632262
rect 430580 632198 430632 632204
rect 440516 632256 440568 632262
rect 440516 632198 440568 632204
rect 457260 632256 457312 632262
rect 457260 632198 457312 632204
rect 468576 632256 468628 632262
rect 468576 632198 468628 632204
rect 268292 632188 268344 632194
rect 268292 632130 268344 632136
rect 279424 632188 279476 632194
rect 279424 632130 279476 632136
rect 295800 632188 295852 632194
rect 295800 632130 295852 632136
rect 305644 632188 305696 632194
rect 305644 632130 305696 632136
rect 322388 632188 322440 632194
rect 322388 632130 322440 632136
rect 336004 632188 336056 632194
rect 336004 632130 336056 632136
rect 349804 632188 349856 632194
rect 349804 632130 349856 632136
rect 359556 632188 359608 632194
rect 359556 632130 359608 632136
rect 376300 632188 376352 632194
rect 376300 632130 376352 632136
rect 386512 632188 386564 632194
rect 386512 632130 386564 632136
rect 403348 632188 403400 632194
rect 403348 632130 403400 632136
rect 253204 632120 253256 632126
rect 253204 632062 253256 632068
rect 251824 608592 251876 608598
rect 251824 608534 251876 608540
rect 253216 608462 253244 632062
rect 268304 629898 268332 632130
rect 278044 632120 278096 632126
rect 278044 632062 278096 632068
rect 278056 629898 278084 632062
rect 268304 629870 268686 629898
rect 278056 629870 278346 629898
rect 258184 629326 259026 629354
rect 256606 620256 256662 620265
rect 256606 620191 256662 620200
rect 253938 619032 253994 619041
rect 253938 618967 253994 618976
rect 253952 611318 253980 618967
rect 256620 611318 256648 620191
rect 253940 611312 253992 611318
rect 253940 611254 253992 611260
rect 256608 611312 256660 611318
rect 256608 611254 256660 611260
rect 258184 608462 258212 629326
rect 279436 615494 279464 632130
rect 279516 632120 279568 632126
rect 279516 632062 279568 632068
rect 278792 615466 279464 615494
rect 278792 610722 278820 615466
rect 278346 610694 278820 610722
rect 259012 608598 259040 610028
rect 259000 608592 259052 608598
rect 259000 608534 259052 608540
rect 232044 608456 232096 608462
rect 232044 608398 232096 608404
rect 241704 608456 241756 608462
rect 241704 608398 241756 608404
rect 253204 608456 253256 608462
rect 253204 608398 253256 608404
rect 258172 608456 258224 608462
rect 258172 608398 258224 608404
rect 268672 608394 268700 610028
rect 279528 608394 279556 632062
rect 295812 629898 295840 632130
rect 305552 632120 305604 632126
rect 305552 632062 305604 632068
rect 305564 629898 305592 632062
rect 295734 629870 295840 629898
rect 305394 629870 305592 629898
rect 286074 629338 286180 629354
rect 285772 629332 285824 629338
rect 286074 629332 286192 629338
rect 286074 629326 286140 629332
rect 285772 629274 285824 629280
rect 286140 629274 286192 629280
rect 284206 619712 284262 619721
rect 284206 619647 284262 619656
rect 280158 619576 280214 619585
rect 280158 619511 280214 619520
rect 280172 611250 280200 619511
rect 284220 611250 284248 619647
rect 280160 611244 280212 611250
rect 280160 611186 280212 611192
rect 284208 611244 284260 611250
rect 284208 611186 284260 611192
rect 285784 608394 285812 629274
rect 305656 625154 305684 632130
rect 307024 632120 307076 632126
rect 307024 632062 307076 632068
rect 305472 625126 305684 625154
rect 305472 610722 305500 625126
rect 305394 610694 305500 610722
rect 286060 608462 286088 610028
rect 286048 608456 286100 608462
rect 286048 608398 286100 608404
rect 295720 608394 295748 610028
rect 307036 608394 307064 632062
rect 322400 629898 322428 632130
rect 331956 632120 332008 632126
rect 331956 632062 332008 632068
rect 333244 632120 333296 632126
rect 333244 632062 333296 632068
rect 331968 629898 331996 632062
rect 322400 629870 322690 629898
rect 331968 629870 332350 629898
rect 312004 629326 313030 629354
rect 311806 620256 311862 620265
rect 311806 620191 311862 620200
rect 307758 619576 307814 619585
rect 307758 619511 307814 619520
rect 307772 611318 307800 619511
rect 307760 611312 307812 611318
rect 307760 611254 307812 611260
rect 311820 611182 311848 620191
rect 311808 611176 311860 611182
rect 311808 611118 311860 611124
rect 312004 608394 312032 629326
rect 332350 610706 332640 610722
rect 332350 610700 332652 610706
rect 332350 610694 332600 610700
rect 332600 610642 332652 610648
rect 313016 608462 313044 610028
rect 313004 608456 313056 608462
rect 313004 608398 313056 608404
rect 322676 608394 322704 610028
rect 333256 608394 333284 632062
rect 335358 619576 335414 619585
rect 335358 619511 335414 619520
rect 335372 611250 335400 619511
rect 335360 611244 335412 611250
rect 335360 611186 335412 611192
rect 336016 610706 336044 632130
rect 349816 629898 349844 632130
rect 359464 632120 359516 632126
rect 359464 632062 359516 632068
rect 359476 629898 359504 632062
rect 349738 629870 349844 629898
rect 359398 629870 359504 629898
rect 340078 629338 340184 629354
rect 339592 629332 339644 629338
rect 340078 629332 340196 629338
rect 340078 629326 340144 629332
rect 339592 629274 339644 629280
rect 340144 629274 340196 629280
rect 338026 620256 338082 620265
rect 338026 620191 338082 620200
rect 338040 611318 338068 620191
rect 338028 611312 338080 611318
rect 338028 611254 338080 611260
rect 336004 610700 336056 610706
rect 336004 610642 336056 610648
rect 339604 608394 339632 629274
rect 359568 628810 359596 632130
rect 359740 632120 359792 632126
rect 359740 632062 359792 632068
rect 359476 628782 359596 628810
rect 359476 610722 359504 628782
rect 359752 628538 359780 632062
rect 376312 629898 376340 632130
rect 386052 632120 386104 632126
rect 386052 632062 386104 632068
rect 386064 629898 386092 632062
rect 376312 629870 376694 629898
rect 386064 629870 386354 629898
rect 359398 610694 359504 610722
rect 359568 628510 359780 628538
rect 365824 629326 367034 629354
rect 340064 608462 340092 610028
rect 340052 608456 340104 608462
rect 340052 608398 340104 608404
rect 349724 608394 349752 610028
rect 359568 608394 359596 628510
rect 365626 620256 365682 620265
rect 365626 620191 365682 620200
rect 361578 619032 361634 619041
rect 361578 618967 361634 618976
rect 361592 611182 361620 618967
rect 365640 611250 365668 620191
rect 365628 611244 365680 611250
rect 365628 611186 365680 611192
rect 361580 611176 361632 611182
rect 361580 611118 361632 611124
rect 365824 608394 365852 629326
rect 386524 610722 386552 632130
rect 387064 632120 387116 632126
rect 387064 632062 387116 632068
rect 386354 610694 386552 610722
rect 367020 608462 367048 610028
rect 367008 608456 367060 608462
rect 367008 608398 367060 608404
rect 376680 608394 376708 610028
rect 387076 608394 387104 632062
rect 403360 629898 403388 632130
rect 413008 632120 413060 632126
rect 413008 632062 413060 632068
rect 413020 629898 413048 632062
rect 403360 629870 403650 629898
rect 413020 629870 413310 629898
rect 393424 629326 393990 629354
rect 391846 620256 391902 620265
rect 391846 620191 391902 620200
rect 389178 619576 389234 619585
rect 389178 619511 389234 619520
rect 389192 611318 389220 619511
rect 391860 611318 391888 620191
rect 389180 611312 389232 611318
rect 389180 611254 389232 611260
rect 391848 611312 391900 611318
rect 391848 611254 391900 611260
rect 393424 608394 393452 629326
rect 413480 610722 413508 632198
rect 421288 632188 421340 632194
rect 421288 632130 421340 632136
rect 414664 632120 414716 632126
rect 414664 632062 414716 632068
rect 413402 610694 413508 610722
rect 393976 608462 394004 610028
rect 393964 608456 394016 608462
rect 393964 608398 394016 608404
rect 403728 608394 403756 610028
rect 414676 608394 414704 632062
rect 421300 629898 421328 632130
rect 421038 629870 421328 629898
rect 430592 629898 430620 632198
rect 440240 632120 440292 632126
rect 440240 632062 440292 632068
rect 440252 629898 440280 632062
rect 430592 629870 430698 629898
rect 440252 629870 440358 629898
rect 419446 620256 419502 620265
rect 419446 620191 419502 620200
rect 415398 619576 415454 619585
rect 415398 619511 415454 619520
rect 415412 611250 415440 619511
rect 419460 611250 419488 620191
rect 415400 611244 415452 611250
rect 415400 611186 415452 611192
rect 419448 611244 419500 611250
rect 419448 611186 419500 611192
rect 440528 610722 440556 632198
rect 445024 632188 445076 632194
rect 445024 632130 445076 632136
rect 442264 632120 442316 632126
rect 442264 632062 442316 632068
rect 440358 610694 440556 610722
rect 421024 608462 421052 610028
rect 430684 608462 430712 610028
rect 442276 608462 442304 632062
rect 442998 619576 443054 619585
rect 442998 619511 443054 619520
rect 443012 611318 443040 619511
rect 443000 611312 443052 611318
rect 443000 611254 443052 611260
rect 445036 611182 445064 632130
rect 457272 629898 457300 632198
rect 467012 632120 467064 632126
rect 467012 632062 467064 632068
rect 468484 632120 468536 632126
rect 468484 632062 468536 632068
rect 467024 629898 467052 632062
rect 457272 629870 457654 629898
rect 467024 629870 467314 629898
rect 447244 629326 447994 629354
rect 445666 620256 445722 620265
rect 445666 620191 445722 620200
rect 445680 611318 445708 620191
rect 445668 611312 445720 611318
rect 445668 611254 445720 611260
rect 445024 611176 445076 611182
rect 445024 611118 445076 611124
rect 447244 608462 447272 629326
rect 447692 611176 447744 611182
rect 447692 611118 447744 611124
rect 467656 611176 467708 611182
rect 467656 611118 467708 611124
rect 447704 610722 447732 611118
rect 467668 610722 467696 611118
rect 447704 610694 447994 610722
rect 467406 610694 467696 610722
rect 421012 608456 421064 608462
rect 421012 608398 421064 608404
rect 430672 608456 430724 608462
rect 430672 608398 430724 608404
rect 442264 608456 442316 608462
rect 442264 608398 442316 608404
rect 447232 608456 447284 608462
rect 447232 608398 447284 608404
rect 457732 608394 457760 610028
rect 468496 608394 468524 632062
rect 468588 611182 468616 632198
rect 475396 629898 475424 632266
rect 484400 632256 484452 632262
rect 484400 632198 484452 632204
rect 475042 629870 475424 629898
rect 484412 629898 484440 632198
rect 494520 632188 494572 632194
rect 494520 632130 494572 632136
rect 494060 632120 494112 632126
rect 494060 632062 494112 632068
rect 494072 629898 494100 632062
rect 484412 629870 484702 629898
rect 494072 629870 494362 629898
rect 473266 619712 473322 619721
rect 473266 619647 473322 619656
rect 469218 619032 469274 619041
rect 469218 618967 469274 618976
rect 469232 611250 469260 618967
rect 473280 611250 473308 619647
rect 469220 611244 469272 611250
rect 469220 611186 469272 611192
rect 473268 611244 473320 611250
rect 473268 611186 473320 611192
rect 468576 611176 468628 611182
rect 468576 611118 468628 611124
rect 494532 610722 494560 632130
rect 494362 610694 494560 610722
rect 475028 608462 475056 610028
rect 484688 608462 484716 610028
rect 494716 608598 494744 632266
rect 511356 632188 511408 632194
rect 511356 632130 511408 632136
rect 522304 632188 522356 632194
rect 522304 632130 522356 632136
rect 496084 632120 496136 632126
rect 496084 632062 496136 632068
rect 494704 608592 494756 608598
rect 494704 608534 494756 608540
rect 496096 608462 496124 632062
rect 511368 629898 511396 632130
rect 520924 632120 520976 632126
rect 520924 632062 520976 632068
rect 520936 629898 520964 632062
rect 511368 629870 511658 629898
rect 520936 629870 521318 629898
rect 501064 629326 501998 629354
rect 500866 620256 500922 620265
rect 500866 620191 500922 620200
rect 496818 619576 496874 619585
rect 496818 619511 496874 619520
rect 496832 611318 496860 619511
rect 500880 611318 500908 620191
rect 496820 611312 496872 611318
rect 496820 611254 496872 611260
rect 500868 611312 500920 611318
rect 500868 611254 500920 611260
rect 501064 608462 501092 629326
rect 522316 615494 522344 632130
rect 522396 632120 522448 632126
rect 522396 632062 522448 632068
rect 521856 615466 522344 615494
rect 521856 610722 521884 615466
rect 521410 610694 521884 610722
rect 501984 608598 502012 610028
rect 501972 608592 502024 608598
rect 501972 608534 502024 608540
rect 475016 608456 475068 608462
rect 475016 608398 475068 608404
rect 484676 608456 484728 608462
rect 484676 608398 484728 608404
rect 496084 608456 496136 608462
rect 496084 608398 496136 608404
rect 501052 608456 501104 608462
rect 501052 608398 501104 608404
rect 511736 608394 511764 610028
rect 522408 608394 522436 632062
rect 526444 629944 526496 629950
rect 526444 629886 526496 629892
rect 526456 620401 526484 629886
rect 526442 620392 526498 620401
rect 526442 620327 526498 620336
rect 523038 619576 523094 619585
rect 523038 619511 523094 619520
rect 523052 611250 523080 619511
rect 523040 611244 523092 611250
rect 523040 611186 523092 611192
rect 160652 608388 160704 608394
rect 160652 608330 160704 608336
rect 171784 608388 171836 608394
rect 171784 608330 171836 608336
rect 214656 608388 214708 608394
rect 214656 608330 214708 608336
rect 225604 608388 225656 608394
rect 225604 608330 225656 608336
rect 268660 608388 268712 608394
rect 268660 608330 268712 608336
rect 279516 608388 279568 608394
rect 279516 608330 279568 608336
rect 285772 608388 285824 608394
rect 285772 608330 285824 608336
rect 295708 608388 295760 608394
rect 295708 608330 295760 608336
rect 307024 608388 307076 608394
rect 307024 608330 307076 608336
rect 311992 608388 312044 608394
rect 311992 608330 312044 608336
rect 322664 608388 322716 608394
rect 322664 608330 322716 608336
rect 333244 608388 333296 608394
rect 333244 608330 333296 608336
rect 339592 608388 339644 608394
rect 339592 608330 339644 608336
rect 349712 608388 349764 608394
rect 349712 608330 349764 608336
rect 359556 608388 359608 608394
rect 359556 608330 359608 608336
rect 365812 608388 365864 608394
rect 365812 608330 365864 608336
rect 376668 608388 376720 608394
rect 376668 608330 376720 608336
rect 387064 608388 387116 608394
rect 387064 608330 387116 608336
rect 393412 608388 393464 608394
rect 393412 608330 393464 608336
rect 403716 608388 403768 608394
rect 403716 608330 403768 608336
rect 414664 608388 414716 608394
rect 414664 608330 414716 608336
rect 457720 608388 457772 608394
rect 457720 608330 457772 608336
rect 468484 608388 468536 608394
rect 468484 608330 468536 608336
rect 511724 608388 511776 608394
rect 511724 608330 511776 608336
rect 522396 608388 522448 608394
rect 522396 608330 522448 608336
rect 232044 604716 232096 604722
rect 232044 604658 232096 604664
rect 251824 604716 251876 604722
rect 251824 604658 251876 604664
rect 475016 604716 475068 604722
rect 475016 604658 475068 604664
rect 494704 604716 494756 604722
rect 494704 604658 494756 604664
rect 170496 604648 170548 604654
rect 170496 604590 170548 604596
rect 187700 604648 187752 604654
rect 187700 604590 187752 604596
rect 197452 604648 197504 604654
rect 197452 604590 197504 604596
rect 214656 604648 214708 604654
rect 214656 604590 214708 604596
rect 224500 604648 224552 604654
rect 224500 604590 224552 604596
rect 170312 604580 170364 604586
rect 170312 604522 170364 604528
rect 160652 604512 160704 604518
rect 160652 604454 160704 604460
rect 160664 602956 160692 604454
rect 170324 602956 170352 604522
rect 150544 602262 151018 602290
rect 148966 593192 149022 593201
rect 148966 593127 149022 593136
rect 148980 583710 149008 593127
rect 148968 583704 149020 583710
rect 148968 583646 149020 583652
rect 148324 580916 148376 580922
rect 148324 580858 148376 580864
rect 150544 580854 150572 602262
rect 170508 583574 170536 604590
rect 178040 604580 178092 604586
rect 178040 604522 178092 604528
rect 171784 604512 171836 604518
rect 171784 604454 171836 604460
rect 170220 583568 170272 583574
rect 170496 583568 170548 583574
rect 170272 583516 170338 583522
rect 170220 583510 170338 583516
rect 170496 583510 170548 583516
rect 170232 583494 170338 583510
rect 150728 583086 151018 583114
rect 160572 583086 160678 583114
rect 150532 580848 150584 580854
rect 150532 580790 150584 580796
rect 150728 580786 150756 583086
rect 160572 580786 160600 583086
rect 171796 580786 171824 604454
rect 178052 602956 178080 604522
rect 187712 602956 187740 604590
rect 197360 604512 197412 604518
rect 197360 604454 197412 604460
rect 197372 602956 197400 604454
rect 176566 592648 176622 592657
rect 176566 592583 176622 592592
rect 172518 592512 172574 592521
rect 172518 592447 172574 592456
rect 172532 583642 172560 592447
rect 176580 583642 176608 592583
rect 197464 583794 197492 604590
rect 200764 604580 200816 604586
rect 200764 604522 200816 604528
rect 199384 604512 199436 604518
rect 199384 604454 199436 604460
rect 197386 583766 197492 583794
rect 172520 583636 172572 583642
rect 172520 583578 172572 583584
rect 176568 583636 176620 583642
rect 176568 583578 176620 583584
rect 178066 583086 178172 583114
rect 187726 583086 188016 583114
rect 178144 580854 178172 583086
rect 187988 580854 188016 583086
rect 199396 580854 199424 604454
rect 200118 592512 200174 592521
rect 200118 592447 200174 592456
rect 200132 583710 200160 592447
rect 200120 583704 200172 583710
rect 200120 583646 200172 583652
rect 200776 583574 200804 604522
rect 214668 602956 214696 604590
rect 224316 604512 224368 604518
rect 224316 604454 224368 604460
rect 224328 602956 224356 604454
rect 204364 602262 205022 602290
rect 202786 593192 202842 593201
rect 202786 593127 202842 593136
rect 202800 583710 202828 593127
rect 202788 583704 202840 583710
rect 202788 583646 202840 583652
rect 200764 583568 200816 583574
rect 200764 583510 200816 583516
rect 204364 580854 204392 602262
rect 224512 583794 224540 604590
rect 225604 604512 225656 604518
rect 225604 604454 225656 604460
rect 224342 583766 224540 583794
rect 204628 583568 204680 583574
rect 204680 583516 205022 583522
rect 204628 583510 205022 583516
rect 204640 583494 205022 583510
rect 214682 583086 215064 583114
rect 178132 580848 178184 580854
rect 178132 580790 178184 580796
rect 187976 580848 188028 580854
rect 187976 580790 188028 580796
rect 199384 580848 199436 580854
rect 199384 580790 199436 580796
rect 204352 580848 204404 580854
rect 204352 580790 204404 580796
rect 215036 580786 215064 583086
rect 225616 580786 225644 604454
rect 232056 602956 232084 604658
rect 241704 604648 241756 604654
rect 241704 604590 241756 604596
rect 241716 602956 241744 604590
rect 251456 604580 251508 604586
rect 251456 604522 251508 604528
rect 251364 604512 251416 604518
rect 251364 604454 251416 604460
rect 251376 602956 251404 604454
rect 230386 593192 230442 593201
rect 230386 593127 230442 593136
rect 226338 592512 226394 592521
rect 226338 592447 226394 592456
rect 226352 583642 226380 592447
rect 230400 583642 230428 593127
rect 251468 583794 251496 604522
rect 251390 583766 251496 583794
rect 226340 583636 226392 583642
rect 226340 583578 226392 583584
rect 230388 583636 230440 583642
rect 230388 583578 230440 583584
rect 231872 583086 232070 583114
rect 241730 583086 242112 583114
rect 231872 580854 231900 583086
rect 242084 580854 242112 583086
rect 251836 580990 251864 604658
rect 413468 604648 413520 604654
rect 413468 604590 413520 604596
rect 430672 604648 430724 604654
rect 430672 604590 430724 604596
rect 440516 604648 440568 604654
rect 440516 604590 440568 604596
rect 457628 604648 457680 604654
rect 457628 604590 457680 604596
rect 468576 604648 468628 604654
rect 468576 604590 468628 604596
rect 268660 604580 268712 604586
rect 268660 604522 268712 604528
rect 279516 604580 279568 604586
rect 279516 604522 279568 604528
rect 295708 604580 295760 604586
rect 295708 604522 295760 604528
rect 305460 604580 305512 604586
rect 305460 604522 305512 604528
rect 322664 604580 322716 604586
rect 322664 604522 322716 604528
rect 336004 604580 336056 604586
rect 336004 604522 336056 604528
rect 349712 604580 349764 604586
rect 349712 604522 349764 604528
rect 359464 604580 359516 604586
rect 359464 604522 359516 604528
rect 376668 604580 376720 604586
rect 376668 604522 376720 604528
rect 386512 604580 386564 604586
rect 386512 604522 386564 604528
rect 403624 604580 403676 604586
rect 403624 604522 403676 604528
rect 253204 604512 253256 604518
rect 253204 604454 253256 604460
rect 251824 580984 251876 580990
rect 251824 580926 251876 580932
rect 253216 580854 253244 604454
rect 268672 602956 268700 604522
rect 278320 604512 278372 604518
rect 278320 604454 278372 604460
rect 279424 604512 279476 604518
rect 279424 604454 279476 604460
rect 278332 602956 278360 604454
rect 258184 602262 259026 602290
rect 256606 593192 256662 593201
rect 256606 593127 256662 593136
rect 253938 592104 253994 592113
rect 253938 592039 253994 592048
rect 253952 583710 253980 592039
rect 256620 583710 256648 593127
rect 253940 583704 253992 583710
rect 253940 583646 253992 583652
rect 256608 583704 256660 583710
rect 256608 583646 256660 583652
rect 258184 580854 258212 602262
rect 278780 584792 278832 584798
rect 278780 584734 278832 584740
rect 278792 583658 278820 584734
rect 278346 583630 278820 583658
rect 258736 583086 259026 583114
rect 268686 583086 268976 583114
rect 258736 580990 258764 583086
rect 258724 580984 258776 580990
rect 258724 580926 258776 580932
rect 231860 580848 231912 580854
rect 231860 580790 231912 580796
rect 242072 580848 242124 580854
rect 242072 580790 242124 580796
rect 253204 580848 253256 580854
rect 253204 580790 253256 580796
rect 258172 580848 258224 580854
rect 258172 580790 258224 580796
rect 268948 580786 268976 583086
rect 279436 580786 279464 604454
rect 279528 584798 279556 604522
rect 285784 603078 286088 603106
rect 284206 592648 284262 592657
rect 284206 592583 284262 592592
rect 280158 592512 280214 592521
rect 280158 592447 280214 592456
rect 279516 584792 279568 584798
rect 279516 584734 279568 584740
rect 280172 583642 280200 592447
rect 284220 583642 284248 592583
rect 280160 583636 280212 583642
rect 280160 583578 280212 583584
rect 284208 583636 284260 583642
rect 284208 583578 284260 583584
rect 285784 580786 285812 603078
rect 286060 602956 286088 603078
rect 295720 602956 295748 604522
rect 305368 604512 305420 604518
rect 305368 604454 305420 604460
rect 305380 602956 305408 604454
rect 305472 583794 305500 604522
rect 307024 604512 307076 604518
rect 307024 604454 307076 604460
rect 305394 583766 305500 583794
rect 286074 583086 286180 583114
rect 295734 583086 296024 583114
rect 286152 580854 286180 583086
rect 286140 580848 286192 580854
rect 286140 580790 286192 580796
rect 295996 580786 296024 583086
rect 307036 580786 307064 604454
rect 322676 602956 322704 604522
rect 332324 604512 332376 604518
rect 332324 604454 332376 604460
rect 333244 604512 333296 604518
rect 333244 604454 333296 604460
rect 332336 602956 332364 604454
rect 312004 602262 313030 602290
rect 311806 593192 311862 593201
rect 311806 593127 311862 593136
rect 307758 592512 307814 592521
rect 307758 592447 307814 592456
rect 307772 583710 307800 592447
rect 307760 583704 307812 583710
rect 307760 583646 307812 583652
rect 311820 583574 311848 593127
rect 311808 583568 311860 583574
rect 311808 583510 311860 583516
rect 312004 580786 312032 602262
rect 332600 583704 332652 583710
rect 332350 583652 332600 583658
rect 332350 583646 332652 583652
rect 332350 583630 332640 583646
rect 312648 583086 313030 583114
rect 322690 583086 322888 583114
rect 312648 580854 312676 583086
rect 312636 580848 312688 580854
rect 312636 580790 312688 580796
rect 322860 580786 322888 583086
rect 333256 580786 333284 604454
rect 335358 592512 335414 592521
rect 335358 592447 335414 592456
rect 335372 583642 335400 592447
rect 336016 583710 336044 604522
rect 339604 603078 340092 603106
rect 338026 593192 338082 593201
rect 338026 593127 338082 593136
rect 338040 583710 338068 593127
rect 336004 583704 336056 583710
rect 336004 583646 336056 583652
rect 338028 583704 338080 583710
rect 338028 583646 338080 583652
rect 335360 583636 335412 583642
rect 335360 583578 335412 583584
rect 339604 580786 339632 603078
rect 340064 602956 340092 603078
rect 349724 602956 349752 604522
rect 359372 604512 359424 604518
rect 359372 604454 359424 604460
rect 359384 602956 359412 604454
rect 359476 583794 359504 604522
rect 359556 604512 359608 604518
rect 359556 604454 359608 604460
rect 359398 583766 359504 583794
rect 340078 583086 340184 583114
rect 349738 583086 350120 583114
rect 340156 580854 340184 583086
rect 340144 580848 340196 580854
rect 340144 580790 340196 580796
rect 350092 580786 350120 583086
rect 359568 580786 359596 604454
rect 376680 602956 376708 604522
rect 386328 604512 386380 604518
rect 386328 604454 386380 604460
rect 386340 602956 386368 604454
rect 365824 602262 367034 602290
rect 365626 593192 365682 593201
rect 365626 593127 365682 593136
rect 361578 592104 361634 592113
rect 361578 592039 361634 592048
rect 361592 583574 361620 592039
rect 365640 583642 365668 593127
rect 365628 583636 365680 583642
rect 365628 583578 365680 583584
rect 361580 583568 361632 583574
rect 361580 583510 361632 583516
rect 365824 580786 365852 602262
rect 386524 583794 386552 604522
rect 387064 604512 387116 604518
rect 387064 604454 387116 604460
rect 386354 583766 386552 583794
rect 366744 583086 367034 583114
rect 376588 583086 376694 583114
rect 366744 580854 366772 583086
rect 366732 580848 366784 580854
rect 366732 580790 366784 580796
rect 376588 580786 376616 583086
rect 387076 580786 387104 604454
rect 403636 602956 403664 604522
rect 413284 604512 413336 604518
rect 413284 604454 413336 604460
rect 413296 602956 413324 604454
rect 393424 602262 393990 602290
rect 391846 592648 391902 592657
rect 391846 592583 391902 592592
rect 389178 592512 389234 592521
rect 389178 592447 389234 592456
rect 389192 583710 389220 592447
rect 391860 583710 391888 592583
rect 389180 583704 389232 583710
rect 389180 583646 389232 583652
rect 391848 583704 391900 583710
rect 391848 583646 391900 583652
rect 393424 580786 393452 602262
rect 413480 583794 413508 604590
rect 421012 604580 421064 604586
rect 421012 604522 421064 604528
rect 414664 604512 414716 604518
rect 414664 604454 414716 604460
rect 413402 583766 413508 583794
rect 393608 583086 393990 583114
rect 403742 583086 404032 583114
rect 393608 580854 393636 583086
rect 393596 580848 393648 580854
rect 393596 580790 393648 580796
rect 404004 580786 404032 583086
rect 414676 580786 414704 604454
rect 421024 602956 421052 604522
rect 430684 602956 430712 604590
rect 440332 604512 440384 604518
rect 440332 604454 440384 604460
rect 440344 602956 440372 604454
rect 419446 593192 419502 593201
rect 419446 593127 419502 593136
rect 415398 592512 415454 592521
rect 415398 592447 415454 592456
rect 415412 583642 415440 592447
rect 419460 583642 419488 593127
rect 440528 583794 440556 604590
rect 445024 604580 445076 604586
rect 445024 604522 445076 604528
rect 442264 604512 442316 604518
rect 442264 604454 442316 604460
rect 440358 583766 440556 583794
rect 415400 583636 415452 583642
rect 415400 583578 415452 583584
rect 419448 583636 419500 583642
rect 419448 583578 419500 583584
rect 420932 583086 421038 583114
rect 430698 583086 431080 583114
rect 420932 580854 420960 583086
rect 431052 580854 431080 583086
rect 442276 580854 442304 604454
rect 442998 592512 443054 592521
rect 442998 592447 443054 592456
rect 443012 583710 443040 592447
rect 445036 583778 445064 604522
rect 457640 602956 457668 604590
rect 467288 604512 467340 604518
rect 467288 604454 467340 604460
rect 468484 604512 468536 604518
rect 468484 604454 468536 604460
rect 467300 602956 467328 604454
rect 447244 602262 447994 602290
rect 445666 593192 445722 593201
rect 445666 593127 445722 593136
rect 445024 583772 445076 583778
rect 445024 583714 445076 583720
rect 445680 583710 445708 593127
rect 443000 583704 443052 583710
rect 443000 583646 443052 583652
rect 445668 583704 445720 583710
rect 445668 583646 445720 583652
rect 447244 580854 447272 602262
rect 447692 583772 447744 583778
rect 447692 583714 447744 583720
rect 447704 583658 447732 583714
rect 447704 583630 447994 583658
rect 467656 583568 467708 583574
rect 467406 583516 467656 583522
rect 467406 583510 467708 583516
rect 467406 583494 467696 583510
rect 457746 583086 458128 583114
rect 420920 580848 420972 580854
rect 420920 580790 420972 580796
rect 431040 580848 431092 580854
rect 431040 580790 431092 580796
rect 442264 580848 442316 580854
rect 442264 580790 442316 580796
rect 447232 580848 447284 580854
rect 447232 580790 447284 580796
rect 458100 580786 458128 583086
rect 468496 580786 468524 604454
rect 468588 583574 468616 604590
rect 475028 602956 475056 604658
rect 484676 604648 484728 604654
rect 484676 604590 484728 604596
rect 484688 602956 484716 604590
rect 494520 604580 494572 604586
rect 494520 604522 494572 604528
rect 494336 604512 494388 604518
rect 494336 604454 494388 604460
rect 494348 602956 494376 604454
rect 473266 592648 473322 592657
rect 473266 592583 473322 592592
rect 469218 592104 469274 592113
rect 469218 592039 469274 592048
rect 469232 583642 469260 592039
rect 473280 583642 473308 592583
rect 494532 583794 494560 604522
rect 494362 583766 494560 583794
rect 469220 583636 469272 583642
rect 469220 583578 469272 583584
rect 473268 583636 473320 583642
rect 473268 583578 473320 583584
rect 468576 583568 468628 583574
rect 468576 583510 468628 583516
rect 474752 583086 475042 583114
rect 484702 583086 484992 583114
rect 474752 580854 474780 583086
rect 484964 580854 484992 583086
rect 494716 580990 494744 604658
rect 511632 604580 511684 604586
rect 511632 604522 511684 604528
rect 522304 604580 522356 604586
rect 522304 604522 522356 604528
rect 496084 604512 496136 604518
rect 496084 604454 496136 604460
rect 494704 580984 494756 580990
rect 494704 580926 494756 580932
rect 496096 580854 496124 604454
rect 511644 602956 511672 604522
rect 521292 604512 521344 604518
rect 521292 604454 521344 604460
rect 521304 602956 521332 604454
rect 501064 602262 501998 602290
rect 500866 593192 500922 593201
rect 500866 593127 500922 593136
rect 496818 592512 496874 592521
rect 496818 592447 496874 592456
rect 496832 583710 496860 592447
rect 500880 583710 500908 593127
rect 496820 583704 496872 583710
rect 496820 583646 496872 583652
rect 500868 583704 500920 583710
rect 500868 583646 500920 583652
rect 501064 580854 501092 602262
rect 522316 586514 522344 604522
rect 522396 604512 522448 604518
rect 522396 604454 522448 604460
rect 521856 586486 522344 586514
rect 521856 583658 521884 586486
rect 521410 583630 521884 583658
rect 501616 583086 501998 583114
rect 511750 583086 511948 583114
rect 501616 580990 501644 583086
rect 501604 580984 501656 580990
rect 501604 580926 501656 580932
rect 474740 580848 474792 580854
rect 474740 580790 474792 580796
rect 484952 580848 485004 580854
rect 484952 580790 485004 580796
rect 496084 580848 496136 580854
rect 496084 580790 496136 580796
rect 501052 580848 501104 580854
rect 501052 580790 501104 580796
rect 511920 580786 511948 583086
rect 522408 580786 522436 604454
rect 526444 602404 526496 602410
rect 526444 602346 526496 602352
rect 526456 593337 526484 602346
rect 526442 593328 526498 593337
rect 526442 593263 526498 593272
rect 523038 592512 523094 592521
rect 523038 592447 523094 592456
rect 523052 583642 523080 592447
rect 523040 583636 523092 583642
rect 523040 583578 523092 583584
rect 150716 580780 150768 580786
rect 150716 580722 150768 580728
rect 160560 580780 160612 580786
rect 160560 580722 160612 580728
rect 171784 580780 171836 580786
rect 171784 580722 171836 580728
rect 215024 580780 215076 580786
rect 215024 580722 215076 580728
rect 225604 580780 225656 580786
rect 225604 580722 225656 580728
rect 268936 580780 268988 580786
rect 268936 580722 268988 580728
rect 279424 580780 279476 580786
rect 279424 580722 279476 580728
rect 285772 580780 285824 580786
rect 285772 580722 285824 580728
rect 295984 580780 296036 580786
rect 295984 580722 296036 580728
rect 307024 580780 307076 580786
rect 307024 580722 307076 580728
rect 311992 580780 312044 580786
rect 311992 580722 312044 580728
rect 322848 580780 322900 580786
rect 322848 580722 322900 580728
rect 333244 580780 333296 580786
rect 333244 580722 333296 580728
rect 339592 580780 339644 580786
rect 339592 580722 339644 580728
rect 350080 580780 350132 580786
rect 350080 580722 350132 580728
rect 359556 580780 359608 580786
rect 359556 580722 359608 580728
rect 365812 580780 365864 580786
rect 365812 580722 365864 580728
rect 376576 580780 376628 580786
rect 376576 580722 376628 580728
rect 387064 580780 387116 580786
rect 387064 580722 387116 580728
rect 393412 580780 393464 580786
rect 393412 580722 393464 580728
rect 403992 580780 404044 580786
rect 403992 580722 404044 580728
rect 414664 580780 414716 580786
rect 414664 580722 414716 580728
rect 458088 580780 458140 580786
rect 458088 580722 458140 580728
rect 468484 580780 468536 580786
rect 468484 580722 468536 580728
rect 511908 580780 511960 580786
rect 511908 580722 511960 580728
rect 522396 580780 522448 580786
rect 522396 580722 522448 580728
rect 149704 578536 149756 578542
rect 149704 578478 149756 578484
rect 148966 566264 149022 566273
rect 148966 566199 149022 566208
rect 148980 557530 149008 566199
rect 148968 557524 149020 557530
rect 148968 557466 149020 557472
rect 146944 554736 146996 554742
rect 146944 554678 146996 554684
rect 124036 554668 124088 554674
rect 124036 554610 124088 554616
rect 133696 554668 133748 554674
rect 133696 554610 133748 554616
rect 144276 554668 144328 554674
rect 144276 554610 144328 554616
rect 79692 554600 79744 554606
rect 79692 554542 79744 554548
rect 90364 554600 90416 554606
rect 90364 554542 90416 554548
rect 106648 554600 106700 554606
rect 106648 554542 106700 554548
rect 116584 554600 116636 554606
rect 116584 554542 116636 554548
rect 122932 554600 122984 554606
rect 122932 554542 122984 554548
rect 146944 550928 146996 550934
rect 146944 550870 146996 550876
rect 52644 550860 52696 550866
rect 52644 550802 52696 550808
rect 43076 550656 43128 550662
rect 43076 550598 43128 550604
rect 43088 548964 43116 550598
rect 52656 548964 52684 550802
rect 62488 550792 62540 550798
rect 62488 550734 62540 550740
rect 79692 550792 79744 550798
rect 79692 550734 79744 550740
rect 90456 550792 90508 550798
rect 90456 550734 90508 550740
rect 106648 550792 106700 550798
rect 106648 550734 106700 550740
rect 116492 550792 116544 550798
rect 116492 550734 116544 550740
rect 133696 550792 133748 550798
rect 133696 550734 133748 550740
rect 62304 550724 62356 550730
rect 62304 550666 62356 550672
rect 62316 548964 62344 550666
rect 37924 548548 37976 548554
rect 37924 548490 37976 548496
rect 41326 539200 41382 539209
rect 41326 539135 41382 539144
rect 37922 538248 37978 538257
rect 37922 538183 37978 538192
rect 36820 526992 36872 526998
rect 36820 526934 36872 526940
rect 36820 523252 36872 523258
rect 36820 523194 36872 523200
rect 36832 502314 36860 523194
rect 37936 522306 37964 538183
rect 41340 529854 41368 539135
rect 41328 529848 41380 529854
rect 41328 529790 41380 529796
rect 62500 529666 62528 550734
rect 64144 550724 64196 550730
rect 64144 550666 64196 550672
rect 62764 550656 62816 550662
rect 62764 550598 62816 550604
rect 62422 529638 62528 529666
rect 42812 529094 43010 529122
rect 52762 529094 53144 529122
rect 42812 527066 42840 529094
rect 53116 527134 53144 529094
rect 53104 527128 53156 527134
rect 53104 527070 53156 527076
rect 62776 527066 62804 550598
rect 64156 527134 64184 550666
rect 79704 548964 79732 550734
rect 89352 550724 89404 550730
rect 89352 550666 89404 550672
rect 90364 550724 90416 550730
rect 90364 550666 90416 550672
rect 89364 548964 89392 550666
rect 69124 548270 70058 548298
rect 68926 538656 68982 538665
rect 68926 538591 68982 538600
rect 64878 538520 64934 538529
rect 64878 538455 64934 538464
rect 64892 529922 64920 538455
rect 64880 529916 64932 529922
rect 64880 529858 64932 529864
rect 68940 529786 68968 538591
rect 68928 529780 68980 529786
rect 68928 529722 68980 529728
rect 69124 527134 69152 548270
rect 89720 533656 89772 533662
rect 89720 533598 89772 533604
rect 89732 529666 89760 533598
rect 89378 529638 89760 529666
rect 69768 529094 70058 529122
rect 79718 529094 80008 529122
rect 64144 527128 64196 527134
rect 64144 527070 64196 527076
rect 69112 527128 69164 527134
rect 69112 527070 69164 527076
rect 69768 527066 69796 529094
rect 42800 527060 42852 527066
rect 42800 527002 42852 527008
rect 62764 527060 62816 527066
rect 62764 527002 62816 527008
rect 69756 527060 69808 527066
rect 69756 527002 69808 527008
rect 79980 526998 80008 529094
rect 90376 526998 90404 550666
rect 90468 533662 90496 550734
rect 106660 548964 106688 550734
rect 116308 550724 116360 550730
rect 116308 550666 116360 550672
rect 116320 548964 116348 550666
rect 96724 548270 97014 548298
rect 95146 539200 95202 539209
rect 95146 539135 95202 539144
rect 91098 538520 91154 538529
rect 91098 538455 91154 538464
rect 90456 533656 90508 533662
rect 90456 533598 90508 533604
rect 91112 529854 91140 538455
rect 95160 529922 95188 539135
rect 95148 529916 95200 529922
rect 95148 529858 95200 529864
rect 91100 529848 91152 529854
rect 91100 529790 91152 529796
rect 96724 527134 96752 548270
rect 116228 529650 116334 529666
rect 116504 529650 116532 550734
rect 116584 550724 116636 550730
rect 116584 550666 116636 550672
rect 116216 529644 116334 529650
rect 116268 529638 116334 529644
rect 116492 529644 116544 529650
rect 116216 529586 116268 529592
rect 116492 529586 116544 529592
rect 96816 529094 97014 529122
rect 106568 529094 106674 529122
rect 96712 527128 96764 527134
rect 96712 527070 96764 527076
rect 96816 527066 96844 529094
rect 96804 527060 96856 527066
rect 96804 527002 96856 527008
rect 106568 526998 106596 529094
rect 116596 526998 116624 550666
rect 133708 548964 133736 550734
rect 143356 550724 143408 550730
rect 143356 550666 143408 550672
rect 144276 550724 144328 550730
rect 144276 550666 144328 550672
rect 143368 548964 143396 550666
rect 144184 550656 144236 550662
rect 144184 550598 144236 550604
rect 122944 548270 124062 548298
rect 122746 539200 122802 539209
rect 122746 539135 122802 539144
rect 118698 538520 118754 538529
rect 118698 538455 118754 538464
rect 118712 529786 118740 538455
rect 122760 529854 122788 539135
rect 122748 529848 122800 529854
rect 122748 529790 122800 529796
rect 118700 529780 118752 529786
rect 118700 529722 118752 529728
rect 79968 526992 80020 526998
rect 79968 526934 80020 526940
rect 90364 526992 90416 526998
rect 90364 526934 90416 526940
rect 106556 526992 106608 526998
rect 106556 526934 106608 526940
rect 116584 526992 116636 526998
rect 116584 526934 116636 526940
rect 122944 526930 122972 548270
rect 144196 538214 144224 550598
rect 143736 538186 144224 538214
rect 143736 529666 143764 538186
rect 143382 529638 143764 529666
rect 123680 529094 124062 529122
rect 133722 529094 133828 529122
rect 123680 527066 123708 529094
rect 123668 527060 123720 527066
rect 123668 527002 123720 527008
rect 133800 526998 133828 529094
rect 144288 526998 144316 550666
rect 146298 538384 146354 538393
rect 146298 538319 146354 538328
rect 146312 529922 146340 538319
rect 146300 529916 146352 529922
rect 146300 529858 146352 529864
rect 133788 526992 133840 526998
rect 133788 526934 133840 526940
rect 144276 526992 144328 526998
rect 144276 526934 144328 526940
rect 122932 526924 122984 526930
rect 122932 526866 122984 526872
rect 52460 523252 52512 523258
rect 52460 523194 52512 523200
rect 43352 523048 43404 523054
rect 43352 522990 43404 522996
rect 37924 522300 37976 522306
rect 37924 522242 37976 522248
rect 43364 521914 43392 522990
rect 43102 521886 43392 521914
rect 52472 521914 52500 523194
rect 62488 523184 62540 523190
rect 62488 523126 62540 523132
rect 79324 523184 79376 523190
rect 79324 523126 79376 523132
rect 90456 523184 90508 523190
rect 90456 523126 90508 523132
rect 106372 523184 106424 523190
rect 106372 523126 106424 523132
rect 116492 523184 116544 523190
rect 116492 523126 116544 523132
rect 133420 523184 133472 523190
rect 133420 523126 133472 523132
rect 144184 523184 144236 523190
rect 144184 523126 144236 523132
rect 62120 523116 62172 523122
rect 62120 523058 62172 523064
rect 62132 521914 62160 523058
rect 52472 521886 52670 521914
rect 62132 521886 62330 521914
rect 41328 520396 41380 520402
rect 41328 520338 41380 520344
rect 41340 512417 41368 520338
rect 41326 512408 41382 512417
rect 41326 512343 41382 512352
rect 37922 511048 37978 511057
rect 37922 510983 37978 510992
rect 36820 502308 36872 502314
rect 36820 502250 36872 502256
rect 36728 500676 36780 500682
rect 36728 500618 36780 500624
rect 36728 497072 36780 497078
rect 36728 497014 36780 497020
rect 36740 475998 36768 497014
rect 36820 496936 36872 496942
rect 36820 496878 36872 496884
rect 36728 475992 36780 475998
rect 36728 475934 36780 475940
rect 36832 473210 36860 496878
rect 37936 494766 37964 510983
rect 62500 502738 62528 523126
rect 64144 523116 64196 523122
rect 64144 523058 64196 523064
rect 62764 523048 62816 523054
rect 62764 522990 62816 522996
rect 62422 502710 62528 502738
rect 42996 500886 43024 502044
rect 52748 500954 52776 502044
rect 52736 500948 52788 500954
rect 52736 500890 52788 500896
rect 62776 500886 62804 522990
rect 64156 500954 64184 523058
rect 79336 521914 79364 523126
rect 89076 523116 89128 523122
rect 89076 523058 89128 523064
rect 90364 523116 90416 523122
rect 90364 523058 90416 523064
rect 89088 521914 89116 523058
rect 79336 521886 79718 521914
rect 89088 521886 89378 521914
rect 69124 521206 70058 521234
rect 68928 520464 68980 520470
rect 68928 520406 68980 520412
rect 64880 520328 64932 520334
rect 64880 520270 64932 520276
rect 64892 511737 64920 520270
rect 68940 512961 68968 520406
rect 68926 512952 68982 512961
rect 68926 512887 68982 512896
rect 64878 511728 64934 511737
rect 64878 511663 64934 511672
rect 69124 500954 69152 521206
rect 89720 505640 89772 505646
rect 89720 505582 89772 505588
rect 89732 502738 89760 505582
rect 89378 502710 89760 502738
rect 64144 500948 64196 500954
rect 64144 500890 64196 500896
rect 69112 500948 69164 500954
rect 69112 500890 69164 500896
rect 70044 500886 70072 502044
rect 42984 500880 43036 500886
rect 42984 500822 43036 500828
rect 62764 500880 62816 500886
rect 62764 500822 62816 500828
rect 70032 500880 70084 500886
rect 70032 500822 70084 500828
rect 79704 500818 79732 502044
rect 90376 500818 90404 523058
rect 90468 505646 90496 523126
rect 106384 521914 106412 523126
rect 115940 523116 115992 523122
rect 115940 523058 115992 523064
rect 115952 521914 115980 523058
rect 106384 521886 106674 521914
rect 115952 521886 116334 521914
rect 96724 521206 97014 521234
rect 91100 520396 91152 520402
rect 91100 520338 91152 520344
rect 91112 511737 91140 520338
rect 91098 511728 91154 511737
rect 91098 511663 91154 511672
rect 90456 505640 90508 505646
rect 90456 505582 90508 505588
rect 96724 500954 96752 521206
rect 96896 520328 96948 520334
rect 96896 520270 96948 520276
rect 96908 512961 96936 520270
rect 96894 512952 96950 512961
rect 96894 512887 96950 512896
rect 96712 500948 96764 500954
rect 96712 500890 96764 500896
rect 97000 500886 97028 502044
rect 96988 500880 97040 500886
rect 96988 500822 97040 500828
rect 106660 500818 106688 502044
rect 116320 501922 116348 502044
rect 116504 501922 116532 523126
rect 116584 523116 116636 523122
rect 116584 523058 116636 523064
rect 116320 501894 116532 501922
rect 116596 500818 116624 523058
rect 133432 521914 133460 523126
rect 142988 523116 143040 523122
rect 142988 523058 143040 523064
rect 143000 521914 143028 523058
rect 133432 521886 133722 521914
rect 143000 521886 143382 521914
rect 122944 521206 124062 521234
rect 118700 520464 118752 520470
rect 118700 520406 118752 520412
rect 118712 511737 118740 520406
rect 122748 520396 122800 520402
rect 122748 520338 122800 520344
rect 122760 512417 122788 520338
rect 122746 512408 122802 512417
rect 122746 512343 122802 512352
rect 118698 511728 118754 511737
rect 118698 511663 118754 511672
rect 122944 500818 122972 521206
rect 144196 509234 144224 523126
rect 144276 523116 144328 523122
rect 144276 523058 144328 523064
rect 143736 509206 144224 509234
rect 143736 502738 143764 509206
rect 143382 502710 143764 502738
rect 124048 500886 124076 502044
rect 133708 500886 133736 502044
rect 144288 500886 144316 523058
rect 146300 520328 146352 520334
rect 146300 520270 146352 520276
rect 146312 512009 146340 520270
rect 146298 512000 146354 512009
rect 146298 511935 146354 511944
rect 146956 500954 146984 550870
rect 148966 539200 149022 539209
rect 148966 539135 149022 539144
rect 148980 529922 149008 539135
rect 148968 529916 149020 529922
rect 148968 529858 149020 529864
rect 149716 527066 149744 578478
rect 232320 578468 232372 578474
rect 232320 578410 232372 578416
rect 251824 578468 251876 578474
rect 251824 578410 251876 578416
rect 475384 578468 475436 578474
rect 475384 578410 475436 578416
rect 494704 578468 494756 578474
rect 494704 578410 494756 578416
rect 160284 578400 160336 578406
rect 160284 578342 160336 578348
rect 170496 578400 170548 578406
rect 170496 578342 170548 578348
rect 187792 578400 187844 578406
rect 187792 578342 187844 578348
rect 197544 578400 197596 578406
rect 197544 578342 197596 578348
rect 214380 578400 214432 578406
rect 214380 578342 214432 578348
rect 224500 578400 224552 578406
rect 224500 578342 224552 578348
rect 160296 575906 160324 578342
rect 170036 578332 170088 578338
rect 170036 578274 170088 578280
rect 170048 575906 170076 578274
rect 160296 575878 160678 575906
rect 170048 575878 170338 575906
rect 150544 575334 151018 575362
rect 150544 554674 150572 575334
rect 150532 554668 150584 554674
rect 150532 554610 150584 554616
rect 151004 554606 151032 556036
rect 150992 554600 151044 554606
rect 150992 554542 151044 554548
rect 160664 554538 160692 556036
rect 170324 555914 170352 556036
rect 170508 555914 170536 578342
rect 178408 578332 178460 578338
rect 178408 578274 178460 578280
rect 171784 578264 171836 578270
rect 171784 578206 171836 578212
rect 170324 555886 170536 555914
rect 171796 554538 171824 578206
rect 178420 575906 178448 578274
rect 187804 575906 187832 578342
rect 197452 578264 197504 578270
rect 197452 578206 197504 578212
rect 197464 575906 197492 578206
rect 178066 575878 178448 575906
rect 187726 575878 187832 575906
rect 197386 575878 197492 575906
rect 197556 567194 197584 578342
rect 200764 578332 200816 578338
rect 200764 578274 200816 578280
rect 199384 578264 199436 578270
rect 199384 578206 199436 578212
rect 197464 567166 197584 567194
rect 176566 565856 176622 565865
rect 176566 565791 176622 565800
rect 172518 565584 172574 565593
rect 172518 565519 172574 565528
rect 172532 557462 172560 565519
rect 176580 557462 176608 565791
rect 172520 557456 172572 557462
rect 172520 557398 172572 557404
rect 176568 557456 176620 557462
rect 176568 557398 176620 557404
rect 197464 556730 197492 567166
rect 197386 556702 197492 556730
rect 178052 554606 178080 556036
rect 187712 554606 187740 556036
rect 199396 554606 199424 578206
rect 200118 565584 200174 565593
rect 200118 565519 200174 565528
rect 200132 557530 200160 565519
rect 200120 557524 200172 557530
rect 200120 557466 200172 557472
rect 200776 554742 200804 578274
rect 214392 575906 214420 578342
rect 223948 578264 224000 578270
rect 223948 578206 224000 578212
rect 223960 575906 223988 578206
rect 214392 575878 214682 575906
rect 223960 575878 224342 575906
rect 204364 575334 205022 575362
rect 202786 566264 202842 566273
rect 202786 566199 202842 566208
rect 202800 557530 202828 566199
rect 202788 557524 202840 557530
rect 202788 557466 202840 557472
rect 200764 554736 200816 554742
rect 200764 554678 200816 554684
rect 204364 554606 204392 575334
rect 224512 556730 224540 578342
rect 225604 578264 225656 578270
rect 225604 578206 225656 578212
rect 224342 556702 224540 556730
rect 205008 554742 205036 556036
rect 204996 554736 205048 554742
rect 204996 554678 205048 554684
rect 178040 554600 178092 554606
rect 178040 554542 178092 554548
rect 187700 554600 187752 554606
rect 187700 554542 187752 554548
rect 199384 554600 199436 554606
rect 199384 554542 199436 554548
rect 204352 554600 204404 554606
rect 204352 554542 204404 554548
rect 214668 554538 214696 556036
rect 225616 554538 225644 578206
rect 232332 575906 232360 578410
rect 241612 578400 241664 578406
rect 241612 578342 241664 578348
rect 232070 575878 232360 575906
rect 241624 575906 241652 578342
rect 251456 578332 251508 578338
rect 251456 578274 251508 578280
rect 251272 578264 251324 578270
rect 251272 578206 251324 578212
rect 251284 575906 251312 578206
rect 241624 575878 241730 575906
rect 251284 575878 251390 575906
rect 230386 566264 230442 566273
rect 230386 566199 230442 566208
rect 226338 565584 226394 565593
rect 226338 565519 226394 565528
rect 226352 557462 226380 565519
rect 230400 557462 230428 566199
rect 226340 557456 226392 557462
rect 226340 557398 226392 557404
rect 230388 557456 230440 557462
rect 230388 557398 230440 557404
rect 251468 556730 251496 578274
rect 251390 556702 251496 556730
rect 232056 554606 232084 556036
rect 241716 554606 241744 556036
rect 251836 554742 251864 578410
rect 413468 578400 413520 578406
rect 413468 578342 413520 578348
rect 430580 578400 430632 578406
rect 430580 578342 430632 578348
rect 440516 578400 440568 578406
rect 440516 578342 440568 578348
rect 457260 578400 457312 578406
rect 457260 578342 457312 578348
rect 468484 578400 468536 578406
rect 468484 578342 468536 578348
rect 268292 578332 268344 578338
rect 268292 578274 268344 578280
rect 279424 578332 279476 578338
rect 279424 578274 279476 578280
rect 295800 578332 295852 578338
rect 295800 578274 295852 578280
rect 305552 578332 305604 578338
rect 305552 578274 305604 578280
rect 322388 578332 322440 578338
rect 322388 578274 322440 578280
rect 336004 578332 336056 578338
rect 336004 578274 336056 578280
rect 349804 578332 349856 578338
rect 349804 578274 349856 578280
rect 359648 578332 359700 578338
rect 359648 578274 359700 578280
rect 376300 578332 376352 578338
rect 376300 578274 376352 578280
rect 386512 578332 386564 578338
rect 386512 578274 386564 578280
rect 403348 578332 403400 578338
rect 403348 578274 403400 578280
rect 253204 578264 253256 578270
rect 253204 578206 253256 578212
rect 251824 554736 251876 554742
rect 251824 554678 251876 554684
rect 253216 554606 253244 578206
rect 268304 575906 268332 578274
rect 278044 578264 278096 578270
rect 278044 578206 278096 578212
rect 278056 575906 278084 578206
rect 268304 575878 268686 575906
rect 278056 575878 278346 575906
rect 258184 575334 259026 575362
rect 256606 566264 256662 566273
rect 256606 566199 256662 566208
rect 253938 565040 253994 565049
rect 253938 564975 253994 564984
rect 253952 557530 253980 564975
rect 256620 557530 256648 566199
rect 253940 557524 253992 557530
rect 253940 557466 253992 557472
rect 256608 557524 256660 557530
rect 256608 557466 256660 557472
rect 258184 554606 258212 575334
rect 279436 557534 279464 578274
rect 279516 578264 279568 578270
rect 279516 578206 279568 578212
rect 278792 557506 279464 557534
rect 278792 556730 278820 557506
rect 278346 556702 278820 556730
rect 259012 554742 259040 556036
rect 259000 554736 259052 554742
rect 259000 554678 259052 554684
rect 232044 554600 232096 554606
rect 232044 554542 232096 554548
rect 241704 554600 241756 554606
rect 241704 554542 241756 554548
rect 253204 554600 253256 554606
rect 253204 554542 253256 554548
rect 258172 554600 258224 554606
rect 258172 554542 258224 554548
rect 268672 554538 268700 556036
rect 279528 554538 279556 578206
rect 295812 575906 295840 578274
rect 305460 578264 305512 578270
rect 305460 578206 305512 578212
rect 305472 575906 305500 578206
rect 295734 575878 295840 575906
rect 305394 575878 305500 575906
rect 286074 575470 286180 575498
rect 286152 575414 286180 575470
rect 285772 575408 285824 575414
rect 285772 575350 285824 575356
rect 286140 575408 286192 575414
rect 286140 575350 286192 575356
rect 284206 565856 284262 565865
rect 284206 565791 284262 565800
rect 280158 565584 280214 565593
rect 280158 565519 280214 565528
rect 280172 557462 280200 565519
rect 284220 557462 284248 565791
rect 280160 557456 280212 557462
rect 280160 557398 280212 557404
rect 284208 557456 284260 557462
rect 284208 557398 284260 557404
rect 285784 554538 285812 575350
rect 305564 567194 305592 578274
rect 307024 578264 307076 578270
rect 307024 578206 307076 578212
rect 305472 567166 305592 567194
rect 305472 556730 305500 567166
rect 305394 556702 305500 556730
rect 286060 554606 286088 556036
rect 286048 554600 286100 554606
rect 286048 554542 286100 554548
rect 295720 554538 295748 556036
rect 307036 554538 307064 578206
rect 322400 575906 322428 578274
rect 331956 578264 332008 578270
rect 331956 578206 332008 578212
rect 333244 578264 333296 578270
rect 333244 578206 333296 578212
rect 331968 575906 331996 578206
rect 322400 575878 322690 575906
rect 331968 575878 332350 575906
rect 312004 575334 313030 575362
rect 311806 566264 311862 566273
rect 311806 566199 311862 566208
rect 307758 565584 307814 565593
rect 307758 565519 307814 565528
rect 307772 557530 307800 565519
rect 307760 557524 307812 557530
rect 307760 557466 307812 557472
rect 311820 557394 311848 566199
rect 311808 557388 311860 557394
rect 311808 557330 311860 557336
rect 312004 554538 312032 575334
rect 313016 554606 313044 556036
rect 313004 554600 313056 554606
rect 313004 554542 313056 554548
rect 322676 554538 322704 556036
rect 332336 554742 332364 556036
rect 332324 554736 332376 554742
rect 332324 554678 332376 554684
rect 333256 554538 333284 578206
rect 335358 565584 335414 565593
rect 335358 565519 335414 565528
rect 335372 557462 335400 565519
rect 335360 557456 335412 557462
rect 335360 557398 335412 557404
rect 336016 554742 336044 578274
rect 349816 575906 349844 578274
rect 359464 578264 359516 578270
rect 359464 578206 359516 578212
rect 359476 575906 359504 578206
rect 349738 575878 349844 575906
rect 359398 575878 359504 575906
rect 340078 575346 340184 575362
rect 339592 575340 339644 575346
rect 340078 575340 340196 575346
rect 340078 575334 340144 575340
rect 339592 575282 339644 575288
rect 340144 575282 340196 575288
rect 338026 566264 338082 566273
rect 338026 566199 338082 566208
rect 338040 557530 338068 566199
rect 338028 557524 338080 557530
rect 338028 557466 338080 557472
rect 336004 554736 336056 554742
rect 336004 554678 336056 554684
rect 339604 554538 339632 575282
rect 359660 570466 359688 578274
rect 359740 578264 359792 578270
rect 359740 578206 359792 578212
rect 359476 570438 359688 570466
rect 359476 556730 359504 570438
rect 359752 567202 359780 578206
rect 376312 575906 376340 578274
rect 386052 578264 386104 578270
rect 386052 578206 386104 578212
rect 386064 575906 386092 578206
rect 376312 575878 376694 575906
rect 386064 575878 386354 575906
rect 359398 556702 359504 556730
rect 359568 567174 359780 567202
rect 365824 575334 367034 575362
rect 340064 554606 340092 556036
rect 340052 554600 340104 554606
rect 340052 554542 340104 554548
rect 349724 554538 349752 556036
rect 359568 554538 359596 567174
rect 365626 566264 365682 566273
rect 365626 566199 365682 566208
rect 361578 565040 361634 565049
rect 361578 564975 361634 564984
rect 361592 557394 361620 564975
rect 365640 557462 365668 566199
rect 365628 557456 365680 557462
rect 365628 557398 365680 557404
rect 361580 557388 361632 557394
rect 361580 557330 361632 557336
rect 365824 554538 365852 575334
rect 386524 556730 386552 578274
rect 387064 578264 387116 578270
rect 387064 578206 387116 578212
rect 386354 556702 386552 556730
rect 367020 554606 367048 556036
rect 367008 554600 367060 554606
rect 367008 554542 367060 554548
rect 376680 554538 376708 556036
rect 387076 554538 387104 578206
rect 403360 575906 403388 578274
rect 412916 578264 412968 578270
rect 412916 578206 412968 578212
rect 412928 575906 412956 578206
rect 403360 575878 403650 575906
rect 412928 575878 413310 575906
rect 393424 575334 393990 575362
rect 391846 566264 391902 566273
rect 391846 566199 391902 566208
rect 389178 565584 389234 565593
rect 389178 565519 389234 565528
rect 389192 557530 389220 565519
rect 391860 557530 391888 566199
rect 389180 557524 389232 557530
rect 389180 557466 389232 557472
rect 391848 557524 391900 557530
rect 391848 557466 391900 557472
rect 393424 554538 393452 575334
rect 413480 556730 413508 578342
rect 421288 578332 421340 578338
rect 421288 578274 421340 578280
rect 414664 578264 414716 578270
rect 414664 578206 414716 578212
rect 413402 556702 413508 556730
rect 393976 554606 394004 556036
rect 393964 554600 394016 554606
rect 393964 554542 394016 554548
rect 403728 554538 403756 556036
rect 414676 554538 414704 578206
rect 421300 575906 421328 578274
rect 421038 575878 421328 575906
rect 430592 575906 430620 578342
rect 440240 578264 440292 578270
rect 440240 578206 440292 578212
rect 440252 575906 440280 578206
rect 430592 575878 430698 575906
rect 440252 575878 440358 575906
rect 419446 566264 419502 566273
rect 419446 566199 419502 566208
rect 415398 565584 415454 565593
rect 415398 565519 415454 565528
rect 415412 557462 415440 565519
rect 419460 557462 419488 566199
rect 415400 557456 415452 557462
rect 415400 557398 415452 557404
rect 419448 557456 419500 557462
rect 419448 557398 419500 557404
rect 440528 556730 440556 578342
rect 446404 578332 446456 578338
rect 446404 578274 446456 578280
rect 442264 578264 442316 578270
rect 442264 578206 442316 578212
rect 440358 556702 440556 556730
rect 421024 554606 421052 556036
rect 430684 554606 430712 556036
rect 442276 554606 442304 578206
rect 445666 566264 445722 566273
rect 445666 566199 445722 566208
rect 442998 565584 443054 565593
rect 442998 565519 443054 565528
rect 443012 557530 443040 565519
rect 445680 557530 445708 566199
rect 443000 557524 443052 557530
rect 443000 557466 443052 557472
rect 445668 557524 445720 557530
rect 445668 557466 445720 557472
rect 446416 556782 446444 578274
rect 457272 575906 457300 578342
rect 467012 578264 467064 578270
rect 467012 578206 467064 578212
rect 467024 575906 467052 578206
rect 457272 575878 457654 575906
rect 467024 575878 467314 575906
rect 447244 575334 447994 575362
rect 446404 556776 446456 556782
rect 446404 556718 446456 556724
rect 447244 554606 447272 575334
rect 468496 557534 468524 578342
rect 468576 578264 468628 578270
rect 468576 578206 468628 578212
rect 467760 557506 468524 557534
rect 447692 556776 447744 556782
rect 467760 556730 467788 557506
rect 447744 556724 447994 556730
rect 447692 556718 447994 556724
rect 447704 556702 447994 556718
rect 467406 556702 467788 556730
rect 421012 554600 421064 554606
rect 421012 554542 421064 554548
rect 430672 554600 430724 554606
rect 430672 554542 430724 554548
rect 442264 554600 442316 554606
rect 442264 554542 442316 554548
rect 447232 554600 447284 554606
rect 447232 554542 447284 554548
rect 457732 554538 457760 556036
rect 468588 554538 468616 578206
rect 475396 575906 475424 578410
rect 484400 578400 484452 578406
rect 484400 578342 484452 578348
rect 475042 575878 475424 575906
rect 484412 575906 484440 578342
rect 494520 578332 494572 578338
rect 494520 578274 494572 578280
rect 494060 578264 494112 578270
rect 494060 578206 494112 578212
rect 494072 575906 494100 578206
rect 484412 575878 484702 575906
rect 494072 575878 494362 575906
rect 473266 565856 473322 565865
rect 473266 565791 473322 565800
rect 469218 565040 469274 565049
rect 469218 564975 469274 564984
rect 469232 557462 469260 564975
rect 473280 557462 473308 565791
rect 469220 557456 469272 557462
rect 469220 557398 469272 557404
rect 473268 557456 473320 557462
rect 473268 557398 473320 557404
rect 494532 556730 494560 578274
rect 494362 556702 494560 556730
rect 475028 554606 475056 556036
rect 484688 554606 484716 556036
rect 494716 554742 494744 578410
rect 511356 578332 511408 578338
rect 511356 578274 511408 578280
rect 522396 578332 522448 578338
rect 522396 578274 522448 578280
rect 496084 578264 496136 578270
rect 496084 578206 496136 578212
rect 494704 554736 494756 554742
rect 494704 554678 494756 554684
rect 496096 554606 496124 578206
rect 511368 575906 511396 578274
rect 520924 578264 520976 578270
rect 520924 578206 520976 578212
rect 522304 578264 522356 578270
rect 522304 578206 522356 578212
rect 520936 575906 520964 578206
rect 511368 575878 511658 575906
rect 520936 575878 521318 575906
rect 501064 575334 501998 575362
rect 500866 566264 500922 566273
rect 500866 566199 500922 566208
rect 496818 565584 496874 565593
rect 496818 565519 496874 565528
rect 496832 557530 496860 565519
rect 500880 557530 500908 566199
rect 496820 557524 496872 557530
rect 496820 557466 496872 557472
rect 500868 557524 500920 557530
rect 500868 557466 500920 557472
rect 501064 554606 501092 575334
rect 521752 556776 521804 556782
rect 521410 556724 521752 556730
rect 521410 556718 521804 556724
rect 521410 556702 521792 556718
rect 501984 554742 502012 556036
rect 501972 554736 502024 554742
rect 501972 554678 502024 554684
rect 475016 554600 475068 554606
rect 475016 554542 475068 554548
rect 484676 554600 484728 554606
rect 484676 554542 484728 554548
rect 496084 554600 496136 554606
rect 496084 554542 496136 554548
rect 501052 554600 501104 554606
rect 501052 554542 501104 554548
rect 511736 554538 511764 556036
rect 522316 554538 522344 578206
rect 522408 556782 522436 578274
rect 526444 576156 526496 576162
rect 526444 576098 526496 576104
rect 526456 566409 526484 576098
rect 526442 566400 526498 566409
rect 526442 566335 526498 566344
rect 523038 565584 523094 565593
rect 523038 565519 523094 565528
rect 523052 557462 523080 565519
rect 523040 557456 523092 557462
rect 523040 557398 523092 557404
rect 522396 556776 522448 556782
rect 522396 556718 522448 556724
rect 160652 554532 160704 554538
rect 160652 554474 160704 554480
rect 171784 554532 171836 554538
rect 171784 554474 171836 554480
rect 214656 554532 214708 554538
rect 214656 554474 214708 554480
rect 225604 554532 225656 554538
rect 225604 554474 225656 554480
rect 268660 554532 268712 554538
rect 268660 554474 268712 554480
rect 279516 554532 279568 554538
rect 279516 554474 279568 554480
rect 285772 554532 285824 554538
rect 285772 554474 285824 554480
rect 295708 554532 295760 554538
rect 295708 554474 295760 554480
rect 307024 554532 307076 554538
rect 307024 554474 307076 554480
rect 311992 554532 312044 554538
rect 311992 554474 312044 554480
rect 322664 554532 322716 554538
rect 322664 554474 322716 554480
rect 333244 554532 333296 554538
rect 333244 554474 333296 554480
rect 339592 554532 339644 554538
rect 339592 554474 339644 554480
rect 349712 554532 349764 554538
rect 349712 554474 349764 554480
rect 359556 554532 359608 554538
rect 359556 554474 359608 554480
rect 365812 554532 365864 554538
rect 365812 554474 365864 554480
rect 376668 554532 376720 554538
rect 376668 554474 376720 554480
rect 387064 554532 387116 554538
rect 387064 554474 387116 554480
rect 393412 554532 393464 554538
rect 393412 554474 393464 554480
rect 403716 554532 403768 554538
rect 403716 554474 403768 554480
rect 414664 554532 414716 554538
rect 414664 554474 414716 554480
rect 457720 554532 457772 554538
rect 457720 554474 457772 554480
rect 468576 554532 468628 554538
rect 468576 554474 468628 554480
rect 511724 554532 511776 554538
rect 511724 554474 511776 554480
rect 522304 554532 522356 554538
rect 522304 554474 522356 554480
rect 232044 550860 232096 550866
rect 232044 550802 232096 550808
rect 251824 550860 251876 550866
rect 251824 550802 251876 550808
rect 475016 550860 475068 550866
rect 475016 550802 475068 550808
rect 494704 550860 494756 550866
rect 494704 550802 494756 550808
rect 170496 550792 170548 550798
rect 170496 550734 170548 550740
rect 187700 550792 187752 550798
rect 187700 550734 187752 550740
rect 197452 550792 197504 550798
rect 197452 550734 197504 550740
rect 214656 550792 214708 550798
rect 214656 550734 214708 550740
rect 224500 550792 224552 550798
rect 224500 550734 224552 550740
rect 170312 550724 170364 550730
rect 170312 550666 170364 550672
rect 160652 550656 160704 550662
rect 160652 550598 160704 550604
rect 160664 548964 160692 550598
rect 170324 548964 170352 550666
rect 150544 548270 151018 548298
rect 149704 527060 149756 527066
rect 149704 527002 149756 527008
rect 150544 526998 150572 548270
rect 170232 529650 170338 529666
rect 170508 529650 170536 550734
rect 178040 550724 178092 550730
rect 178040 550666 178092 550672
rect 171784 550656 171836 550662
rect 171784 550598 171836 550604
rect 170220 529644 170338 529650
rect 170272 529638 170338 529644
rect 170496 529644 170548 529650
rect 170220 529586 170272 529592
rect 170496 529586 170548 529592
rect 150728 529094 151018 529122
rect 160572 529094 160678 529122
rect 150532 526992 150584 526998
rect 150532 526934 150584 526940
rect 150728 526930 150756 529094
rect 160572 526930 160600 529094
rect 171796 526930 171824 550598
rect 178052 548964 178080 550666
rect 187712 548964 187740 550734
rect 197360 550656 197412 550662
rect 197360 550598 197412 550604
rect 197372 548964 197400 550598
rect 176566 538656 176622 538665
rect 176566 538591 176622 538600
rect 172518 538520 172574 538529
rect 172518 538455 172574 538464
rect 172532 529854 172560 538455
rect 176580 529854 176608 538591
rect 172520 529848 172572 529854
rect 172520 529790 172572 529796
rect 176568 529848 176620 529854
rect 176568 529790 176620 529796
rect 197464 529666 197492 550734
rect 200764 550724 200816 550730
rect 200764 550666 200816 550672
rect 199384 550656 199436 550662
rect 199384 550598 199436 550604
rect 197386 529638 197492 529666
rect 178066 529094 178172 529122
rect 187726 529094 188016 529122
rect 178144 526998 178172 529094
rect 187988 526998 188016 529094
rect 199396 526998 199424 550598
rect 200118 538520 200174 538529
rect 200118 538455 200174 538464
rect 200132 529922 200160 538455
rect 200120 529916 200172 529922
rect 200120 529858 200172 529864
rect 200776 527134 200804 550666
rect 214668 548964 214696 550734
rect 224316 550656 224368 550662
rect 224316 550598 224368 550604
rect 224328 548964 224356 550598
rect 204364 548270 205022 548298
rect 202786 539200 202842 539209
rect 202786 539135 202842 539144
rect 202800 529922 202828 539135
rect 202788 529916 202840 529922
rect 202788 529858 202840 529864
rect 200764 527128 200816 527134
rect 200764 527070 200816 527076
rect 204364 526998 204392 548270
rect 224512 529666 224540 550734
rect 225604 550656 225656 550662
rect 225604 550598 225656 550604
rect 224342 529638 224540 529666
rect 204640 529094 205022 529122
rect 214682 529094 215064 529122
rect 204640 527134 204668 529094
rect 204628 527128 204680 527134
rect 204628 527070 204680 527076
rect 178132 526992 178184 526998
rect 178132 526934 178184 526940
rect 187976 526992 188028 526998
rect 187976 526934 188028 526940
rect 199384 526992 199436 526998
rect 199384 526934 199436 526940
rect 204352 526992 204404 526998
rect 204352 526934 204404 526940
rect 215036 526930 215064 529094
rect 225616 526930 225644 550598
rect 232056 548964 232084 550802
rect 241704 550792 241756 550798
rect 241704 550734 241756 550740
rect 241716 548964 241744 550734
rect 251456 550724 251508 550730
rect 251456 550666 251508 550672
rect 251364 550656 251416 550662
rect 251364 550598 251416 550604
rect 251376 548964 251404 550598
rect 230386 539200 230442 539209
rect 230386 539135 230442 539144
rect 226338 538520 226394 538529
rect 226338 538455 226394 538464
rect 226352 529854 226380 538455
rect 230400 529854 230428 539135
rect 226340 529848 226392 529854
rect 226340 529790 226392 529796
rect 230388 529848 230440 529854
rect 230388 529790 230440 529796
rect 251468 529666 251496 550666
rect 251390 529638 251496 529666
rect 231964 529094 232070 529122
rect 241730 529094 242112 529122
rect 231964 526998 231992 529094
rect 242084 526998 242112 529094
rect 251836 527134 251864 550802
rect 413468 550792 413520 550798
rect 413468 550734 413520 550740
rect 430672 550792 430724 550798
rect 430672 550734 430724 550740
rect 440516 550792 440568 550798
rect 440516 550734 440568 550740
rect 457628 550792 457680 550798
rect 457628 550734 457680 550740
rect 468484 550792 468536 550798
rect 468484 550734 468536 550740
rect 268660 550724 268712 550730
rect 268660 550666 268712 550672
rect 279516 550724 279568 550730
rect 279516 550666 279568 550672
rect 295708 550724 295760 550730
rect 295708 550666 295760 550672
rect 305460 550724 305512 550730
rect 305460 550666 305512 550672
rect 322664 550724 322716 550730
rect 322664 550666 322716 550672
rect 334624 550724 334676 550730
rect 334624 550666 334676 550672
rect 349712 550724 349764 550730
rect 349712 550666 349764 550672
rect 359464 550724 359516 550730
rect 359464 550666 359516 550672
rect 376668 550724 376720 550730
rect 376668 550666 376720 550672
rect 386512 550724 386564 550730
rect 386512 550666 386564 550672
rect 403624 550724 403676 550730
rect 403624 550666 403676 550672
rect 253204 550656 253256 550662
rect 253204 550598 253256 550604
rect 251824 527128 251876 527134
rect 251824 527070 251876 527076
rect 253216 526998 253244 550598
rect 268672 548964 268700 550666
rect 278320 550656 278372 550662
rect 278320 550598 278372 550604
rect 279424 550656 279476 550662
rect 279424 550598 279476 550604
rect 278332 548964 278360 550598
rect 258184 548270 259026 548298
rect 256606 539200 256662 539209
rect 256606 539135 256662 539144
rect 253938 538384 253994 538393
rect 253938 538319 253994 538328
rect 253952 529922 253980 538319
rect 256620 529922 256648 539135
rect 253940 529916 253992 529922
rect 253940 529858 253992 529864
rect 256608 529916 256660 529922
rect 256608 529858 256660 529864
rect 258184 526998 258212 548270
rect 278688 529848 278740 529854
rect 278688 529790 278740 529796
rect 278700 529666 278728 529790
rect 278346 529638 278728 529666
rect 258736 529094 259026 529122
rect 268686 529094 268976 529122
rect 258736 527134 258764 529094
rect 258724 527128 258776 527134
rect 258724 527070 258776 527076
rect 231952 526992 232004 526998
rect 231952 526934 232004 526940
rect 242072 526992 242124 526998
rect 242072 526934 242124 526940
rect 253204 526992 253256 526998
rect 253204 526934 253256 526940
rect 258172 526992 258224 526998
rect 258172 526934 258224 526940
rect 268948 526930 268976 529094
rect 279436 526930 279464 550598
rect 279528 529854 279556 550666
rect 285784 549086 286088 549114
rect 284206 538656 284262 538665
rect 284206 538591 284262 538600
rect 280158 538520 280214 538529
rect 280158 538455 280214 538464
rect 279516 529848 279568 529854
rect 279516 529790 279568 529796
rect 280172 529786 280200 538455
rect 284220 529854 284248 538591
rect 284208 529848 284260 529854
rect 284208 529790 284260 529796
rect 280160 529780 280212 529786
rect 280160 529722 280212 529728
rect 285784 526998 285812 549086
rect 286060 548964 286088 549086
rect 295720 548964 295748 550666
rect 305368 550656 305420 550662
rect 305368 550598 305420 550604
rect 305380 548964 305408 550598
rect 305472 529666 305500 550666
rect 307024 550656 307076 550662
rect 307024 550598 307076 550604
rect 305394 529638 305500 529666
rect 286074 529094 286180 529122
rect 295734 529094 296024 529122
rect 285772 526992 285824 526998
rect 285772 526934 285824 526940
rect 286152 526930 286180 529094
rect 295996 526930 296024 529094
rect 307036 526930 307064 550598
rect 322676 548964 322704 550666
rect 332324 550656 332376 550662
rect 332324 550598 332376 550604
rect 333244 550656 333296 550662
rect 333244 550598 333296 550604
rect 332336 548964 332364 550598
rect 312004 548270 313030 548298
rect 311806 539200 311862 539209
rect 311806 539135 311862 539144
rect 307758 538520 307814 538529
rect 307758 538455 307814 538464
rect 307772 529922 307800 538455
rect 307760 529916 307812 529922
rect 307760 529858 307812 529864
rect 311820 529786 311848 539135
rect 311808 529780 311860 529786
rect 311808 529722 311860 529728
rect 312004 526930 312032 548270
rect 332508 529916 332560 529922
rect 332508 529858 332560 529864
rect 332520 529666 332548 529858
rect 332350 529638 332548 529666
rect 312648 529094 313030 529122
rect 322690 529094 322888 529122
rect 312648 526998 312676 529094
rect 312636 526992 312688 526998
rect 312636 526934 312688 526940
rect 322860 526930 322888 529094
rect 333256 526930 333284 550598
rect 334636 529922 334664 550666
rect 339604 549086 340092 549114
rect 338026 539200 338082 539209
rect 338026 539135 338082 539144
rect 335358 538520 335414 538529
rect 335358 538455 335414 538464
rect 334624 529916 334676 529922
rect 334624 529858 334676 529864
rect 335372 529854 335400 538455
rect 338040 529922 338068 539135
rect 338028 529916 338080 529922
rect 338028 529858 338080 529864
rect 335360 529848 335412 529854
rect 335360 529790 335412 529796
rect 339604 526930 339632 549086
rect 340064 548964 340092 549086
rect 349724 548964 349752 550666
rect 359372 550656 359424 550662
rect 359372 550598 359424 550604
rect 359384 548964 359412 550598
rect 359476 529666 359504 550666
rect 359556 550656 359608 550662
rect 359556 550598 359608 550604
rect 359398 529638 359504 529666
rect 340078 529094 340184 529122
rect 349738 529094 350120 529122
rect 340156 526998 340184 529094
rect 340144 526992 340196 526998
rect 340144 526934 340196 526940
rect 350092 526930 350120 529094
rect 359568 526930 359596 550598
rect 376680 548964 376708 550666
rect 386328 550656 386380 550662
rect 386328 550598 386380 550604
rect 386340 548964 386368 550598
rect 365824 548270 367034 548298
rect 365626 539200 365682 539209
rect 365626 539135 365682 539144
rect 361578 538384 361634 538393
rect 361578 538319 361634 538328
rect 361592 529786 361620 538319
rect 365640 529854 365668 539135
rect 365628 529848 365680 529854
rect 365628 529790 365680 529796
rect 361580 529780 361632 529786
rect 361580 529722 361632 529728
rect 365824 526930 365852 548270
rect 386524 529666 386552 550666
rect 387064 550656 387116 550662
rect 387064 550598 387116 550604
rect 386354 529638 386552 529666
rect 366744 529094 367034 529122
rect 376588 529094 376694 529122
rect 366744 526998 366772 529094
rect 366732 526992 366784 526998
rect 366732 526934 366784 526940
rect 376588 526930 376616 529094
rect 387076 526930 387104 550598
rect 403636 548964 403664 550666
rect 413284 550656 413336 550662
rect 413284 550598 413336 550604
rect 413296 548964 413324 550598
rect 393424 548270 393990 548298
rect 391846 539200 391902 539209
rect 391846 539135 391902 539144
rect 389178 538520 389234 538529
rect 389178 538455 389234 538464
rect 389192 529922 389220 538455
rect 391860 529922 391888 539135
rect 389180 529916 389232 529922
rect 389180 529858 389232 529864
rect 391848 529916 391900 529922
rect 391848 529858 391900 529864
rect 393424 526930 393452 548270
rect 413480 529666 413508 550734
rect 421012 550724 421064 550730
rect 421012 550666 421064 550672
rect 414664 550656 414716 550662
rect 414664 550598 414716 550604
rect 413402 529638 413508 529666
rect 393608 529094 393990 529122
rect 403742 529094 404032 529122
rect 393608 526998 393636 529094
rect 393596 526992 393648 526998
rect 393596 526934 393648 526940
rect 404004 526930 404032 529094
rect 414676 526930 414704 550598
rect 421024 548964 421052 550666
rect 430684 548964 430712 550734
rect 440332 550656 440384 550662
rect 440332 550598 440384 550604
rect 440344 548964 440372 550598
rect 419446 539200 419502 539209
rect 419446 539135 419502 539144
rect 415398 538520 415454 538529
rect 415398 538455 415454 538464
rect 415412 529854 415440 538455
rect 419460 529854 419488 539135
rect 415400 529848 415452 529854
rect 415400 529790 415452 529796
rect 419448 529848 419500 529854
rect 419448 529790 419500 529796
rect 440528 529666 440556 550734
rect 443644 550724 443696 550730
rect 443644 550666 443696 550672
rect 442264 550656 442316 550662
rect 442264 550598 442316 550604
rect 440358 529638 440556 529666
rect 420932 529094 421038 529122
rect 430698 529094 431080 529122
rect 420932 526998 420960 529094
rect 431052 526998 431080 529094
rect 442276 526998 442304 550598
rect 442998 538520 443054 538529
rect 442998 538455 443054 538464
rect 443012 529922 443040 538455
rect 443000 529916 443052 529922
rect 443000 529858 443052 529864
rect 443656 527134 443684 550666
rect 457640 548964 457668 550734
rect 467288 550656 467340 550662
rect 467288 550598 467340 550604
rect 467300 548964 467328 550598
rect 447244 548270 447994 548298
rect 445666 539200 445722 539209
rect 445666 539135 445722 539144
rect 445680 529922 445708 539135
rect 445668 529916 445720 529922
rect 445668 529858 445720 529864
rect 443644 527128 443696 527134
rect 443644 527070 443696 527076
rect 447244 526998 447272 548270
rect 468496 538214 468524 550734
rect 468576 550656 468628 550662
rect 468576 550598 468628 550604
rect 467852 538186 468524 538214
rect 467852 529666 467880 538186
rect 467406 529638 467880 529666
rect 447704 529094 447994 529122
rect 457746 529094 458128 529122
rect 447704 527134 447732 529094
rect 447692 527128 447744 527134
rect 447692 527070 447744 527076
rect 420920 526992 420972 526998
rect 420920 526934 420972 526940
rect 431040 526992 431092 526998
rect 431040 526934 431092 526940
rect 442264 526992 442316 526998
rect 442264 526934 442316 526940
rect 447232 526992 447284 526998
rect 447232 526934 447284 526940
rect 458100 526930 458128 529094
rect 468588 526930 468616 550598
rect 475028 548964 475056 550802
rect 484676 550792 484728 550798
rect 484676 550734 484728 550740
rect 484688 548964 484716 550734
rect 494520 550724 494572 550730
rect 494520 550666 494572 550672
rect 494336 550656 494388 550662
rect 494336 550598 494388 550604
rect 494348 548964 494376 550598
rect 473266 538656 473322 538665
rect 473266 538591 473322 538600
rect 469218 538384 469274 538393
rect 469218 538319 469274 538328
rect 469232 529854 469260 538319
rect 473280 529854 473308 538591
rect 469220 529848 469272 529854
rect 469220 529790 469272 529796
rect 473268 529848 473320 529854
rect 473268 529790 473320 529796
rect 494532 529666 494560 550666
rect 494362 529638 494560 529666
rect 474752 529094 475042 529122
rect 484702 529094 484992 529122
rect 474752 526998 474780 529094
rect 484964 526998 484992 529094
rect 494716 527134 494744 550802
rect 511632 550724 511684 550730
rect 511632 550666 511684 550672
rect 522304 550724 522356 550730
rect 522304 550666 522356 550672
rect 496084 550656 496136 550662
rect 496084 550598 496136 550604
rect 494704 527128 494756 527134
rect 494704 527070 494756 527076
rect 496096 526998 496124 550598
rect 511644 548964 511672 550666
rect 521292 550656 521344 550662
rect 521292 550598 521344 550604
rect 521304 548964 521332 550598
rect 501064 548270 501998 548298
rect 500866 539200 500922 539209
rect 500866 539135 500922 539144
rect 496818 538520 496874 538529
rect 496818 538455 496874 538464
rect 496832 529922 496860 538455
rect 500880 529922 500908 539135
rect 496820 529916 496872 529922
rect 496820 529858 496872 529864
rect 500868 529916 500920 529922
rect 500868 529858 500920 529864
rect 501064 526998 501092 548270
rect 522316 538214 522344 550666
rect 522396 550656 522448 550662
rect 522396 550598 522448 550604
rect 521856 538186 522344 538214
rect 521856 529666 521884 538186
rect 521410 529638 521884 529666
rect 501616 529094 501998 529122
rect 511750 529094 511856 529122
rect 501616 527134 501644 529094
rect 501604 527128 501656 527134
rect 501604 527070 501656 527076
rect 474740 526992 474792 526998
rect 474740 526934 474792 526940
rect 484952 526992 485004 526998
rect 484952 526934 485004 526940
rect 496084 526992 496136 526998
rect 496084 526934 496136 526940
rect 501052 526992 501104 526998
rect 501052 526934 501104 526940
rect 511828 526930 511856 529094
rect 522408 526930 522436 550598
rect 526444 548548 526496 548554
rect 526444 548490 526496 548496
rect 526456 539345 526484 548490
rect 526442 539336 526498 539345
rect 526442 539271 526498 539280
rect 523038 538520 523094 538529
rect 523038 538455 523094 538464
rect 523052 529854 523080 538455
rect 523040 529848 523092 529854
rect 523040 529790 523092 529796
rect 150716 526924 150768 526930
rect 150716 526866 150768 526872
rect 160560 526924 160612 526930
rect 160560 526866 160612 526872
rect 171784 526924 171836 526930
rect 171784 526866 171836 526872
rect 215024 526924 215076 526930
rect 215024 526866 215076 526872
rect 225604 526924 225656 526930
rect 225604 526866 225656 526872
rect 268936 526924 268988 526930
rect 268936 526866 268988 526872
rect 279424 526924 279476 526930
rect 279424 526866 279476 526872
rect 286140 526924 286192 526930
rect 286140 526866 286192 526872
rect 295984 526924 296036 526930
rect 295984 526866 296036 526872
rect 307024 526924 307076 526930
rect 307024 526866 307076 526872
rect 311992 526924 312044 526930
rect 311992 526866 312044 526872
rect 322848 526924 322900 526930
rect 322848 526866 322900 526872
rect 333244 526924 333296 526930
rect 333244 526866 333296 526872
rect 339592 526924 339644 526930
rect 339592 526866 339644 526872
rect 350080 526924 350132 526930
rect 350080 526866 350132 526872
rect 359556 526924 359608 526930
rect 359556 526866 359608 526872
rect 365812 526924 365864 526930
rect 365812 526866 365864 526872
rect 376576 526924 376628 526930
rect 376576 526866 376628 526872
rect 387064 526924 387116 526930
rect 387064 526866 387116 526872
rect 393412 526924 393464 526930
rect 393412 526866 393464 526872
rect 403992 526924 404044 526930
rect 403992 526866 404044 526872
rect 414664 526924 414716 526930
rect 414664 526866 414716 526872
rect 458088 526924 458140 526930
rect 458088 526866 458140 526872
rect 468576 526924 468628 526930
rect 468576 526866 468628 526872
rect 511816 526924 511868 526930
rect 511816 526866 511868 526872
rect 522396 526924 522448 526930
rect 522396 526866 522448 526872
rect 527100 525774 527128 674183
rect 550652 673713 550680 683198
rect 550638 673704 550694 673713
rect 550638 673639 550694 673648
rect 529032 662250 529060 664020
rect 529020 662244 529072 662250
rect 529020 662186 529072 662192
rect 529020 658980 529072 658986
rect 529020 658922 529072 658928
rect 529032 656948 529060 658922
rect 538680 658368 538732 658374
rect 538680 658310 538732 658316
rect 538692 656948 538720 658310
rect 548340 658300 548392 658306
rect 548340 658242 548392 658248
rect 548352 656948 548380 658242
rect 550640 655580 550692 655586
rect 550640 655522 550692 655528
rect 550652 646649 550680 655522
rect 550638 646640 550694 646649
rect 550638 646575 550694 646584
rect 528664 637078 529046 637106
rect 538416 637078 538706 637106
rect 547984 637078 548366 637106
rect 528664 634642 528692 637078
rect 528652 634636 528704 634642
rect 528652 634578 528704 634584
rect 538416 634506 538444 637078
rect 547984 634710 548012 637078
rect 547972 634704 548024 634710
rect 547972 634646 548024 634652
rect 538404 634500 538456 634506
rect 538404 634442 538456 634448
rect 528744 632732 528796 632738
rect 528744 632674 528796 632680
rect 528756 629898 528784 632674
rect 538404 632188 538456 632194
rect 538404 632130 538456 632136
rect 538416 629898 538444 632130
rect 548064 632120 548116 632126
rect 548064 632062 548116 632068
rect 548076 629898 548104 632062
rect 528756 629870 529046 629898
rect 538416 629870 538706 629898
rect 548076 629870 548366 629898
rect 550638 619576 550694 619585
rect 550638 619511 550694 619520
rect 550652 611318 550680 619511
rect 550640 611312 550692 611318
rect 550640 611254 550692 611260
rect 529032 608462 529060 610028
rect 529020 608456 529072 608462
rect 529020 608398 529072 608404
rect 538692 608326 538720 610028
rect 548352 608530 548380 610028
rect 548340 608524 548392 608530
rect 548340 608466 548392 608472
rect 538680 608320 538732 608326
rect 538680 608262 538732 608268
rect 529020 605124 529072 605130
rect 529020 605066 529072 605072
rect 529032 602956 529060 605066
rect 538680 604580 538732 604586
rect 538680 604522 538732 604528
rect 538692 602956 538720 604522
rect 548340 604512 548392 604518
rect 548340 604454 548392 604460
rect 548352 602956 548380 604454
rect 550638 592104 550694 592113
rect 550638 592039 550694 592048
rect 550652 583710 550680 592039
rect 550640 583704 550692 583710
rect 550640 583646 550692 583652
rect 528756 583086 529046 583114
rect 538416 583086 538706 583114
rect 548076 583086 548366 583114
rect 528756 580854 528784 583086
rect 528744 580848 528796 580854
rect 528744 580790 528796 580796
rect 538416 580718 538444 583086
rect 548076 580922 548104 583086
rect 548064 580916 548116 580922
rect 548064 580858 548116 580864
rect 538404 580712 538456 580718
rect 538404 580654 538456 580660
rect 528652 578944 528704 578950
rect 528652 578886 528704 578892
rect 528664 575906 528692 578886
rect 538404 578332 538456 578338
rect 538404 578274 538456 578280
rect 538416 575906 538444 578274
rect 547972 578264 548024 578270
rect 547972 578206 548024 578212
rect 547984 575906 548012 578206
rect 528664 575878 529046 575906
rect 538416 575878 538706 575906
rect 547984 575878 548366 575906
rect 550638 565584 550694 565593
rect 550638 565519 550694 565528
rect 550652 557530 550680 565519
rect 550640 557524 550692 557530
rect 550640 557466 550692 557472
rect 529032 554606 529060 556036
rect 529020 554600 529072 554606
rect 529020 554542 529072 554548
rect 538692 554470 538720 556036
rect 548352 554674 548380 556036
rect 548340 554668 548392 554674
rect 548340 554610 548392 554616
rect 538680 554464 538732 554470
rect 538680 554406 538732 554412
rect 529020 551336 529072 551342
rect 529020 551278 529072 551284
rect 529032 548964 529060 551278
rect 538680 550724 538732 550730
rect 538680 550666 538732 550672
rect 538692 548964 538720 550666
rect 548340 550656 548392 550662
rect 548340 550598 548392 550604
rect 548352 548964 548380 550598
rect 550638 538520 550694 538529
rect 550638 538455 550694 538464
rect 550652 529922 550680 538455
rect 550640 529916 550692 529922
rect 550640 529858 550692 529864
rect 528664 529094 529046 529122
rect 538416 529094 538706 529122
rect 547984 529094 548366 529122
rect 528664 526998 528692 529094
rect 528652 526992 528704 526998
rect 528652 526934 528704 526940
rect 538416 526862 538444 529094
rect 547984 527066 548012 529094
rect 547972 527060 548024 527066
rect 547972 527002 548024 527008
rect 538404 526856 538456 526862
rect 538404 526798 538456 526804
rect 527088 525768 527140 525774
rect 527088 525710 527140 525716
rect 579804 525768 579856 525774
rect 579804 525710 579856 525716
rect 579816 524521 579844 525710
rect 579802 524512 579858 524521
rect 579802 524447 579858 524456
rect 528744 523728 528796 523734
rect 528744 523670 528796 523676
rect 149704 523320 149756 523326
rect 149704 523262 149756 523268
rect 148968 520328 149020 520334
rect 148968 520270 149020 520276
rect 148980 512417 149008 520270
rect 148966 512408 149022 512417
rect 148966 512343 149022 512352
rect 146944 500948 146996 500954
rect 146944 500890 146996 500896
rect 124036 500880 124088 500886
rect 124036 500822 124088 500828
rect 133696 500880 133748 500886
rect 133696 500822 133748 500828
rect 144276 500880 144328 500886
rect 144276 500822 144328 500828
rect 79692 500812 79744 500818
rect 79692 500754 79744 500760
rect 90364 500812 90416 500818
rect 90364 500754 90416 500760
rect 106648 500812 106700 500818
rect 106648 500754 106700 500760
rect 116584 500812 116636 500818
rect 116584 500754 116636 500760
rect 122932 500812 122984 500818
rect 122932 500754 122984 500760
rect 146944 497140 146996 497146
rect 146944 497082 146996 497088
rect 52644 497072 52696 497078
rect 52644 497014 52696 497020
rect 43076 496868 43128 496874
rect 43076 496810 43128 496816
rect 43088 494972 43116 496810
rect 52656 494972 52684 497014
rect 62488 497004 62540 497010
rect 62488 496946 62540 496952
rect 79692 497004 79744 497010
rect 79692 496946 79744 496952
rect 90364 497004 90416 497010
rect 90364 496946 90416 496952
rect 106648 497004 106700 497010
rect 106648 496946 106700 496952
rect 116492 497004 116544 497010
rect 116492 496946 116544 496952
rect 133696 497004 133748 497010
rect 133696 496946 133748 496952
rect 62304 496936 62356 496942
rect 62304 496878 62356 496884
rect 62316 494972 62344 496878
rect 37924 494760 37976 494766
rect 37924 494702 37976 494708
rect 41328 494080 41380 494086
rect 41328 494022 41380 494028
rect 41340 485353 41368 494022
rect 41326 485344 41382 485353
rect 41326 485279 41382 485288
rect 37922 484936 37978 484945
rect 37922 484871 37978 484880
rect 36820 473204 36872 473210
rect 36820 473146 36872 473152
rect 36636 473068 36688 473074
rect 36636 473010 36688 473016
rect 36728 469328 36780 469334
rect 36728 469270 36780 469276
rect 36636 466540 36688 466546
rect 36636 466482 36688 466488
rect 36544 445460 36596 445466
rect 36544 445402 36596 445408
rect 16028 443692 16080 443698
rect 16028 443634 16080 443640
rect 25688 443284 25740 443290
rect 25688 443226 25740 443232
rect 25700 440980 25728 443226
rect 13728 440292 13780 440298
rect 13728 440234 13780 440240
rect 15212 440286 16054 440314
rect 35374 440286 35940 440314
rect 13740 431361 13768 440234
rect 13726 431352 13782 431361
rect 13726 431287 13782 431296
rect 15212 419422 15240 440286
rect 35912 431954 35940 440286
rect 35912 431926 36584 431954
rect 35624 422272 35676 422278
rect 35624 422214 35676 422220
rect 35636 421682 35664 422214
rect 35374 421654 35664 421682
rect 16054 421110 16344 421138
rect 25714 421110 26096 421138
rect 15200 419416 15252 419422
rect 15200 419358 15252 419364
rect 16316 416090 16344 421110
rect 26068 419354 26096 421110
rect 26056 419348 26108 419354
rect 26056 419290 26108 419296
rect 16304 416084 16356 416090
rect 16304 416026 16356 416032
rect 25964 415744 26016 415750
rect 25964 415686 26016 415692
rect 25976 413930 26004 415686
rect 25714 413902 26004 413930
rect 15212 413222 16054 413250
rect 35374 413222 35664 413250
rect 13726 404288 13782 404297
rect 13726 404223 13782 404232
rect 13740 394670 13768 404223
rect 13728 394664 13780 394670
rect 13728 394606 13780 394612
rect 15212 391882 15240 413222
rect 35636 412690 35664 413222
rect 35624 412684 35676 412690
rect 35624 412626 35676 412632
rect 35374 394602 35664 394618
rect 35374 394596 35676 394602
rect 35374 394590 35624 394596
rect 35624 394538 35676 394544
rect 15200 391876 15252 391882
rect 15200 391818 15252 391824
rect 16040 389842 16068 394060
rect 25700 391814 25728 394060
rect 25688 391808 25740 391814
rect 25688 391750 25740 391756
rect 36556 391678 36584 431926
rect 36648 419218 36676 466482
rect 36740 445738 36768 469270
rect 37936 468518 37964 484871
rect 62500 475674 62528 496946
rect 64144 496936 64196 496942
rect 64144 496878 64196 496884
rect 62764 496868 62816 496874
rect 62764 496810 62816 496816
rect 62422 475646 62528 475674
rect 42812 475102 43010 475130
rect 52762 475102 53144 475130
rect 42812 473278 42840 475102
rect 53116 473278 53144 475102
rect 62776 473346 62804 496810
rect 62764 473340 62816 473346
rect 62764 473282 62816 473288
rect 64156 473278 64184 496878
rect 79704 494972 79732 496946
rect 89352 496936 89404 496942
rect 89352 496878 89404 496884
rect 89364 494972 89392 496878
rect 69124 494278 70058 494306
rect 68928 494148 68980 494154
rect 68928 494090 68980 494096
rect 68940 485761 68968 494090
rect 68926 485752 68982 485761
rect 68926 485687 68982 485696
rect 64878 484528 64934 484537
rect 64878 484463 64934 484472
rect 64892 476066 64920 484463
rect 64880 476060 64932 476066
rect 64880 476002 64932 476008
rect 69124 473278 69152 494278
rect 90376 480254 90404 496946
rect 90456 496936 90508 496942
rect 90456 496878 90508 496884
rect 89824 480226 90404 480254
rect 89824 475674 89852 480226
rect 89378 475646 89852 475674
rect 69768 475102 70058 475130
rect 79718 475102 80008 475130
rect 69768 473346 69796 475102
rect 69756 473340 69808 473346
rect 69756 473282 69808 473288
rect 42800 473272 42852 473278
rect 42800 473214 42852 473220
rect 53104 473272 53156 473278
rect 53104 473214 53156 473220
rect 64144 473272 64196 473278
rect 64144 473214 64196 473220
rect 69112 473272 69164 473278
rect 69112 473214 69164 473220
rect 79980 473210 80008 475102
rect 90468 473210 90496 496878
rect 106660 494972 106688 496946
rect 116308 496936 116360 496942
rect 116308 496878 116360 496884
rect 116320 494972 116348 496878
rect 96724 494278 97014 494306
rect 91100 494080 91152 494086
rect 91100 494022 91152 494028
rect 91112 484673 91140 494022
rect 95146 485208 95202 485217
rect 95146 485143 95202 485152
rect 91098 484664 91154 484673
rect 91098 484599 91154 484608
rect 95160 476066 95188 485143
rect 95148 476060 95200 476066
rect 95148 476002 95200 476008
rect 96724 473346 96752 494278
rect 116228 475658 116334 475674
rect 116504 475658 116532 496946
rect 116584 496936 116636 496942
rect 116584 496878 116636 496884
rect 116216 475652 116334 475658
rect 116268 475646 116334 475652
rect 116492 475652 116544 475658
rect 116216 475594 116268 475600
rect 116492 475594 116544 475600
rect 96816 475102 97014 475130
rect 106568 475102 106674 475130
rect 96712 473340 96764 473346
rect 96712 473282 96764 473288
rect 96816 473278 96844 475102
rect 96804 473272 96856 473278
rect 96804 473214 96856 473220
rect 106568 473210 106596 475102
rect 116596 473210 116624 496878
rect 133708 494972 133736 496946
rect 143356 496936 143408 496942
rect 143356 496878 143408 496884
rect 144276 496936 144328 496942
rect 144276 496878 144328 496884
rect 143368 494972 143396 496878
rect 144184 496868 144236 496874
rect 144184 496810 144236 496816
rect 122944 494278 124062 494306
rect 118700 494148 118752 494154
rect 118700 494090 118752 494096
rect 122748 494148 122800 494154
rect 122748 494090 122800 494096
rect 118712 484673 118740 494090
rect 122760 485353 122788 494090
rect 122746 485344 122802 485353
rect 122746 485279 122802 485288
rect 118698 484664 118754 484673
rect 118698 484599 118754 484608
rect 79968 473204 80020 473210
rect 79968 473146 80020 473152
rect 90456 473204 90508 473210
rect 90456 473146 90508 473152
rect 106556 473204 106608 473210
rect 106556 473146 106608 473152
rect 116584 473204 116636 473210
rect 116584 473146 116636 473152
rect 122944 473142 122972 494278
rect 144196 480254 144224 496810
rect 143736 480226 144224 480254
rect 143736 475674 143764 480226
rect 143382 475646 143764 475674
rect 123680 475102 124062 475130
rect 133722 475102 133828 475130
rect 123680 473278 123708 475102
rect 123668 473272 123720 473278
rect 123668 473214 123720 473220
rect 133800 473210 133828 475102
rect 144288 473210 144316 496878
rect 146298 484528 146354 484537
rect 146298 484463 146354 484472
rect 146312 476066 146340 484463
rect 146300 476060 146352 476066
rect 146300 476002 146352 476008
rect 133788 473204 133840 473210
rect 133788 473146 133840 473152
rect 144276 473204 144328 473210
rect 144276 473146 144328 473152
rect 122932 473136 122984 473142
rect 122932 473078 122984 473084
rect 52460 469464 52512 469470
rect 52460 469406 52512 469412
rect 43352 469260 43404 469266
rect 43352 469202 43404 469208
rect 37924 468512 37976 468518
rect 37924 468454 37976 468460
rect 43364 467922 43392 469202
rect 43102 467894 43392 467922
rect 52472 467922 52500 469406
rect 62488 469396 62540 469402
rect 62488 469338 62540 469344
rect 79324 469396 79376 469402
rect 79324 469338 79376 469344
rect 90456 469396 90508 469402
rect 90456 469338 90508 469344
rect 106372 469396 106424 469402
rect 106372 469338 106424 469344
rect 116492 469396 116544 469402
rect 116492 469338 116544 469344
rect 133420 469396 133472 469402
rect 133420 469338 133472 469344
rect 144276 469396 144328 469402
rect 144276 469338 144328 469344
rect 62120 469328 62172 469334
rect 62120 469270 62172 469276
rect 62132 467922 62160 469270
rect 52472 467894 52670 467922
rect 62132 467894 62330 467922
rect 41328 466540 41380 466546
rect 41328 466482 41380 466488
rect 41340 458425 41368 466482
rect 41326 458416 41382 458425
rect 41326 458351 41382 458360
rect 37922 457056 37978 457065
rect 37922 456991 37978 457000
rect 36728 445732 36780 445738
rect 36728 445674 36780 445680
rect 36728 443216 36780 443222
rect 36728 443158 36780 443164
rect 36740 422278 36768 443158
rect 36820 443080 36872 443086
rect 36820 443022 36872 443028
rect 36728 422272 36780 422278
rect 36728 422214 36780 422220
rect 36832 419354 36860 443022
rect 37936 440910 37964 456991
rect 62500 448746 62528 469338
rect 64144 469328 64196 469334
rect 64144 469270 64196 469276
rect 62764 469260 62816 469266
rect 62764 469202 62816 469208
rect 62422 448718 62528 448746
rect 42996 445670 43024 448052
rect 52748 445670 52776 448052
rect 62776 445738 62804 469202
rect 62764 445732 62816 445738
rect 62764 445674 62816 445680
rect 64156 445670 64184 469270
rect 79336 467922 79364 469338
rect 89076 469328 89128 469334
rect 89076 469270 89128 469276
rect 90364 469328 90416 469334
rect 90364 469270 90416 469276
rect 89088 467922 89116 469270
rect 79336 467894 79718 467922
rect 89088 467894 89378 467922
rect 69124 467214 70058 467242
rect 68928 466608 68980 466614
rect 68928 466550 68980 466556
rect 64880 466472 64932 466478
rect 64880 466414 64932 466420
rect 64892 457745 64920 466414
rect 68940 458969 68968 466550
rect 68926 458960 68982 458969
rect 68926 458895 68982 458904
rect 64878 457736 64934 457745
rect 64878 457671 64934 457680
rect 69124 445670 69152 467214
rect 89720 448520 89772 448526
rect 89378 448468 89720 448474
rect 89378 448462 89772 448468
rect 89378 448446 89760 448462
rect 70044 445738 70072 448052
rect 70032 445732 70084 445738
rect 70032 445674 70084 445680
rect 42984 445664 43036 445670
rect 42984 445606 43036 445612
rect 52736 445664 52788 445670
rect 52736 445606 52788 445612
rect 64144 445664 64196 445670
rect 64144 445606 64196 445612
rect 69112 445664 69164 445670
rect 69112 445606 69164 445612
rect 79704 445602 79732 448052
rect 90376 445602 90404 469270
rect 90468 448526 90496 469338
rect 106384 467922 106412 469338
rect 115940 469328 115992 469334
rect 115940 469270 115992 469276
rect 115952 467922 115980 469270
rect 106384 467894 106674 467922
rect 115952 467894 116334 467922
rect 96724 467214 97014 467242
rect 91100 466540 91152 466546
rect 91100 466482 91152 466488
rect 91112 457745 91140 466482
rect 95148 466472 95200 466478
rect 95148 466414 95200 466420
rect 95160 458425 95188 466414
rect 95146 458416 95202 458425
rect 95146 458351 95202 458360
rect 91098 457736 91154 457745
rect 91098 457671 91154 457680
rect 90456 448520 90508 448526
rect 90456 448462 90508 448468
rect 96724 445738 96752 467214
rect 96712 445732 96764 445738
rect 96712 445674 96764 445680
rect 97000 445670 97028 448052
rect 96988 445664 97040 445670
rect 96988 445606 97040 445612
rect 106660 445602 106688 448052
rect 116320 447930 116348 448052
rect 116504 447930 116532 469338
rect 116584 469328 116636 469334
rect 116584 469270 116636 469276
rect 116320 447902 116532 447930
rect 116596 445602 116624 469270
rect 133432 467922 133460 469338
rect 142988 469328 143040 469334
rect 142988 469270 143040 469276
rect 144184 469328 144236 469334
rect 144184 469270 144236 469276
rect 143000 467922 143028 469270
rect 133432 467894 133722 467922
rect 143000 467894 143382 467922
rect 122944 467214 124062 467242
rect 118700 466608 118752 466614
rect 118700 466550 118752 466556
rect 118712 457745 118740 466550
rect 122748 466540 122800 466546
rect 122748 466482 122800 466488
rect 122760 458425 122788 466482
rect 122746 458416 122802 458425
rect 122746 458351 122802 458360
rect 118698 457736 118754 457745
rect 118698 457671 118754 457680
rect 122944 445602 122972 467214
rect 143632 449676 143684 449682
rect 143632 449618 143684 449624
rect 143644 448746 143672 449618
rect 143382 448718 143672 448746
rect 124048 445670 124076 448052
rect 133708 445670 133736 448052
rect 144196 445670 144224 469270
rect 144288 449682 144316 469338
rect 146300 466472 146352 466478
rect 146300 466414 146352 466420
rect 146312 458153 146340 466414
rect 146298 458144 146354 458153
rect 146298 458079 146354 458088
rect 144276 449676 144328 449682
rect 144276 449618 144328 449624
rect 146956 445738 146984 497082
rect 148968 494080 149020 494086
rect 148968 494022 149020 494028
rect 148980 485353 149008 494022
rect 148966 485344 149022 485353
rect 148966 485279 149022 485288
rect 149716 473278 149744 523262
rect 232320 523252 232372 523258
rect 232320 523194 232372 523200
rect 251824 523252 251876 523258
rect 251824 523194 251876 523200
rect 475384 523252 475436 523258
rect 475384 523194 475436 523200
rect 494704 523252 494756 523258
rect 494704 523194 494756 523200
rect 160284 523184 160336 523190
rect 160284 523126 160336 523132
rect 170496 523184 170548 523190
rect 170496 523126 170548 523132
rect 187792 523184 187844 523190
rect 187792 523126 187844 523132
rect 197544 523184 197596 523190
rect 197544 523126 197596 523132
rect 214380 523184 214432 523190
rect 214380 523126 214432 523132
rect 224500 523184 224552 523190
rect 224500 523126 224552 523132
rect 160296 521914 160324 523126
rect 170036 523116 170088 523122
rect 170036 523058 170088 523064
rect 170048 521914 170076 523058
rect 160296 521886 160678 521914
rect 170048 521886 170338 521914
rect 150544 521206 151018 521234
rect 150544 500818 150572 521206
rect 151004 500886 151032 502044
rect 150992 500880 151044 500886
rect 150992 500822 151044 500828
rect 150532 500812 150584 500818
rect 150532 500754 150584 500760
rect 160664 500750 160692 502044
rect 170324 501922 170352 502044
rect 170508 501922 170536 523126
rect 178408 523116 178460 523122
rect 178408 523058 178460 523064
rect 171784 523048 171836 523054
rect 171784 522990 171836 522996
rect 170324 501894 170536 501922
rect 171796 500750 171824 522990
rect 178420 521914 178448 523058
rect 187804 521914 187832 523126
rect 197452 523048 197504 523054
rect 197452 522990 197504 522996
rect 197464 521914 197492 522990
rect 178066 521886 178448 521914
rect 187726 521886 187832 521914
rect 197386 521886 197492 521914
rect 172520 520396 172572 520402
rect 172520 520338 172572 520344
rect 176568 520396 176620 520402
rect 176568 520338 176620 520344
rect 172532 511737 172560 520338
rect 176580 512961 176608 520338
rect 176566 512952 176622 512961
rect 176566 512887 176622 512896
rect 172518 511728 172574 511737
rect 172518 511663 172574 511672
rect 197556 509234 197584 523126
rect 200764 523116 200816 523122
rect 200764 523058 200816 523064
rect 199384 523048 199436 523054
rect 199384 522990 199436 522996
rect 197464 509206 197584 509234
rect 197464 502738 197492 509206
rect 197386 502710 197492 502738
rect 178052 500818 178080 502044
rect 187712 500818 187740 502044
rect 199396 500818 199424 522990
rect 200120 520328 200172 520334
rect 200120 520270 200172 520276
rect 200132 511737 200160 520270
rect 200118 511728 200174 511737
rect 200118 511663 200174 511672
rect 200776 500954 200804 523058
rect 214392 521914 214420 523126
rect 223948 523048 224000 523054
rect 223948 522990 224000 522996
rect 223960 521914 223988 522990
rect 214392 521886 214682 521914
rect 223960 521886 224342 521914
rect 204364 521206 205022 521234
rect 200764 500948 200816 500954
rect 200764 500890 200816 500896
rect 204364 500818 204392 521206
rect 204904 520328 204956 520334
rect 204904 520270 204956 520276
rect 204916 512961 204944 520270
rect 204902 512952 204958 512961
rect 204902 512887 204958 512896
rect 224512 502738 224540 523126
rect 225604 523048 225656 523054
rect 225604 522990 225656 522996
rect 224342 502710 224540 502738
rect 205008 500954 205036 502044
rect 204996 500948 205048 500954
rect 204996 500890 205048 500896
rect 178040 500812 178092 500818
rect 178040 500754 178092 500760
rect 187700 500812 187752 500818
rect 187700 500754 187752 500760
rect 199384 500812 199436 500818
rect 199384 500754 199436 500760
rect 204352 500812 204404 500818
rect 204352 500754 204404 500760
rect 214668 500750 214696 502044
rect 225616 500750 225644 522990
rect 232332 521914 232360 523194
rect 241520 523184 241572 523190
rect 241520 523126 241572 523132
rect 232070 521886 232360 521914
rect 241532 521914 241560 523126
rect 251456 523116 251508 523122
rect 251456 523058 251508 523064
rect 251180 523048 251232 523054
rect 251180 522990 251232 522996
rect 251192 521914 251220 522990
rect 241532 521886 241730 521914
rect 251192 521886 251390 521914
rect 226340 520396 226392 520402
rect 226340 520338 226392 520344
rect 231860 520396 231912 520402
rect 231860 520338 231912 520344
rect 226352 511737 226380 520338
rect 231872 518906 231900 520338
rect 230388 518900 230440 518906
rect 230388 518842 230440 518848
rect 231860 518900 231912 518906
rect 231860 518842 231912 518848
rect 230400 512417 230428 518842
rect 230386 512408 230442 512417
rect 230386 512343 230442 512352
rect 226338 511728 226394 511737
rect 226338 511663 226394 511672
rect 251468 502738 251496 523058
rect 251390 502710 251496 502738
rect 232056 500818 232084 502044
rect 241716 500818 241744 502044
rect 251836 500954 251864 523194
rect 413468 523184 413520 523190
rect 413468 523126 413520 523132
rect 430580 523184 430632 523190
rect 430580 523126 430632 523132
rect 440516 523184 440568 523190
rect 440516 523126 440568 523132
rect 457260 523184 457312 523190
rect 457260 523126 457312 523132
rect 468484 523184 468536 523190
rect 468484 523126 468536 523132
rect 268292 523116 268344 523122
rect 268292 523058 268344 523064
rect 279516 523116 279568 523122
rect 279516 523058 279568 523064
rect 295800 523116 295852 523122
rect 295800 523058 295852 523064
rect 305552 523116 305604 523122
rect 305552 523058 305604 523064
rect 322388 523116 322440 523122
rect 322388 523058 322440 523064
rect 334624 523116 334676 523122
rect 334624 523058 334676 523064
rect 349804 523116 349856 523122
rect 349804 523058 349856 523064
rect 359556 523116 359608 523122
rect 359556 523058 359608 523064
rect 376300 523116 376352 523122
rect 376300 523058 376352 523064
rect 386512 523116 386564 523122
rect 386512 523058 386564 523064
rect 403348 523116 403400 523122
rect 403348 523058 403400 523064
rect 253204 523048 253256 523054
rect 253204 522990 253256 522996
rect 251824 500948 251876 500954
rect 251824 500890 251876 500896
rect 253216 500818 253244 522990
rect 268304 521914 268332 523058
rect 278044 523048 278096 523054
rect 278044 522990 278096 522996
rect 279424 523048 279476 523054
rect 279424 522990 279476 522996
rect 278056 521914 278084 522990
rect 268304 521886 268686 521914
rect 278056 521886 278346 521914
rect 258184 521206 259026 521234
rect 253940 520328 253992 520334
rect 253940 520270 253992 520276
rect 256608 520328 256660 520334
rect 256608 520270 256660 520276
rect 253952 512009 253980 520270
rect 256620 512417 256648 520270
rect 256606 512408 256662 512417
rect 256606 512343 256662 512352
rect 253938 512000 253994 512009
rect 253938 511935 253994 511944
rect 258184 500818 258212 521206
rect 278688 503668 278740 503674
rect 278688 503610 278740 503616
rect 278700 502738 278728 503610
rect 278346 502710 278728 502738
rect 259012 500954 259040 502044
rect 259000 500948 259052 500954
rect 259000 500890 259052 500896
rect 232044 500812 232096 500818
rect 232044 500754 232096 500760
rect 241704 500812 241756 500818
rect 241704 500754 241756 500760
rect 253204 500812 253256 500818
rect 253204 500754 253256 500760
rect 258172 500812 258224 500818
rect 258172 500754 258224 500760
rect 268672 500750 268700 502044
rect 279436 500750 279464 522990
rect 279528 503674 279556 523058
rect 295812 521914 295840 523058
rect 305460 523048 305512 523054
rect 305460 522990 305512 522996
rect 305472 521914 305500 522990
rect 295734 521886 295840 521914
rect 305394 521886 305500 521914
rect 286074 521478 286180 521506
rect 286152 521422 286180 521478
rect 285772 521416 285824 521422
rect 285772 521358 285824 521364
rect 286140 521416 286192 521422
rect 286140 521358 286192 521364
rect 280160 520396 280212 520402
rect 280160 520338 280212 520344
rect 284208 520396 284260 520402
rect 284208 520338 284260 520344
rect 280172 511737 280200 520338
rect 284220 512961 284248 520338
rect 284206 512952 284262 512961
rect 284206 512887 284262 512896
rect 280158 511728 280214 511737
rect 280158 511663 280214 511672
rect 279516 503668 279568 503674
rect 279516 503610 279568 503616
rect 285784 500818 285812 521358
rect 305564 509234 305592 523058
rect 307024 523048 307076 523054
rect 307024 522990 307076 522996
rect 305472 509206 305592 509234
rect 305472 502738 305500 509206
rect 305394 502710 305500 502738
rect 285772 500812 285824 500818
rect 285772 500754 285824 500760
rect 286060 500750 286088 502044
rect 295720 500750 295748 502044
rect 307036 500750 307064 522990
rect 322400 521914 322428 523058
rect 331956 523048 332008 523054
rect 331956 522990 332008 522996
rect 333244 523048 333296 523054
rect 333244 522990 333296 522996
rect 331968 521914 331996 522990
rect 322400 521886 322690 521914
rect 331968 521886 332350 521914
rect 312004 521206 313030 521234
rect 311808 520464 311860 520470
rect 311808 520406 311860 520412
rect 307760 520328 307812 520334
rect 307760 520270 307812 520276
rect 307772 511737 307800 520270
rect 311820 512417 311848 520406
rect 311806 512408 311862 512417
rect 311806 512343 311862 512352
rect 307758 511728 307814 511737
rect 307758 511663 307814 511672
rect 312004 500750 312032 521206
rect 332508 503668 332560 503674
rect 332508 503610 332560 503616
rect 332520 502738 332548 503610
rect 332350 502710 332548 502738
rect 313016 500818 313044 502044
rect 313004 500812 313056 500818
rect 313004 500754 313056 500760
rect 322676 500750 322704 502044
rect 333256 500750 333284 522990
rect 334636 503674 334664 523058
rect 349816 521914 349844 523058
rect 359464 523048 359516 523054
rect 359464 522990 359516 522996
rect 359476 521914 359504 522990
rect 349738 521886 349844 521914
rect 359398 521886 359504 521914
rect 340078 521354 340184 521370
rect 339592 521348 339644 521354
rect 340078 521348 340196 521354
rect 340078 521342 340144 521348
rect 339592 521290 339644 521296
rect 340144 521290 340196 521296
rect 335360 520396 335412 520402
rect 335360 520338 335412 520344
rect 335372 511737 335400 520338
rect 335358 511728 335414 511737
rect 335358 511663 335414 511672
rect 334624 503668 334676 503674
rect 334624 503610 334676 503616
rect 339604 500750 339632 521290
rect 359568 521098 359596 523058
rect 359740 523048 359792 523054
rect 359740 522990 359792 522996
rect 359476 521070 359596 521098
rect 339868 520328 339920 520334
rect 339868 520270 339920 520276
rect 339880 512961 339908 520270
rect 339866 512952 339922 512961
rect 339866 512887 339922 512896
rect 359476 502738 359504 521070
rect 359752 520826 359780 522990
rect 376312 521914 376340 523058
rect 386052 523048 386104 523054
rect 386052 522990 386104 522996
rect 386064 521914 386092 522990
rect 376312 521886 376694 521914
rect 386064 521886 386354 521914
rect 359398 502710 359504 502738
rect 359568 520798 359780 520826
rect 365824 521206 367034 521234
rect 340064 500818 340092 502044
rect 340052 500812 340104 500818
rect 340052 500754 340104 500760
rect 349724 500750 349752 502044
rect 359568 500750 359596 520798
rect 361580 520464 361632 520470
rect 361580 520406 361632 520412
rect 361592 512009 361620 520406
rect 365628 520396 365680 520402
rect 365628 520338 365680 520344
rect 365640 512417 365668 520338
rect 365626 512408 365682 512417
rect 365626 512343 365682 512352
rect 361578 512000 361634 512009
rect 361578 511935 361634 511944
rect 365824 500750 365852 521206
rect 386524 502738 386552 523058
rect 387064 523048 387116 523054
rect 387064 522990 387116 522996
rect 386354 502710 386552 502738
rect 367020 500818 367048 502044
rect 367008 500812 367060 500818
rect 367008 500754 367060 500760
rect 376680 500750 376708 502044
rect 387076 500750 387104 522990
rect 403360 521914 403388 523058
rect 412916 523048 412968 523054
rect 412916 522990 412968 522996
rect 412928 521914 412956 522990
rect 403360 521886 403650 521914
rect 412928 521886 413310 521914
rect 393424 521206 393990 521234
rect 389180 520328 389232 520334
rect 389180 520270 389232 520276
rect 391848 520328 391900 520334
rect 391848 520270 391900 520276
rect 389192 511737 389220 520270
rect 391860 512961 391888 520270
rect 391846 512952 391902 512961
rect 391846 512887 391902 512896
rect 389178 511728 389234 511737
rect 389178 511663 389234 511672
rect 393424 500750 393452 521206
rect 413480 502738 413508 523126
rect 421288 523116 421340 523122
rect 421288 523058 421340 523064
rect 414664 523048 414716 523054
rect 414664 522990 414716 522996
rect 413402 502710 413508 502738
rect 393976 500818 394004 502044
rect 393964 500812 394016 500818
rect 393964 500754 394016 500760
rect 403728 500750 403756 502044
rect 414676 500750 414704 522990
rect 421300 521914 421328 523058
rect 421038 521886 421328 521914
rect 430592 521914 430620 523126
rect 440240 523048 440292 523054
rect 440240 522990 440292 522996
rect 440252 521914 440280 522990
rect 430592 521886 430698 521914
rect 440252 521886 440358 521914
rect 415400 520396 415452 520402
rect 415400 520338 415452 520344
rect 419448 520396 419500 520402
rect 419448 520338 419500 520344
rect 415412 511737 415440 520338
rect 419460 512417 419488 520338
rect 419446 512408 419502 512417
rect 419446 512343 419502 512352
rect 415398 511728 415454 511737
rect 415398 511663 415454 511672
rect 440528 502738 440556 523126
rect 443644 523116 443696 523122
rect 443644 523058 443696 523064
rect 442264 523048 442316 523054
rect 442264 522990 442316 522996
rect 440358 502710 440556 502738
rect 421024 500818 421052 502044
rect 430684 500818 430712 502044
rect 442276 500818 442304 522990
rect 443000 520328 443052 520334
rect 443000 520270 443052 520276
rect 443012 511873 443040 520270
rect 442998 511864 443054 511873
rect 442998 511799 443054 511808
rect 443656 500954 443684 523058
rect 457272 521914 457300 523126
rect 467012 523048 467064 523054
rect 467012 522990 467064 522996
rect 467024 521914 467052 522990
rect 457272 521886 457654 521914
rect 467024 521886 467314 521914
rect 447244 521206 447994 521234
rect 445668 520328 445720 520334
rect 445668 520270 445720 520276
rect 445680 512417 445708 520270
rect 445666 512408 445722 512417
rect 445666 512343 445722 512352
rect 443644 500948 443696 500954
rect 443644 500890 443696 500896
rect 447244 500818 447272 521206
rect 468496 509234 468524 523126
rect 468576 523048 468628 523054
rect 468576 522990 468628 522996
rect 467852 509206 468524 509234
rect 467852 502874 467880 509206
rect 467760 502846 467880 502874
rect 467760 502738 467788 502846
rect 467406 502710 467788 502738
rect 447980 500954 448008 502044
rect 447968 500948 448020 500954
rect 447968 500890 448020 500896
rect 421012 500812 421064 500818
rect 421012 500754 421064 500760
rect 430672 500812 430724 500818
rect 430672 500754 430724 500760
rect 442264 500812 442316 500818
rect 442264 500754 442316 500760
rect 447232 500812 447284 500818
rect 447232 500754 447284 500760
rect 457732 500750 457760 502044
rect 468588 500750 468616 522990
rect 475396 521914 475424 523194
rect 484400 523184 484452 523190
rect 484400 523126 484452 523132
rect 475042 521886 475424 521914
rect 484412 521914 484440 523126
rect 494520 523116 494572 523122
rect 494520 523058 494572 523064
rect 494060 523048 494112 523054
rect 494060 522990 494112 522996
rect 494072 521914 494100 522990
rect 484412 521886 484702 521914
rect 494072 521886 494362 521914
rect 469220 520396 469272 520402
rect 469220 520338 469272 520344
rect 474832 520396 474884 520402
rect 474832 520338 474884 520344
rect 469232 512009 469260 520338
rect 474844 518906 474872 520338
rect 473268 518900 473320 518906
rect 473268 518842 473320 518848
rect 474832 518900 474884 518906
rect 474832 518842 474884 518848
rect 473280 512961 473308 518842
rect 473266 512952 473322 512961
rect 473266 512887 473322 512896
rect 469218 512000 469274 512009
rect 469218 511935 469274 511944
rect 494532 502738 494560 523058
rect 494362 502710 494560 502738
rect 475028 500818 475056 502044
rect 484688 500818 484716 502044
rect 494716 500954 494744 523194
rect 511356 523116 511408 523122
rect 511356 523058 511408 523064
rect 522396 523116 522448 523122
rect 522396 523058 522448 523064
rect 496084 523048 496136 523054
rect 496084 522990 496136 522996
rect 494704 500948 494756 500954
rect 494704 500890 494756 500896
rect 496096 500818 496124 522990
rect 511368 521914 511396 523058
rect 520924 523048 520976 523054
rect 520924 522990 520976 522996
rect 522304 523048 522356 523054
rect 522304 522990 522356 522996
rect 520936 521914 520964 522990
rect 511368 521886 511658 521914
rect 520936 521886 521318 521914
rect 501064 521206 501998 521234
rect 496820 520328 496872 520334
rect 496820 520270 496872 520276
rect 500868 520328 500920 520334
rect 500868 520270 500920 520276
rect 496832 511737 496860 520270
rect 500880 512961 500908 520270
rect 500866 512952 500922 512961
rect 500866 512887 500922 512896
rect 496818 511728 496874 511737
rect 496818 511663 496874 511672
rect 501064 500818 501092 521206
rect 521752 505640 521804 505646
rect 521752 505582 521804 505588
rect 521764 502738 521792 505582
rect 521410 502710 521792 502738
rect 501984 500954 502012 502044
rect 501972 500948 502024 500954
rect 501972 500890 502024 500896
rect 475016 500812 475068 500818
rect 475016 500754 475068 500760
rect 484676 500812 484728 500818
rect 484676 500754 484728 500760
rect 496084 500812 496136 500818
rect 496084 500754 496136 500760
rect 501052 500812 501104 500818
rect 501052 500754 501104 500760
rect 511736 500750 511764 502044
rect 522316 500750 522344 522990
rect 522408 505646 522436 523058
rect 526444 522300 526496 522306
rect 526444 522242 526496 522248
rect 523040 520396 523092 520402
rect 523040 520338 523092 520344
rect 523052 511737 523080 520338
rect 526456 512417 526484 522242
rect 528756 521914 528784 523670
rect 538404 523116 538456 523122
rect 538404 523058 538456 523064
rect 538416 521914 538444 523058
rect 548064 523048 548116 523054
rect 548064 522990 548116 522996
rect 548076 521914 548104 522990
rect 528756 521886 529046 521914
rect 538416 521886 538706 521914
rect 548076 521886 548366 521914
rect 550640 520328 550692 520334
rect 550640 520270 550692 520276
rect 526442 512408 526498 512417
rect 526442 512343 526498 512352
rect 550652 512009 550680 520270
rect 550638 512000 550694 512009
rect 550638 511935 550694 511944
rect 523038 511728 523094 511737
rect 523038 511663 523094 511672
rect 580262 511320 580318 511329
rect 580262 511255 580318 511264
rect 522396 505640 522448 505646
rect 522396 505582 522448 505588
rect 529032 500818 529060 502044
rect 529020 500812 529072 500818
rect 529020 500754 529072 500760
rect 160652 500744 160704 500750
rect 160652 500686 160704 500692
rect 171784 500744 171836 500750
rect 171784 500686 171836 500692
rect 214656 500744 214708 500750
rect 214656 500686 214708 500692
rect 225604 500744 225656 500750
rect 225604 500686 225656 500692
rect 268660 500744 268712 500750
rect 268660 500686 268712 500692
rect 279424 500744 279476 500750
rect 279424 500686 279476 500692
rect 286048 500744 286100 500750
rect 286048 500686 286100 500692
rect 295708 500744 295760 500750
rect 295708 500686 295760 500692
rect 307024 500744 307076 500750
rect 307024 500686 307076 500692
rect 311992 500744 312044 500750
rect 311992 500686 312044 500692
rect 322664 500744 322716 500750
rect 322664 500686 322716 500692
rect 333244 500744 333296 500750
rect 333244 500686 333296 500692
rect 339592 500744 339644 500750
rect 339592 500686 339644 500692
rect 349712 500744 349764 500750
rect 349712 500686 349764 500692
rect 359556 500744 359608 500750
rect 359556 500686 359608 500692
rect 365812 500744 365864 500750
rect 365812 500686 365864 500692
rect 376668 500744 376720 500750
rect 376668 500686 376720 500692
rect 387064 500744 387116 500750
rect 387064 500686 387116 500692
rect 393412 500744 393464 500750
rect 393412 500686 393464 500692
rect 403716 500744 403768 500750
rect 403716 500686 403768 500692
rect 414664 500744 414716 500750
rect 414664 500686 414716 500692
rect 457720 500744 457772 500750
rect 457720 500686 457772 500692
rect 468576 500744 468628 500750
rect 468576 500686 468628 500692
rect 511724 500744 511776 500750
rect 511724 500686 511776 500692
rect 522304 500744 522356 500750
rect 522304 500686 522356 500692
rect 538692 500682 538720 502044
rect 548352 500886 548380 502044
rect 548340 500880 548392 500886
rect 548340 500822 548392 500828
rect 538680 500676 538732 500682
rect 538680 500618 538732 500624
rect 529020 497480 529072 497486
rect 529020 497422 529072 497428
rect 232044 497072 232096 497078
rect 232044 497014 232096 497020
rect 251824 497072 251876 497078
rect 251824 497014 251876 497020
rect 475016 497072 475068 497078
rect 475016 497014 475068 497020
rect 494704 497072 494756 497078
rect 494704 497014 494756 497020
rect 170496 497004 170548 497010
rect 170496 496946 170548 496952
rect 187700 497004 187752 497010
rect 187700 496946 187752 496952
rect 197452 497004 197504 497010
rect 197452 496946 197504 496952
rect 214656 497004 214708 497010
rect 214656 496946 214708 496952
rect 224500 497004 224552 497010
rect 224500 496946 224552 496952
rect 170312 496936 170364 496942
rect 170312 496878 170364 496884
rect 160652 496868 160704 496874
rect 160652 496810 160704 496816
rect 160664 494972 160692 496810
rect 170324 494972 170352 496878
rect 150544 494278 151018 494306
rect 149704 473272 149756 473278
rect 149704 473214 149756 473220
rect 150544 473210 150572 494278
rect 170232 475658 170338 475674
rect 170508 475658 170536 496946
rect 178040 496936 178092 496942
rect 178040 496878 178092 496884
rect 171784 496868 171836 496874
rect 171784 496810 171836 496816
rect 170220 475652 170338 475658
rect 170272 475646 170338 475652
rect 170496 475652 170548 475658
rect 170220 475594 170272 475600
rect 170496 475594 170548 475600
rect 150728 475102 151018 475130
rect 160572 475102 160678 475130
rect 150532 473204 150584 473210
rect 150532 473146 150584 473152
rect 150728 473142 150756 475102
rect 160572 473142 160600 475102
rect 171796 473142 171824 496810
rect 178052 494972 178080 496878
rect 187712 494972 187740 496946
rect 197360 496868 197412 496874
rect 197360 496810 197412 496816
rect 197372 494972 197400 496810
rect 172520 494148 172572 494154
rect 172520 494090 172572 494096
rect 172532 484673 172560 494090
rect 172518 484664 172574 484673
rect 172518 484599 172574 484608
rect 176566 484664 176622 484673
rect 176566 484599 176622 484608
rect 176580 476066 176608 484599
rect 176568 476060 176620 476066
rect 176568 476002 176620 476008
rect 197464 475674 197492 496946
rect 200764 496936 200816 496942
rect 200764 496878 200816 496884
rect 199384 496868 199436 496874
rect 199384 496810 199436 496816
rect 197386 475646 197492 475674
rect 178066 475102 178172 475130
rect 187726 475102 188016 475130
rect 178144 473210 178172 475102
rect 187988 473210 188016 475102
rect 199396 473210 199424 496810
rect 200120 494080 200172 494086
rect 200120 494022 200172 494028
rect 200132 484673 200160 494022
rect 200118 484664 200174 484673
rect 200118 484599 200174 484608
rect 200776 473346 200804 496878
rect 214668 494972 214696 496946
rect 224316 496868 224368 496874
rect 224316 496810 224368 496816
rect 224328 494972 224356 496810
rect 204364 494278 205022 494306
rect 202788 494080 202840 494086
rect 202788 494022 202840 494028
rect 202800 485353 202828 494022
rect 202786 485344 202842 485353
rect 202786 485279 202842 485288
rect 200764 473340 200816 473346
rect 200764 473282 200816 473288
rect 204364 473210 204392 494278
rect 224512 475674 224540 496946
rect 225604 496868 225656 496874
rect 225604 496810 225656 496816
rect 224342 475646 224540 475674
rect 204640 475102 205022 475130
rect 214682 475102 215064 475130
rect 204640 473346 204668 475102
rect 204628 473340 204680 473346
rect 204628 473282 204680 473288
rect 178132 473204 178184 473210
rect 178132 473146 178184 473152
rect 187976 473204 188028 473210
rect 187976 473146 188028 473152
rect 199384 473204 199436 473210
rect 199384 473146 199436 473152
rect 204352 473204 204404 473210
rect 204352 473146 204404 473152
rect 215036 473142 215064 475102
rect 225616 473142 225644 496810
rect 232056 494972 232084 497014
rect 241704 497004 241756 497010
rect 241704 496946 241756 496952
rect 241716 494972 241744 496946
rect 251456 496936 251508 496942
rect 251456 496878 251508 496884
rect 251364 496868 251416 496874
rect 251364 496810 251416 496816
rect 251376 494972 251404 496810
rect 230388 494148 230440 494154
rect 230388 494090 230440 494096
rect 230400 485353 230428 494090
rect 230386 485344 230442 485353
rect 230386 485279 230442 485288
rect 226338 484528 226394 484537
rect 226338 484463 226394 484472
rect 226352 476066 226380 484463
rect 226340 476060 226392 476066
rect 226340 476002 226392 476008
rect 251468 475674 251496 496878
rect 251390 475646 251496 475674
rect 231872 475102 232070 475130
rect 241730 475102 242112 475130
rect 231872 473210 231900 475102
rect 242084 473210 242112 475102
rect 251836 473346 251864 497014
rect 413468 497004 413520 497010
rect 413468 496946 413520 496952
rect 430672 497004 430724 497010
rect 430672 496946 430724 496952
rect 440516 497004 440568 497010
rect 440516 496946 440568 496952
rect 457628 497004 457680 497010
rect 457628 496946 457680 496952
rect 468576 497004 468628 497010
rect 468576 496946 468628 496952
rect 268660 496936 268712 496942
rect 268660 496878 268712 496884
rect 279516 496936 279568 496942
rect 279516 496878 279568 496884
rect 295708 496936 295760 496942
rect 295708 496878 295760 496884
rect 305460 496936 305512 496942
rect 305460 496878 305512 496884
rect 322664 496936 322716 496942
rect 322664 496878 322716 496884
rect 334624 496936 334676 496942
rect 334624 496878 334676 496884
rect 349712 496936 349764 496942
rect 349712 496878 349764 496884
rect 359464 496936 359516 496942
rect 359464 496878 359516 496884
rect 376668 496936 376720 496942
rect 376668 496878 376720 496884
rect 386512 496936 386564 496942
rect 386512 496878 386564 496884
rect 403624 496936 403676 496942
rect 403624 496878 403676 496884
rect 253204 496868 253256 496874
rect 253204 496810 253256 496816
rect 251824 473340 251876 473346
rect 251824 473282 251876 473288
rect 253216 473210 253244 496810
rect 268672 494972 268700 496878
rect 278320 496868 278372 496874
rect 278320 496810 278372 496816
rect 279424 496868 279476 496874
rect 279424 496810 279476 496816
rect 278332 494972 278360 496810
rect 258184 494278 259026 494306
rect 253940 494080 253992 494086
rect 253940 494022 253992 494028
rect 253952 485217 253980 494022
rect 253938 485208 253994 485217
rect 253938 485143 253994 485152
rect 256606 485208 256662 485217
rect 256606 485143 256662 485152
rect 256620 476066 256648 485143
rect 256608 476060 256660 476066
rect 256608 476002 256660 476008
rect 258184 473210 258212 494278
rect 278688 475992 278740 475998
rect 278688 475934 278740 475940
rect 278700 475674 278728 475934
rect 278346 475646 278728 475674
rect 258736 475102 259026 475130
rect 268686 475102 268976 475130
rect 258736 473346 258764 475102
rect 258724 473340 258776 473346
rect 258724 473282 258776 473288
rect 231860 473204 231912 473210
rect 231860 473146 231912 473152
rect 242072 473204 242124 473210
rect 242072 473146 242124 473152
rect 253204 473204 253256 473210
rect 253204 473146 253256 473152
rect 258172 473204 258224 473210
rect 258172 473146 258224 473152
rect 268948 473142 268976 475102
rect 279436 473142 279464 496810
rect 279528 475998 279556 496878
rect 285784 495094 286088 495122
rect 280160 494148 280212 494154
rect 280160 494090 280212 494096
rect 280172 484673 280200 494090
rect 284208 494080 284260 494086
rect 284208 494022 284260 494028
rect 284220 485761 284248 494022
rect 284206 485752 284262 485761
rect 284206 485687 284262 485696
rect 280158 484664 280214 484673
rect 280158 484599 280214 484608
rect 279516 475992 279568 475998
rect 279516 475934 279568 475940
rect 285784 473142 285812 495094
rect 286060 494972 286088 495094
rect 295720 494972 295748 496878
rect 305368 496868 305420 496874
rect 305368 496810 305420 496816
rect 305380 494972 305408 496810
rect 305472 475674 305500 496878
rect 307024 496868 307076 496874
rect 307024 496810 307076 496816
rect 305394 475646 305500 475674
rect 286074 475102 286180 475130
rect 295734 475102 296024 475130
rect 286152 473210 286180 475102
rect 286140 473204 286192 473210
rect 286140 473146 286192 473152
rect 295996 473142 296024 475102
rect 307036 473142 307064 496810
rect 322676 494972 322704 496878
rect 332324 496868 332376 496874
rect 332324 496810 332376 496816
rect 333244 496868 333296 496874
rect 333244 496810 333296 496816
rect 332336 494972 332364 496810
rect 312004 494278 313030 494306
rect 311808 494148 311860 494154
rect 311808 494090 311860 494096
rect 311820 485353 311848 494090
rect 311806 485344 311862 485353
rect 311806 485279 311862 485288
rect 307758 484528 307814 484537
rect 307758 484463 307814 484472
rect 307772 476066 307800 484463
rect 307760 476060 307812 476066
rect 307760 476002 307812 476008
rect 312004 473142 312032 494278
rect 332508 476060 332560 476066
rect 332508 476002 332560 476008
rect 332520 475674 332548 476002
rect 332350 475646 332548 475674
rect 312648 475102 313030 475130
rect 322690 475102 322888 475130
rect 312648 473210 312676 475102
rect 312636 473204 312688 473210
rect 312636 473146 312688 473152
rect 322860 473142 322888 475102
rect 333256 473142 333284 496810
rect 334636 476066 334664 496878
rect 339604 495094 340092 495122
rect 335360 494080 335412 494086
rect 335360 494022 335412 494028
rect 335372 484673 335400 494022
rect 338026 485208 338082 485217
rect 338026 485143 338082 485152
rect 335358 484664 335414 484673
rect 335358 484599 335414 484608
rect 338040 476066 338068 485143
rect 334624 476060 334676 476066
rect 334624 476002 334676 476008
rect 338028 476060 338080 476066
rect 338028 476002 338080 476008
rect 339604 473142 339632 495094
rect 340064 494972 340092 495094
rect 349724 494972 349752 496878
rect 359372 496868 359424 496874
rect 359372 496810 359424 496816
rect 359384 494972 359412 496810
rect 359476 475674 359504 496878
rect 359556 496868 359608 496874
rect 359556 496810 359608 496816
rect 359398 475646 359504 475674
rect 340078 475102 340184 475130
rect 349738 475102 350120 475130
rect 340156 473210 340184 475102
rect 340144 473204 340196 473210
rect 340144 473146 340196 473152
rect 350092 473142 350120 475102
rect 359568 473142 359596 496810
rect 376680 494972 376708 496878
rect 386328 496868 386380 496874
rect 386328 496810 386380 496816
rect 386340 494972 386368 496810
rect 365824 494278 367034 494306
rect 361580 494148 361632 494154
rect 361580 494090 361632 494096
rect 361592 485217 361620 494090
rect 365628 494080 365680 494086
rect 365628 494022 365680 494028
rect 365640 485353 365668 494022
rect 365626 485344 365682 485353
rect 365626 485279 365682 485288
rect 361578 485208 361634 485217
rect 361578 485143 361634 485152
rect 365824 473142 365852 494278
rect 386524 475674 386552 496878
rect 387064 496868 387116 496874
rect 387064 496810 387116 496816
rect 386354 475646 386552 475674
rect 366744 475102 367034 475130
rect 376588 475102 376694 475130
rect 366744 473210 366772 475102
rect 366732 473204 366784 473210
rect 366732 473146 366784 473152
rect 376588 473142 376616 475102
rect 387076 473142 387104 496810
rect 403636 494972 403664 496878
rect 413284 496868 413336 496874
rect 413284 496810 413336 496816
rect 413296 494972 413324 496810
rect 393424 494278 393990 494306
rect 391846 485208 391902 485217
rect 391846 485143 391902 485152
rect 389178 484528 389234 484537
rect 389178 484463 389234 484472
rect 389192 476066 389220 484463
rect 391860 476066 391888 485143
rect 389180 476060 389232 476066
rect 389180 476002 389232 476008
rect 391848 476060 391900 476066
rect 391848 476002 391900 476008
rect 393424 473142 393452 494278
rect 413480 475674 413508 496946
rect 421012 496936 421064 496942
rect 421012 496878 421064 496884
rect 414664 496868 414716 496874
rect 414664 496810 414716 496816
rect 413402 475646 413508 475674
rect 393608 475102 393990 475130
rect 403742 475102 404032 475130
rect 393608 473210 393636 475102
rect 393596 473204 393648 473210
rect 393596 473146 393648 473152
rect 404004 473142 404032 475102
rect 414676 473142 414704 496810
rect 421024 494972 421052 496878
rect 430684 494972 430712 496946
rect 440332 496868 440384 496874
rect 440332 496810 440384 496816
rect 440344 494972 440372 496810
rect 415400 494080 415452 494086
rect 415400 494022 415452 494028
rect 419448 494080 419500 494086
rect 419448 494022 419500 494028
rect 415412 484673 415440 494022
rect 419460 485353 419488 494022
rect 419446 485344 419502 485353
rect 419446 485279 419502 485288
rect 415398 484664 415454 484673
rect 415398 484599 415454 484608
rect 440528 475674 440556 496946
rect 443644 496936 443696 496942
rect 443644 496878 443696 496884
rect 442264 496868 442316 496874
rect 442264 496810 442316 496816
rect 440358 475646 440556 475674
rect 420932 475102 421038 475130
rect 430698 475102 431080 475130
rect 420932 473210 420960 475102
rect 431052 473210 431080 475102
rect 442276 473210 442304 496810
rect 442998 484528 443054 484537
rect 442998 484463 443054 484472
rect 443012 476066 443040 484463
rect 443000 476060 443052 476066
rect 443000 476002 443052 476008
rect 443656 473346 443684 496878
rect 457640 494972 457668 496946
rect 467288 496868 467340 496874
rect 467288 496810 467340 496816
rect 468484 496868 468536 496874
rect 468484 496810 468536 496816
rect 467300 494972 467328 496810
rect 447244 494278 447994 494306
rect 445666 485208 445722 485217
rect 445666 485143 445722 485152
rect 445680 476066 445708 485143
rect 445668 476060 445720 476066
rect 445668 476002 445720 476008
rect 443644 473340 443696 473346
rect 443644 473282 443696 473288
rect 447244 473210 447272 494278
rect 467656 475992 467708 475998
rect 467656 475934 467708 475940
rect 467668 475674 467696 475934
rect 467406 475646 467696 475674
rect 447704 475102 447994 475130
rect 457746 475102 458128 475130
rect 447704 473346 447732 475102
rect 447692 473340 447744 473346
rect 447692 473282 447744 473288
rect 420920 473204 420972 473210
rect 420920 473146 420972 473152
rect 431040 473204 431092 473210
rect 431040 473146 431092 473152
rect 442264 473204 442316 473210
rect 442264 473146 442316 473152
rect 447232 473204 447284 473210
rect 447232 473146 447284 473152
rect 458100 473142 458128 475102
rect 468496 473142 468524 496810
rect 468588 475998 468616 496946
rect 475028 494972 475056 497014
rect 484676 497004 484728 497010
rect 484676 496946 484728 496952
rect 484688 494972 484716 496946
rect 494520 496936 494572 496942
rect 494520 496878 494572 496884
rect 494336 496868 494388 496874
rect 494336 496810 494388 496816
rect 494348 494972 494376 496810
rect 469220 494080 469272 494086
rect 469220 494022 469272 494028
rect 473268 494080 473320 494086
rect 473268 494022 473320 494028
rect 469232 485217 469260 494022
rect 473280 485761 473308 494022
rect 473266 485752 473322 485761
rect 473266 485687 473322 485696
rect 469218 485208 469274 485217
rect 469218 485143 469274 485152
rect 468576 475992 468628 475998
rect 468576 475934 468628 475940
rect 494532 475674 494560 496878
rect 494362 475646 494560 475674
rect 474752 475102 475042 475130
rect 484702 475102 484992 475130
rect 474752 473210 474780 475102
rect 484964 473210 484992 475102
rect 494716 473346 494744 497014
rect 511632 496936 511684 496942
rect 511632 496878 511684 496884
rect 522396 496936 522448 496942
rect 522396 496878 522448 496884
rect 496084 496868 496136 496874
rect 496084 496810 496136 496816
rect 494704 473340 494756 473346
rect 494704 473282 494756 473288
rect 496096 473210 496124 496810
rect 511644 494972 511672 496878
rect 521292 496868 521344 496874
rect 521292 496810 521344 496816
rect 522304 496868 522356 496874
rect 522304 496810 522356 496816
rect 521304 494972 521332 496810
rect 501064 494278 501998 494306
rect 500868 494148 500920 494154
rect 500868 494090 500920 494096
rect 500880 485353 500908 494090
rect 500866 485344 500922 485353
rect 500866 485279 500922 485288
rect 496818 484528 496874 484537
rect 496818 484463 496874 484472
rect 496832 476066 496860 484463
rect 496820 476060 496872 476066
rect 496820 476002 496872 476008
rect 501064 473210 501092 494278
rect 521752 477692 521804 477698
rect 521752 477634 521804 477640
rect 521764 475674 521792 477634
rect 521410 475646 521792 475674
rect 501616 475102 501998 475130
rect 511750 475102 511948 475130
rect 501616 473346 501644 475102
rect 501604 473340 501656 473346
rect 501604 473282 501656 473288
rect 474740 473204 474792 473210
rect 474740 473146 474792 473152
rect 484952 473204 485004 473210
rect 484952 473146 485004 473152
rect 496084 473204 496136 473210
rect 496084 473146 496136 473152
rect 501052 473204 501104 473210
rect 501052 473146 501104 473152
rect 511920 473142 511948 475102
rect 522316 473142 522344 496810
rect 522408 477698 522436 496878
rect 529032 494972 529060 497422
rect 538680 496936 538732 496942
rect 538680 496878 538732 496884
rect 538692 494972 538720 496878
rect 548340 496868 548392 496874
rect 548340 496810 548392 496816
rect 548352 494972 548380 496810
rect 526444 494760 526496 494766
rect 526444 494702 526496 494708
rect 523040 494080 523092 494086
rect 523040 494022 523092 494028
rect 523052 484673 523080 494022
rect 526456 485353 526484 494702
rect 550640 494148 550692 494154
rect 550640 494090 550692 494096
rect 526442 485344 526498 485353
rect 526442 485279 526498 485288
rect 550652 484673 550680 494090
rect 523038 484664 523094 484673
rect 523038 484599 523094 484608
rect 550638 484664 550694 484673
rect 550638 484599 550694 484608
rect 522396 477692 522448 477698
rect 522396 477634 522448 477640
rect 528664 475102 529046 475130
rect 538416 475102 538706 475130
rect 547984 475102 548366 475130
rect 528664 473210 528692 475102
rect 528652 473204 528704 473210
rect 528652 473146 528704 473152
rect 150716 473136 150768 473142
rect 150716 473078 150768 473084
rect 160560 473136 160612 473142
rect 160560 473078 160612 473084
rect 171784 473136 171836 473142
rect 171784 473078 171836 473084
rect 215024 473136 215076 473142
rect 215024 473078 215076 473084
rect 225604 473136 225656 473142
rect 225604 473078 225656 473084
rect 268936 473136 268988 473142
rect 268936 473078 268988 473084
rect 279424 473136 279476 473142
rect 279424 473078 279476 473084
rect 285772 473136 285824 473142
rect 285772 473078 285824 473084
rect 295984 473136 296036 473142
rect 295984 473078 296036 473084
rect 307024 473136 307076 473142
rect 307024 473078 307076 473084
rect 311992 473136 312044 473142
rect 311992 473078 312044 473084
rect 322848 473136 322900 473142
rect 322848 473078 322900 473084
rect 333244 473136 333296 473142
rect 333244 473078 333296 473084
rect 339592 473136 339644 473142
rect 339592 473078 339644 473084
rect 350080 473136 350132 473142
rect 350080 473078 350132 473084
rect 359556 473136 359608 473142
rect 359556 473078 359608 473084
rect 365812 473136 365864 473142
rect 365812 473078 365864 473084
rect 376576 473136 376628 473142
rect 376576 473078 376628 473084
rect 387064 473136 387116 473142
rect 387064 473078 387116 473084
rect 393412 473136 393464 473142
rect 393412 473078 393464 473084
rect 403992 473136 404044 473142
rect 403992 473078 404044 473084
rect 414664 473136 414716 473142
rect 414664 473078 414716 473084
rect 458088 473136 458140 473142
rect 458088 473078 458140 473084
rect 468484 473136 468536 473142
rect 468484 473078 468536 473084
rect 511908 473136 511960 473142
rect 511908 473078 511960 473084
rect 522304 473136 522356 473142
rect 522304 473078 522356 473084
rect 538416 473074 538444 475102
rect 547984 473278 548012 475102
rect 547972 473272 548024 473278
rect 547972 473214 548024 473220
rect 538404 473068 538456 473074
rect 538404 473010 538456 473016
rect 528744 469872 528796 469878
rect 528744 469814 528796 469820
rect 149704 469532 149756 469538
rect 149704 469474 149756 469480
rect 148968 466472 149020 466478
rect 148968 466414 149020 466420
rect 148980 458425 149008 466414
rect 148966 458416 149022 458425
rect 148966 458351 149022 458360
rect 146944 445732 146996 445738
rect 146944 445674 146996 445680
rect 124036 445664 124088 445670
rect 124036 445606 124088 445612
rect 133696 445664 133748 445670
rect 133696 445606 133748 445612
rect 144184 445664 144236 445670
rect 144184 445606 144236 445612
rect 79692 445596 79744 445602
rect 79692 445538 79744 445544
rect 90364 445596 90416 445602
rect 90364 445538 90416 445544
rect 106648 445596 106700 445602
rect 106648 445538 106700 445544
rect 116584 445596 116636 445602
rect 116584 445538 116636 445544
rect 122932 445596 122984 445602
rect 122932 445538 122984 445544
rect 146944 443284 146996 443290
rect 146944 443226 146996 443232
rect 52644 443216 52696 443222
rect 52644 443158 52696 443164
rect 43352 443012 43404 443018
rect 43352 442954 43404 442960
rect 43364 440994 43392 442954
rect 43102 440966 43392 440994
rect 52656 440980 52684 443158
rect 62488 443148 62540 443154
rect 62488 443090 62540 443096
rect 79692 443148 79744 443154
rect 79692 443090 79744 443096
rect 90456 443148 90508 443154
rect 90456 443090 90508 443096
rect 106648 443148 106700 443154
rect 106648 443090 106700 443096
rect 116492 443148 116544 443154
rect 116492 443090 116544 443096
rect 133696 443148 133748 443154
rect 133696 443090 133748 443096
rect 62304 443080 62356 443086
rect 62304 443022 62356 443028
rect 62316 440980 62344 443022
rect 37924 440904 37976 440910
rect 37924 440846 37976 440852
rect 41328 440360 41380 440366
rect 41328 440302 41380 440308
rect 41340 431361 41368 440302
rect 41326 431352 41382 431361
rect 41326 431287 41382 431296
rect 37922 430944 37978 430953
rect 37922 430879 37978 430888
rect 36820 419348 36872 419354
rect 36820 419290 36872 419296
rect 36636 419212 36688 419218
rect 36636 419154 36688 419160
rect 36728 415676 36780 415682
rect 36728 415618 36780 415624
rect 36636 412684 36688 412690
rect 36636 412626 36688 412632
rect 36544 391672 36596 391678
rect 36544 391614 36596 391620
rect 16028 389836 16080 389842
rect 16028 389778 16080 389784
rect 25964 389496 26016 389502
rect 25964 389438 26016 389444
rect 25976 386866 26004 389438
rect 25714 386838 26004 386866
rect 35374 386430 36032 386458
rect 15580 386294 16054 386322
rect 13726 377224 13782 377233
rect 13726 377159 13782 377168
rect 13740 368490 13768 377159
rect 15580 373994 15608 386294
rect 36004 383654 36032 386430
rect 36004 383626 36584 383654
rect 15212 373966 15608 373994
rect 13728 368484 13780 368490
rect 13728 368426 13780 368432
rect 15212 365634 15240 373966
rect 16054 367118 16160 367146
rect 25714 367118 26096 367146
rect 35374 367118 35664 367146
rect 15200 365628 15252 365634
rect 15200 365570 15252 365576
rect 16132 362234 16160 367118
rect 26068 365566 26096 367118
rect 35636 367062 35664 367118
rect 35624 367056 35676 367062
rect 35624 366998 35676 367004
rect 26056 365560 26108 365566
rect 26056 365502 26108 365508
rect 16120 362228 16172 362234
rect 16120 362170 16172 362176
rect 25688 361888 25740 361894
rect 25688 361830 25740 361836
rect 25700 359924 25728 361830
rect 15212 359230 16054 359258
rect 35374 359230 35664 359258
rect 13726 350296 13782 350305
rect 13726 350231 13782 350240
rect 13740 340882 13768 350231
rect 13728 340876 13780 340882
rect 13728 340818 13780 340824
rect 15212 338026 15240 359230
rect 35636 358834 35664 359230
rect 35624 358828 35676 358834
rect 35624 358770 35676 358776
rect 35624 340808 35676 340814
rect 35374 340756 35624 340762
rect 35374 340750 35676 340756
rect 35374 340734 35664 340750
rect 15200 338020 15252 338026
rect 15200 337962 15252 337968
rect 16040 336054 16068 340068
rect 25700 338094 25728 340068
rect 25688 338088 25740 338094
rect 25688 338030 25740 338036
rect 36556 337822 36584 383626
rect 36648 365430 36676 412626
rect 36740 394602 36768 415618
rect 36820 415540 36872 415546
rect 36820 415482 36872 415488
rect 36728 394596 36780 394602
rect 36728 394538 36780 394544
rect 36832 391814 36860 415482
rect 37936 414730 37964 430879
rect 62500 421682 62528 443090
rect 64144 443080 64196 443086
rect 64144 443022 64196 443028
rect 62764 443012 62816 443018
rect 62764 442954 62816 442960
rect 62422 421654 62528 421682
rect 42812 421110 43010 421138
rect 52762 421110 53144 421138
rect 42812 419422 42840 421110
rect 53116 419490 53144 421110
rect 53104 419484 53156 419490
rect 53104 419426 53156 419432
rect 62776 419422 62804 442954
rect 64156 419490 64184 443022
rect 79704 440980 79732 443090
rect 89352 443080 89404 443086
rect 89352 443022 89404 443028
rect 90364 443080 90416 443086
rect 90364 443022 90416 443028
rect 89364 440980 89392 443022
rect 68928 440428 68980 440434
rect 68928 440370 68980 440376
rect 64880 440292 64932 440298
rect 64880 440234 64932 440240
rect 64892 430681 64920 440234
rect 68940 431633 68968 440370
rect 69124 440286 70058 440314
rect 68926 431624 68982 431633
rect 68926 431559 68982 431568
rect 64878 430672 64934 430681
rect 64878 430607 64934 430616
rect 69124 419490 69152 440286
rect 89720 423836 89772 423842
rect 89720 423778 89772 423784
rect 89732 421682 89760 423778
rect 89378 421654 89760 421682
rect 69768 421110 70058 421138
rect 79718 421110 80008 421138
rect 64144 419484 64196 419490
rect 64144 419426 64196 419432
rect 69112 419484 69164 419490
rect 69112 419426 69164 419432
rect 69768 419422 69796 421110
rect 42800 419416 42852 419422
rect 42800 419358 42852 419364
rect 62764 419416 62816 419422
rect 62764 419358 62816 419364
rect 69756 419416 69808 419422
rect 69756 419358 69808 419364
rect 79980 419354 80008 421110
rect 90376 419354 90404 443022
rect 90468 423842 90496 443090
rect 106660 440980 106688 443090
rect 116308 443080 116360 443086
rect 116308 443022 116360 443028
rect 116320 440980 116348 443022
rect 91100 440360 91152 440366
rect 91100 440302 91152 440308
rect 91112 430681 91140 440302
rect 95148 440292 95200 440298
rect 95148 440234 95200 440240
rect 96724 440286 97014 440314
rect 95160 431361 95188 440234
rect 95146 431352 95202 431361
rect 95146 431287 95202 431296
rect 91098 430672 91154 430681
rect 91098 430607 91154 430616
rect 90456 423836 90508 423842
rect 90456 423778 90508 423784
rect 96724 419490 96752 440286
rect 96816 421110 97014 421138
rect 106568 421110 106674 421138
rect 116228 421110 116334 421138
rect 96712 419484 96764 419490
rect 96712 419426 96764 419432
rect 96816 419422 96844 421110
rect 96804 419416 96856 419422
rect 96804 419358 96856 419364
rect 106568 419354 106596 421110
rect 116228 421002 116256 421110
rect 116504 421002 116532 443090
rect 116584 443080 116636 443086
rect 116584 443022 116636 443028
rect 116228 420974 116532 421002
rect 116596 419354 116624 443022
rect 133708 440980 133736 443090
rect 143356 443080 143408 443086
rect 143356 443022 143408 443028
rect 144276 443080 144328 443086
rect 144276 443022 144328 443028
rect 143368 440980 143396 443022
rect 144184 443012 144236 443018
rect 144184 442954 144236 442960
rect 118700 440428 118752 440434
rect 118700 440370 118752 440376
rect 118712 430681 118740 440370
rect 122748 440360 122800 440366
rect 122748 440302 122800 440308
rect 122760 431361 122788 440302
rect 122944 440286 124062 440314
rect 122746 431352 122802 431361
rect 122746 431287 122802 431296
rect 118698 430672 118754 430681
rect 118698 430607 118754 430616
rect 79968 419348 80020 419354
rect 79968 419290 80020 419296
rect 90364 419348 90416 419354
rect 90364 419290 90416 419296
rect 106556 419348 106608 419354
rect 106556 419290 106608 419296
rect 116584 419348 116636 419354
rect 116584 419290 116636 419296
rect 122944 419286 122972 440286
rect 144196 422294 144224 442954
rect 143736 422266 144224 422294
rect 143736 421682 143764 422266
rect 143382 421654 143764 421682
rect 123680 421110 124062 421138
rect 133722 421110 133828 421138
rect 123680 419422 123708 421110
rect 123668 419416 123720 419422
rect 123668 419358 123720 419364
rect 133800 419354 133828 421110
rect 144288 419354 144316 443022
rect 146300 440292 146352 440298
rect 146300 440234 146352 440240
rect 146312 431225 146340 440234
rect 146298 431216 146354 431225
rect 146298 431151 146354 431160
rect 133788 419348 133840 419354
rect 133788 419290 133840 419296
rect 144276 419348 144328 419354
rect 144276 419290 144328 419296
rect 122932 419280 122984 419286
rect 122932 419222 122984 419228
rect 52460 415676 52512 415682
rect 52460 415618 52512 415624
rect 43352 415608 43404 415614
rect 43352 415550 43404 415556
rect 37924 414724 37976 414730
rect 37924 414666 37976 414672
rect 43364 413930 43392 415550
rect 43102 413902 43392 413930
rect 52472 413930 52500 415618
rect 62764 415608 62816 415614
rect 62764 415550 62816 415556
rect 90456 415608 90508 415614
rect 90456 415550 90508 415556
rect 106372 415608 106424 415614
rect 106372 415550 106424 415556
rect 116492 415608 116544 415614
rect 116492 415550 116544 415556
rect 133420 415608 133472 415614
rect 133420 415550 133472 415556
rect 144276 415608 144328 415614
rect 144276 415550 144328 415556
rect 62120 415540 62172 415546
rect 62120 415482 62172 415488
rect 62132 413930 62160 415482
rect 62488 415472 62540 415478
rect 62488 415414 62540 415420
rect 52472 413902 52670 413930
rect 62132 413902 62330 413930
rect 41326 404288 41382 404297
rect 41326 404223 41382 404232
rect 37922 403064 37978 403073
rect 37922 402999 37978 403008
rect 36820 391808 36872 391814
rect 36820 391750 36872 391756
rect 36820 389428 36872 389434
rect 36820 389370 36872 389376
rect 36728 389292 36780 389298
rect 36728 389234 36780 389240
rect 36740 365566 36768 389234
rect 36832 367062 36860 389370
rect 37936 387122 37964 402999
rect 41340 394602 41368 404223
rect 62500 394754 62528 415414
rect 62422 394726 62528 394754
rect 41328 394596 41380 394602
rect 41328 394538 41380 394544
rect 42996 391882 43024 394060
rect 52748 391950 52776 394060
rect 52736 391944 52788 391950
rect 52736 391886 52788 391892
rect 62776 391882 62804 415550
rect 64144 415540 64196 415546
rect 64144 415482 64196 415488
rect 89076 415540 89128 415546
rect 89076 415482 89128 415488
rect 90364 415540 90416 415546
rect 90364 415482 90416 415488
rect 64156 391950 64184 415482
rect 79324 415472 79376 415478
rect 79324 415414 79376 415420
rect 79336 413930 79364 415414
rect 89088 413930 89116 415482
rect 79336 413902 79718 413930
rect 89088 413902 89378 413930
rect 69124 413222 70058 413250
rect 68926 403744 68982 403753
rect 68926 403679 68982 403688
rect 64878 403608 64934 403617
rect 64878 403543 64934 403552
rect 64892 394670 64920 403543
rect 64880 394664 64932 394670
rect 64880 394606 64932 394612
rect 68940 394534 68968 403679
rect 68928 394528 68980 394534
rect 68928 394470 68980 394476
rect 69124 391950 69152 413222
rect 89720 394664 89772 394670
rect 89378 394612 89720 394618
rect 89378 394606 89772 394612
rect 89378 394590 89760 394606
rect 64144 391944 64196 391950
rect 64144 391886 64196 391892
rect 69112 391944 69164 391950
rect 69112 391886 69164 391892
rect 70044 391882 70072 394060
rect 42984 391876 43036 391882
rect 42984 391818 43036 391824
rect 62764 391876 62816 391882
rect 62764 391818 62816 391824
rect 70032 391876 70084 391882
rect 70032 391818 70084 391824
rect 79704 391814 79732 394060
rect 90376 391814 90404 415482
rect 90468 394670 90496 415550
rect 106384 413930 106412 415550
rect 115940 415540 115992 415546
rect 115940 415482 115992 415488
rect 115952 413930 115980 415482
rect 106384 413902 106674 413930
rect 115952 413902 116334 413930
rect 96724 413222 97014 413250
rect 95146 404288 95202 404297
rect 95146 404223 95202 404232
rect 91098 403608 91154 403617
rect 91098 403543 91154 403552
rect 90456 394664 90508 394670
rect 90456 394606 90508 394612
rect 91112 394602 91140 403543
rect 95160 394670 95188 404223
rect 95148 394664 95200 394670
rect 95148 394606 95200 394612
rect 91100 394596 91152 394602
rect 91100 394538 91152 394544
rect 96724 391950 96752 413222
rect 96712 391944 96764 391950
rect 96712 391886 96764 391892
rect 97000 391882 97028 394060
rect 96988 391876 97040 391882
rect 96988 391818 97040 391824
rect 106660 391814 106688 394060
rect 116320 393938 116348 394060
rect 116504 393938 116532 415550
rect 116584 415540 116636 415546
rect 116584 415482 116636 415488
rect 116320 393910 116532 393938
rect 116596 391814 116624 415482
rect 133432 413930 133460 415550
rect 142988 415540 143040 415546
rect 142988 415482 143040 415488
rect 144184 415540 144236 415546
rect 144184 415482 144236 415488
rect 143000 413930 143028 415482
rect 133432 413902 133722 413930
rect 143000 413902 143382 413930
rect 122944 413222 124062 413250
rect 122746 404288 122802 404297
rect 122746 404223 122802 404232
rect 118698 403608 118754 403617
rect 118698 403543 118754 403552
rect 118712 394534 118740 403543
rect 122760 394602 122788 404223
rect 122748 394596 122800 394602
rect 122748 394538 122800 394544
rect 118700 394528 118752 394534
rect 118700 394470 118752 394476
rect 122944 391814 122972 413222
rect 143632 394664 143684 394670
rect 143382 394612 143632 394618
rect 143382 394606 143684 394612
rect 143382 394590 143672 394606
rect 124048 391882 124076 394060
rect 133708 391882 133736 394060
rect 144196 391882 144224 415482
rect 144288 394670 144316 415550
rect 146298 403336 146354 403345
rect 146298 403271 146354 403280
rect 146312 394670 146340 403271
rect 144276 394664 144328 394670
rect 144276 394606 144328 394612
rect 146300 394664 146352 394670
rect 146300 394606 146352 394612
rect 146956 391882 146984 443226
rect 148968 440292 149020 440298
rect 148968 440234 149020 440240
rect 148980 431361 149008 440234
rect 148966 431352 149022 431361
rect 148966 431287 149022 431296
rect 149716 419422 149744 469474
rect 232320 469464 232372 469470
rect 232320 469406 232372 469412
rect 251824 469464 251876 469470
rect 251824 469406 251876 469412
rect 160284 469396 160336 469402
rect 160284 469338 160336 469344
rect 170496 469396 170548 469402
rect 170496 469338 170548 469344
rect 187792 469396 187844 469402
rect 187792 469338 187844 469344
rect 197544 469396 197596 469402
rect 197544 469338 197596 469344
rect 214380 469396 214432 469402
rect 214380 469338 214432 469344
rect 224500 469396 224552 469402
rect 224500 469338 224552 469344
rect 160296 467922 160324 469338
rect 170036 469328 170088 469334
rect 170036 469270 170088 469276
rect 170048 467922 170076 469270
rect 160296 467894 160678 467922
rect 170048 467894 170338 467922
rect 150544 467214 151018 467242
rect 150544 445602 150572 467214
rect 151004 445670 151032 448052
rect 150992 445664 151044 445670
rect 150992 445606 151044 445612
rect 150532 445596 150584 445602
rect 150532 445538 150584 445544
rect 160664 445534 160692 448052
rect 170324 447930 170352 448052
rect 170508 447930 170536 469338
rect 178408 469328 178460 469334
rect 178408 469270 178460 469276
rect 171784 469260 171836 469266
rect 171784 469202 171836 469208
rect 170324 447902 170536 447930
rect 171796 445534 171824 469202
rect 178420 467922 178448 469270
rect 187804 467922 187832 469338
rect 197452 469260 197504 469266
rect 197452 469202 197504 469208
rect 197464 467922 197492 469202
rect 178066 467894 178448 467922
rect 187726 467894 187832 467922
rect 197386 467894 197492 467922
rect 172520 466540 172572 466546
rect 172520 466482 172572 466488
rect 176568 466540 176620 466546
rect 176568 466482 176620 466488
rect 172532 457745 172560 466482
rect 176580 458969 176608 466482
rect 176566 458960 176622 458969
rect 176566 458895 176622 458904
rect 172518 457736 172574 457745
rect 172518 457671 172574 457680
rect 197556 451274 197584 469338
rect 200764 469328 200816 469334
rect 200764 469270 200816 469276
rect 199384 469260 199436 469266
rect 199384 469202 199436 469208
rect 197464 451246 197584 451274
rect 197464 448746 197492 451246
rect 197386 448718 197492 448746
rect 178052 445602 178080 448052
rect 187712 445602 187740 448052
rect 199396 445602 199424 469202
rect 200120 466472 200172 466478
rect 200120 466414 200172 466420
rect 200132 457745 200160 466414
rect 200118 457736 200174 457745
rect 200118 457671 200174 457680
rect 200776 448526 200804 469270
rect 214392 467922 214420 469338
rect 223948 469260 224000 469266
rect 223948 469202 224000 469208
rect 223960 467922 223988 469202
rect 214392 467894 214682 467922
rect 223960 467894 224342 467922
rect 204364 467214 205022 467242
rect 202788 466472 202840 466478
rect 202788 466414 202840 466420
rect 202800 458425 202828 466414
rect 202786 458416 202842 458425
rect 202786 458351 202842 458360
rect 200764 448520 200816 448526
rect 200764 448462 200816 448468
rect 204364 445602 204392 467214
rect 224512 448746 224540 469338
rect 225604 469260 225656 469266
rect 225604 469202 225656 469208
rect 224342 448718 224540 448746
rect 204628 448520 204680 448526
rect 204680 448468 205022 448474
rect 204628 448462 205022 448468
rect 204640 448446 205022 448462
rect 178040 445596 178092 445602
rect 178040 445538 178092 445544
rect 187700 445596 187752 445602
rect 187700 445538 187752 445544
rect 199384 445596 199436 445602
rect 199384 445538 199436 445544
rect 204352 445596 204404 445602
rect 204352 445538 204404 445544
rect 214668 445534 214696 448052
rect 225616 445534 225644 469202
rect 232332 467922 232360 469406
rect 241520 469396 241572 469402
rect 241520 469338 241572 469344
rect 232070 467894 232360 467922
rect 241532 467922 241560 469338
rect 251456 469328 251508 469334
rect 251456 469270 251508 469276
rect 251180 469260 251232 469266
rect 251180 469202 251232 469208
rect 251192 467922 251220 469202
rect 241532 467894 241730 467922
rect 251192 467894 251390 467922
rect 230388 466608 230440 466614
rect 230388 466550 230440 466556
rect 226340 466540 226392 466546
rect 226340 466482 226392 466488
rect 226352 457745 226380 466482
rect 230400 458425 230428 466550
rect 230386 458416 230442 458425
rect 230386 458351 230442 458360
rect 226338 457736 226394 457745
rect 226338 457671 226394 457680
rect 251468 448746 251496 469270
rect 251390 448718 251496 448746
rect 232056 445602 232084 448052
rect 241716 445602 241744 448052
rect 251836 445738 251864 469406
rect 413468 469396 413520 469402
rect 413468 469338 413520 469344
rect 430580 469396 430632 469402
rect 430580 469338 430632 469344
rect 440516 469396 440568 469402
rect 440516 469338 440568 469344
rect 457260 469396 457312 469402
rect 457260 469338 457312 469344
rect 268292 469328 268344 469334
rect 268292 469270 268344 469276
rect 279516 469328 279568 469334
rect 279516 469270 279568 469276
rect 295800 469328 295852 469334
rect 295800 469270 295852 469276
rect 305552 469328 305604 469334
rect 305552 469270 305604 469276
rect 322388 469328 322440 469334
rect 322388 469270 322440 469276
rect 336004 469328 336056 469334
rect 336004 469270 336056 469276
rect 349804 469328 349856 469334
rect 349804 469270 349856 469276
rect 359556 469328 359608 469334
rect 359556 469270 359608 469276
rect 376300 469328 376352 469334
rect 376300 469270 376352 469276
rect 386512 469328 386564 469334
rect 386512 469270 386564 469276
rect 403348 469328 403400 469334
rect 403348 469270 403400 469276
rect 253204 469260 253256 469266
rect 253204 469202 253256 469208
rect 251824 445732 251876 445738
rect 251824 445674 251876 445680
rect 253216 445602 253244 469202
rect 268304 467922 268332 469270
rect 278044 469260 278096 469266
rect 278044 469202 278096 469208
rect 279424 469260 279476 469266
rect 279424 469202 279476 469208
rect 278056 467922 278084 469202
rect 268304 467894 268686 467922
rect 278056 467894 278346 467922
rect 258184 467214 259026 467242
rect 256608 466540 256660 466546
rect 256608 466482 256660 466488
rect 253940 466472 253992 466478
rect 253940 466414 253992 466420
rect 253952 458153 253980 466414
rect 256620 458425 256648 466482
rect 256606 458416 256662 458425
rect 256606 458351 256662 458360
rect 253938 458144 253994 458153
rect 253938 458079 253994 458088
rect 258184 445602 258212 467214
rect 278688 448520 278740 448526
rect 278346 448468 278688 448474
rect 278346 448462 278740 448468
rect 278346 448446 278728 448462
rect 259012 445738 259040 448052
rect 259000 445732 259052 445738
rect 259000 445674 259052 445680
rect 232044 445596 232096 445602
rect 232044 445538 232096 445544
rect 241704 445596 241756 445602
rect 241704 445538 241756 445544
rect 253204 445596 253256 445602
rect 253204 445538 253256 445544
rect 258172 445596 258224 445602
rect 258172 445538 258224 445544
rect 268672 445534 268700 448052
rect 279436 445534 279464 469202
rect 279528 448526 279556 469270
rect 285784 468030 286180 468058
rect 280160 466608 280212 466614
rect 280160 466550 280212 466556
rect 280172 457745 280200 466550
rect 284208 466472 284260 466478
rect 284208 466414 284260 466420
rect 284220 458969 284248 466414
rect 284206 458960 284262 458969
rect 284206 458895 284262 458904
rect 280158 457736 280214 457745
rect 280158 457671 280214 457680
rect 279516 448520 279568 448526
rect 279516 448462 279568 448468
rect 285784 445602 285812 468030
rect 286152 467922 286180 468030
rect 295812 467922 295840 469270
rect 305460 469260 305512 469266
rect 305460 469202 305512 469208
rect 305472 467922 305500 469202
rect 286074 467894 286180 467922
rect 295734 467894 295840 467922
rect 305394 467894 305500 467922
rect 305564 451274 305592 469270
rect 307024 469260 307076 469266
rect 307024 469202 307076 469208
rect 305472 451246 305592 451274
rect 305472 448746 305500 451246
rect 305394 448718 305500 448746
rect 285772 445596 285824 445602
rect 285772 445538 285824 445544
rect 286060 445534 286088 448052
rect 295720 445534 295748 448052
rect 307036 445534 307064 469202
rect 322400 467922 322428 469270
rect 331956 469260 332008 469266
rect 331956 469202 332008 469208
rect 333244 469260 333296 469266
rect 333244 469202 333296 469208
rect 331968 467922 331996 469202
rect 322400 467894 322690 467922
rect 331968 467894 332350 467922
rect 312004 467214 313030 467242
rect 307760 466540 307812 466546
rect 307760 466482 307812 466488
rect 311808 466540 311860 466546
rect 311808 466482 311860 466488
rect 307772 457745 307800 466482
rect 311820 458425 311848 466482
rect 311806 458416 311862 458425
rect 311806 458351 311862 458360
rect 307758 457736 307814 457745
rect 307758 457671 307814 457680
rect 312004 445534 312032 467214
rect 332600 448520 332652 448526
rect 332350 448468 332600 448474
rect 332350 448462 332652 448468
rect 332350 448446 332640 448462
rect 313016 445602 313044 448052
rect 313004 445596 313056 445602
rect 313004 445538 313056 445544
rect 322676 445534 322704 448052
rect 333256 445534 333284 469202
rect 335360 466472 335412 466478
rect 335360 466414 335412 466420
rect 335372 457745 335400 466414
rect 335358 457736 335414 457745
rect 335358 457671 335414 457680
rect 336016 448526 336044 469270
rect 349816 467922 349844 469270
rect 359464 469260 359516 469266
rect 359464 469202 359516 469208
rect 359476 467922 359504 469202
rect 349738 467894 349844 467922
rect 359398 467894 359504 467922
rect 340078 467362 340184 467378
rect 339592 467356 339644 467362
rect 340078 467356 340196 467362
rect 340078 467350 340144 467356
rect 339592 467298 339644 467304
rect 340144 467298 340196 467304
rect 338028 466472 338080 466478
rect 338028 466414 338080 466420
rect 338040 458425 338068 466414
rect 338026 458416 338082 458425
rect 338026 458351 338082 458360
rect 336004 448520 336056 448526
rect 336004 448462 336056 448468
rect 339604 445534 339632 467298
rect 359568 465202 359596 469270
rect 359740 469260 359792 469266
rect 359740 469202 359792 469208
rect 359476 465174 359596 465202
rect 359476 448746 359504 465174
rect 359752 460986 359780 469202
rect 376312 467922 376340 469270
rect 386052 469260 386104 469266
rect 386052 469202 386104 469208
rect 386064 467922 386092 469202
rect 376312 467894 376694 467922
rect 386064 467894 386354 467922
rect 365824 467214 367034 467242
rect 361580 466540 361632 466546
rect 361580 466482 361632 466488
rect 365628 466540 365680 466546
rect 365628 466482 365680 466488
rect 359398 448718 359504 448746
rect 359568 460958 359780 460986
rect 340064 445602 340092 448052
rect 340052 445596 340104 445602
rect 340052 445538 340104 445544
rect 349724 445534 349752 448052
rect 359568 445534 359596 460958
rect 361592 458153 361620 466482
rect 365640 458425 365668 466482
rect 365626 458416 365682 458425
rect 365626 458351 365682 458360
rect 361578 458144 361634 458153
rect 361578 458079 361634 458088
rect 365824 445602 365852 467214
rect 386524 448746 386552 469270
rect 387064 469260 387116 469266
rect 387064 469202 387116 469208
rect 386354 448718 386552 448746
rect 365812 445596 365864 445602
rect 365812 445538 365864 445544
rect 367020 445534 367048 448052
rect 376680 445534 376708 448052
rect 387076 445534 387104 469202
rect 403360 467922 403388 469270
rect 412916 469260 412968 469266
rect 412916 469202 412968 469208
rect 412928 467922 412956 469202
rect 403360 467894 403650 467922
rect 412928 467894 413310 467922
rect 393424 467214 393990 467242
rect 389180 466472 389232 466478
rect 389180 466414 389232 466420
rect 391848 466472 391900 466478
rect 391848 466414 391900 466420
rect 389192 457745 389220 466414
rect 391860 458969 391888 466414
rect 391846 458960 391902 458969
rect 391846 458895 391902 458904
rect 389178 457736 389234 457745
rect 389178 457671 389234 457680
rect 393424 445534 393452 467214
rect 413480 448746 413508 469338
rect 421288 469328 421340 469334
rect 421288 469270 421340 469276
rect 414664 469260 414716 469266
rect 414664 469202 414716 469208
rect 413402 448718 413508 448746
rect 393976 445602 394004 448052
rect 393964 445596 394016 445602
rect 393964 445538 394016 445544
rect 403728 445534 403756 448052
rect 414676 445534 414704 469202
rect 421300 467922 421328 469270
rect 421038 467894 421328 467922
rect 430592 467922 430620 469338
rect 440240 469260 440292 469266
rect 440240 469202 440292 469208
rect 440252 467922 440280 469202
rect 430592 467894 430698 467922
rect 440252 467894 440358 467922
rect 415400 466540 415452 466546
rect 415400 466482 415452 466488
rect 419448 466540 419500 466546
rect 419448 466482 419500 466488
rect 415412 457745 415440 466482
rect 419460 458425 419488 466482
rect 419446 458416 419502 458425
rect 419446 458351 419502 458360
rect 415398 457736 415454 457745
rect 415398 457671 415454 457680
rect 440528 448746 440556 469338
rect 446404 469328 446456 469334
rect 446404 469270 446456 469276
rect 442264 469260 442316 469266
rect 442264 469202 442316 469208
rect 440358 448718 440556 448746
rect 421024 445602 421052 448052
rect 430684 445602 430712 448052
rect 442276 445602 442304 469202
rect 443000 466472 443052 466478
rect 443000 466414 443052 466420
rect 445668 466472 445720 466478
rect 445668 466414 445720 466420
rect 443012 458153 443040 466414
rect 445680 458425 445708 466414
rect 445666 458416 445722 458425
rect 445666 458351 445722 458360
rect 442998 458144 443054 458153
rect 442998 458079 443054 458088
rect 446416 448526 446444 469270
rect 457272 467922 457300 469338
rect 467472 469328 467524 469334
rect 467472 469270 467524 469276
rect 484400 469328 484452 469334
rect 484400 469270 484452 469276
rect 494520 469328 494572 469334
rect 494520 469270 494572 469276
rect 511356 469328 511408 469334
rect 511356 469270 511408 469276
rect 522304 469328 522356 469334
rect 522304 469270 522356 469276
rect 467012 469260 467064 469266
rect 467012 469202 467064 469208
rect 467024 467922 467052 469202
rect 457272 467894 457654 467922
rect 467024 467894 467314 467922
rect 447244 467214 447994 467242
rect 446404 448520 446456 448526
rect 446404 448462 446456 448468
rect 447244 445602 447272 467214
rect 467484 448746 467512 469270
rect 468484 469260 468536 469266
rect 468484 469202 468536 469208
rect 467406 448718 467512 448746
rect 447692 448520 447744 448526
rect 447744 448468 447994 448474
rect 447692 448462 447994 448468
rect 447704 448446 447994 448462
rect 421012 445596 421064 445602
rect 421012 445538 421064 445544
rect 430672 445596 430724 445602
rect 430672 445538 430724 445544
rect 442264 445596 442316 445602
rect 442264 445538 442316 445544
rect 447232 445596 447284 445602
rect 447232 445538 447284 445544
rect 457732 445534 457760 448052
rect 468496 445534 468524 469202
rect 484412 467922 484440 469270
rect 494060 469260 494112 469266
rect 494060 469202 494112 469208
rect 494072 467922 494100 469202
rect 484412 467894 484702 467922
rect 494072 467894 494362 467922
rect 474844 467214 475042 467242
rect 469220 466540 469272 466546
rect 469220 466482 469272 466488
rect 473268 466540 473320 466546
rect 473268 466482 473320 466488
rect 469232 458153 469260 466482
rect 473280 458969 473308 466482
rect 473266 458960 473322 458969
rect 473266 458895 473322 458904
rect 469218 458144 469274 458153
rect 469218 458079 469274 458088
rect 474844 445534 474872 467214
rect 494532 448746 494560 469270
rect 496084 469260 496136 469266
rect 496084 469202 496136 469208
rect 494362 448718 494560 448746
rect 475028 445602 475056 448052
rect 475016 445596 475068 445602
rect 475016 445538 475068 445544
rect 484688 445534 484716 448052
rect 496096 445534 496124 469202
rect 511368 467922 511396 469270
rect 520924 469260 520976 469266
rect 520924 469202 520976 469208
rect 520936 467922 520964 469202
rect 511368 467894 511658 467922
rect 520936 467894 521318 467922
rect 501064 467214 501998 467242
rect 496820 466472 496872 466478
rect 496820 466414 496872 466420
rect 500868 466472 500920 466478
rect 500868 466414 500920 466420
rect 496832 457745 496860 466414
rect 500880 458969 500908 466414
rect 500866 458960 500922 458969
rect 500866 458895 500922 458904
rect 496818 457736 496874 457745
rect 496818 457671 496874 457680
rect 501064 445602 501092 467214
rect 522316 451274 522344 469270
rect 522396 469260 522448 469266
rect 522396 469202 522448 469208
rect 521856 451246 522344 451274
rect 521856 448474 521884 451246
rect 521410 448446 521884 448474
rect 501052 445596 501104 445602
rect 501052 445538 501104 445544
rect 501984 445534 502012 448052
rect 511736 445534 511764 448052
rect 522408 445534 522436 469202
rect 526444 468512 526496 468518
rect 526444 468454 526496 468460
rect 523040 466540 523092 466546
rect 523040 466482 523092 466488
rect 523052 457745 523080 466482
rect 526456 458425 526484 468454
rect 528756 467922 528784 469814
rect 538404 469328 538456 469334
rect 538404 469270 538456 469276
rect 538416 467922 538444 469270
rect 548064 469260 548116 469266
rect 548064 469202 548116 469208
rect 548076 467922 548104 469202
rect 528756 467894 529046 467922
rect 538416 467894 538706 467922
rect 548076 467894 548366 467922
rect 550640 466472 550692 466478
rect 550640 466414 550692 466420
rect 526442 458416 526498 458425
rect 526442 458351 526498 458360
rect 550652 458153 550680 466414
rect 550638 458144 550694 458153
rect 550638 458079 550694 458088
rect 523038 457736 523094 457745
rect 523038 457671 523094 457680
rect 529032 445602 529060 448052
rect 529020 445596 529072 445602
rect 529020 445538 529072 445544
rect 160652 445528 160704 445534
rect 160652 445470 160704 445476
rect 171784 445528 171836 445534
rect 171784 445470 171836 445476
rect 214656 445528 214708 445534
rect 214656 445470 214708 445476
rect 225604 445528 225656 445534
rect 225604 445470 225656 445476
rect 268660 445528 268712 445534
rect 268660 445470 268712 445476
rect 279424 445528 279476 445534
rect 279424 445470 279476 445476
rect 286048 445528 286100 445534
rect 286048 445470 286100 445476
rect 295708 445528 295760 445534
rect 295708 445470 295760 445476
rect 307024 445528 307076 445534
rect 307024 445470 307076 445476
rect 311992 445528 312044 445534
rect 311992 445470 312044 445476
rect 322664 445528 322716 445534
rect 322664 445470 322716 445476
rect 333244 445528 333296 445534
rect 333244 445470 333296 445476
rect 339592 445528 339644 445534
rect 339592 445470 339644 445476
rect 349712 445528 349764 445534
rect 349712 445470 349764 445476
rect 359556 445528 359608 445534
rect 359556 445470 359608 445476
rect 367008 445528 367060 445534
rect 367008 445470 367060 445476
rect 376668 445528 376720 445534
rect 376668 445470 376720 445476
rect 387064 445528 387116 445534
rect 387064 445470 387116 445476
rect 393412 445528 393464 445534
rect 393412 445470 393464 445476
rect 403716 445528 403768 445534
rect 403716 445470 403768 445476
rect 414664 445528 414716 445534
rect 414664 445470 414716 445476
rect 457720 445528 457772 445534
rect 457720 445470 457772 445476
rect 468484 445528 468536 445534
rect 468484 445470 468536 445476
rect 474832 445528 474884 445534
rect 474832 445470 474884 445476
rect 484676 445528 484728 445534
rect 484676 445470 484728 445476
rect 496084 445528 496136 445534
rect 496084 445470 496136 445476
rect 501972 445528 502024 445534
rect 501972 445470 502024 445476
rect 511724 445528 511776 445534
rect 511724 445470 511776 445476
rect 522396 445528 522448 445534
rect 522396 445470 522448 445476
rect 538692 445466 538720 448052
rect 548352 445670 548380 448052
rect 548340 445664 548392 445670
rect 548340 445606 548392 445612
rect 538680 445460 538732 445466
rect 538680 445402 538732 445408
rect 529020 443692 529072 443698
rect 529020 443634 529072 443640
rect 232044 443216 232096 443222
rect 232044 443158 232096 443164
rect 251824 443216 251876 443222
rect 251824 443158 251876 443164
rect 502064 443216 502116 443222
rect 502064 443158 502116 443164
rect 522488 443216 522540 443222
rect 522488 443158 522540 443164
rect 170496 443148 170548 443154
rect 170496 443090 170548 443096
rect 187700 443148 187752 443154
rect 187700 443090 187752 443096
rect 197452 443148 197504 443154
rect 197452 443090 197504 443096
rect 214656 443148 214708 443154
rect 214656 443090 214708 443096
rect 224500 443148 224552 443154
rect 224500 443090 224552 443096
rect 170312 443080 170364 443086
rect 170312 443022 170364 443028
rect 160652 443012 160704 443018
rect 160652 442954 160704 442960
rect 160664 440980 160692 442954
rect 170324 440980 170352 443022
rect 150544 440286 151018 440314
rect 149704 419416 149756 419422
rect 149704 419358 149756 419364
rect 150544 419354 150572 440286
rect 170232 421666 170338 421682
rect 170508 421666 170536 443090
rect 178040 443080 178092 443086
rect 178040 443022 178092 443028
rect 171784 443012 171836 443018
rect 171784 442954 171836 442960
rect 170220 421660 170338 421666
rect 170272 421654 170338 421660
rect 170496 421660 170548 421666
rect 170220 421602 170272 421608
rect 170496 421602 170548 421608
rect 150728 421110 151018 421138
rect 160572 421110 160678 421138
rect 150532 419348 150584 419354
rect 150532 419290 150584 419296
rect 150728 419286 150756 421110
rect 160572 419286 160600 421110
rect 171796 419286 171824 442954
rect 178052 440980 178080 443022
rect 187712 440980 187740 443090
rect 197360 443012 197412 443018
rect 197360 442954 197412 442960
rect 197372 440980 197400 442954
rect 172520 440360 172572 440366
rect 172520 440302 172572 440308
rect 176568 440360 176620 440366
rect 176568 440302 176620 440308
rect 172532 430681 172560 440302
rect 176580 431633 176608 440302
rect 176566 431624 176622 431633
rect 176566 431559 176622 431568
rect 172518 430672 172574 430681
rect 172518 430607 172574 430616
rect 197464 421682 197492 443090
rect 200764 443080 200816 443086
rect 200764 443022 200816 443028
rect 199384 443012 199436 443018
rect 199384 442954 199436 442960
rect 197386 421654 197492 421682
rect 178066 421110 178172 421138
rect 187726 421110 188016 421138
rect 178144 419354 178172 421110
rect 187988 419354 188016 421110
rect 199396 419354 199424 442954
rect 200120 440292 200172 440298
rect 200120 440234 200172 440240
rect 200132 430681 200160 440234
rect 200118 430672 200174 430681
rect 200118 430607 200174 430616
rect 200776 419490 200804 443022
rect 214668 440980 214696 443090
rect 224316 443012 224368 443018
rect 224316 442954 224368 442960
rect 224328 440980 224356 442954
rect 202788 440292 202840 440298
rect 202788 440234 202840 440240
rect 204364 440286 205022 440314
rect 202800 431361 202828 440234
rect 202786 431352 202842 431361
rect 202786 431287 202842 431296
rect 200764 419484 200816 419490
rect 200764 419426 200816 419432
rect 204364 419354 204392 440286
rect 224512 421682 224540 443090
rect 225604 443012 225656 443018
rect 225604 442954 225656 442960
rect 224342 421654 224540 421682
rect 204640 421110 205022 421138
rect 214682 421110 215064 421138
rect 204640 419490 204668 421110
rect 204628 419484 204680 419490
rect 204628 419426 204680 419432
rect 178132 419348 178184 419354
rect 178132 419290 178184 419296
rect 187976 419348 188028 419354
rect 187976 419290 188028 419296
rect 199384 419348 199436 419354
rect 199384 419290 199436 419296
rect 204352 419348 204404 419354
rect 204352 419290 204404 419296
rect 215036 419286 215064 421110
rect 225616 419286 225644 442954
rect 232056 440980 232084 443158
rect 241704 443148 241756 443154
rect 241704 443090 241756 443096
rect 241716 440980 241744 443090
rect 251456 443080 251508 443086
rect 251456 443022 251508 443028
rect 251364 443012 251416 443018
rect 251364 442954 251416 442960
rect 251376 440980 251404 442954
rect 226340 440360 226392 440366
rect 226340 440302 226392 440308
rect 230388 440360 230440 440366
rect 230388 440302 230440 440308
rect 226352 430681 226380 440302
rect 230400 431361 230428 440302
rect 230386 431352 230442 431361
rect 230386 431287 230442 431296
rect 226338 430672 226394 430681
rect 226338 430607 226394 430616
rect 251468 421682 251496 443022
rect 251390 421654 251496 421682
rect 231872 421110 232070 421138
rect 241730 421110 242112 421138
rect 231872 419354 231900 421110
rect 242084 419354 242112 421110
rect 251836 419490 251864 443158
rect 305460 443148 305512 443154
rect 305460 443090 305512 443096
rect 322664 443148 322716 443154
rect 322664 443090 322716 443096
rect 413468 443148 413520 443154
rect 413468 443090 413520 443096
rect 430672 443148 430724 443154
rect 430672 443090 430724 443096
rect 440516 443148 440568 443154
rect 440516 443090 440568 443096
rect 457260 443148 457312 443154
rect 457260 443090 457312 443096
rect 468576 443148 468628 443154
rect 468576 443090 468628 443096
rect 484676 443148 484728 443154
rect 484676 443090 484728 443096
rect 494520 443148 494572 443154
rect 494520 443090 494572 443096
rect 268660 443080 268712 443086
rect 268660 443022 268712 443028
rect 279516 443080 279568 443086
rect 279516 443022 279568 443028
rect 295708 443080 295760 443086
rect 295708 443022 295760 443028
rect 253204 443012 253256 443018
rect 253204 442954 253256 442960
rect 251824 419484 251876 419490
rect 251824 419426 251876 419432
rect 253216 419354 253244 442954
rect 268672 440980 268700 443022
rect 278320 443012 278372 443018
rect 278320 442954 278372 442960
rect 279424 443012 279476 443018
rect 279424 442954 279476 442960
rect 278332 440980 278360 442954
rect 253940 440292 253992 440298
rect 253940 440234 253992 440240
rect 256608 440292 256660 440298
rect 256608 440234 256660 440240
rect 258184 440286 259026 440314
rect 253952 431225 253980 440234
rect 256620 431361 256648 440234
rect 256606 431352 256662 431361
rect 256606 431287 256662 431296
rect 253938 431216 253994 431225
rect 253938 431151 253994 431160
rect 258184 419354 258212 440286
rect 278688 421728 278740 421734
rect 278346 421676 278688 421682
rect 278346 421670 278740 421676
rect 278346 421654 278728 421670
rect 258736 421110 259026 421138
rect 268686 421110 268976 421138
rect 258736 419490 258764 421110
rect 258724 419484 258776 419490
rect 258724 419426 258776 419432
rect 231860 419348 231912 419354
rect 231860 419290 231912 419296
rect 242072 419348 242124 419354
rect 242072 419290 242124 419296
rect 253204 419348 253256 419354
rect 253204 419290 253256 419296
rect 258172 419348 258224 419354
rect 258172 419290 258224 419296
rect 268948 419286 268976 421110
rect 279436 419286 279464 442954
rect 279528 421734 279556 443022
rect 285784 441102 286088 441130
rect 280160 440360 280212 440366
rect 280160 440302 280212 440308
rect 284208 440360 284260 440366
rect 284208 440302 284260 440308
rect 280172 430681 280200 440302
rect 284220 431633 284248 440302
rect 284206 431624 284262 431633
rect 284206 431559 284262 431568
rect 280158 430672 280214 430681
rect 280158 430607 280214 430616
rect 279516 421728 279568 421734
rect 279516 421670 279568 421676
rect 285784 419354 285812 441102
rect 286060 440980 286088 441102
rect 295720 440980 295748 443022
rect 305368 443012 305420 443018
rect 305368 442954 305420 442960
rect 305380 440980 305408 442954
rect 305472 421682 305500 443090
rect 313004 443080 313056 443086
rect 313004 443022 313056 443028
rect 307024 443012 307076 443018
rect 307024 442954 307076 442960
rect 305394 421654 305500 421682
rect 286074 421110 286180 421138
rect 295734 421110 296024 421138
rect 285772 419348 285824 419354
rect 285772 419290 285824 419296
rect 286152 419286 286180 421110
rect 295996 419286 296024 421110
rect 307036 419286 307064 442954
rect 313016 440980 313044 443022
rect 322676 440980 322704 443090
rect 333336 443080 333388 443086
rect 333336 443022 333388 443028
rect 334624 443080 334676 443086
rect 334624 443022 334676 443028
rect 349712 443080 349764 443086
rect 349712 443022 349764 443028
rect 359464 443080 359516 443086
rect 359464 443022 359516 443028
rect 376668 443080 376720 443086
rect 376668 443022 376720 443028
rect 386512 443080 386564 443086
rect 386512 443022 386564 443028
rect 403348 443080 403400 443086
rect 403348 443022 403400 443028
rect 332324 443012 332376 443018
rect 332324 442954 332376 442960
rect 333244 443012 333296 443018
rect 333244 442954 333296 442960
rect 332336 440980 332364 442954
rect 311808 440428 311860 440434
rect 311808 440370 311860 440376
rect 307760 440292 307812 440298
rect 307760 440234 307812 440240
rect 307772 430681 307800 440234
rect 311820 431361 311848 440370
rect 311806 431352 311862 431361
rect 311806 431287 311862 431296
rect 307758 430672 307814 430681
rect 307758 430607 307814 430616
rect 332508 421728 332560 421734
rect 332350 421676 332508 421682
rect 332350 421670 332560 421676
rect 332350 421654 332548 421670
rect 312648 421110 313030 421138
rect 322690 421110 322888 421138
rect 312648 419354 312676 421110
rect 322860 419354 322888 421110
rect 333256 419354 333284 442954
rect 333348 422958 333376 443022
rect 333336 422952 333388 422958
rect 333336 422894 333388 422900
rect 334636 421734 334664 443022
rect 349724 440980 349752 443022
rect 359372 443012 359424 443018
rect 359372 442954 359424 442960
rect 359384 440980 359412 442954
rect 335360 440360 335412 440366
rect 335360 440302 335412 440308
rect 338028 440360 338080 440366
rect 338028 440302 338080 440308
rect 335372 430681 335400 440302
rect 338040 431361 338068 440302
rect 340078 440298 340184 440314
rect 339592 440292 339644 440298
rect 340078 440292 340196 440298
rect 340078 440286 340144 440292
rect 339592 440234 339644 440240
rect 340144 440234 340196 440240
rect 338026 431352 338082 431361
rect 338026 431287 338082 431296
rect 335358 430672 335414 430681
rect 335358 430607 335414 430616
rect 334624 421728 334676 421734
rect 334624 421670 334676 421676
rect 339604 419354 339632 440234
rect 339868 422952 339920 422958
rect 339868 422894 339920 422900
rect 339880 421002 339908 422894
rect 359476 421682 359504 443022
rect 359556 443012 359608 443018
rect 359556 442954 359608 442960
rect 359398 421654 359504 421682
rect 340078 421110 340184 421138
rect 349738 421110 350120 421138
rect 340156 421002 340184 421110
rect 339880 420974 340184 421002
rect 312636 419348 312688 419354
rect 312636 419290 312688 419296
rect 322848 419348 322900 419354
rect 322848 419290 322900 419296
rect 333244 419348 333296 419354
rect 333244 419290 333296 419296
rect 339592 419348 339644 419354
rect 339592 419290 339644 419296
rect 350092 419286 350120 421110
rect 359568 419286 359596 442954
rect 376680 440980 376708 443022
rect 386328 443012 386380 443018
rect 386328 442954 386380 442960
rect 386340 440980 386368 442954
rect 361580 440428 361632 440434
rect 361580 440370 361632 440376
rect 361592 431225 361620 440370
rect 365628 440360 365680 440366
rect 365628 440302 365680 440308
rect 365640 431361 365668 440302
rect 365824 440286 367034 440314
rect 365626 431352 365682 431361
rect 365626 431287 365682 431296
rect 361578 431216 361634 431225
rect 361578 431151 361634 431160
rect 365824 419354 365852 440286
rect 386524 421682 386552 443022
rect 387064 443012 387116 443018
rect 387064 442954 387116 442960
rect 386354 421654 386552 421682
rect 366744 421110 367034 421138
rect 376588 421110 376694 421138
rect 365812 419348 365864 419354
rect 365812 419290 365864 419296
rect 366744 419286 366772 421110
rect 376588 419286 376616 421110
rect 387076 419286 387104 442954
rect 403360 440994 403388 443022
rect 412916 443012 412968 443018
rect 412916 442954 412968 442960
rect 412928 440994 412956 442954
rect 403360 440966 403650 440994
rect 412928 440966 413310 440994
rect 389180 440292 389232 440298
rect 389180 440234 389232 440240
rect 391848 440292 391900 440298
rect 391848 440234 391900 440240
rect 393424 440286 393990 440314
rect 389192 430681 389220 440234
rect 391860 431361 391888 440234
rect 391846 431352 391902 431361
rect 391846 431287 391902 431296
rect 389178 430672 389234 430681
rect 389178 430607 389234 430616
rect 393424 419286 393452 440286
rect 413480 421682 413508 443090
rect 421012 443080 421064 443086
rect 421012 443022 421064 443028
rect 414664 443012 414716 443018
rect 414664 442954 414716 442960
rect 413402 421654 413508 421682
rect 393608 421110 393990 421138
rect 403742 421110 404032 421138
rect 393608 419354 393636 421110
rect 393596 419348 393648 419354
rect 393596 419290 393648 419296
rect 404004 419286 404032 421110
rect 414676 419286 414704 442954
rect 421024 440980 421052 443022
rect 430684 440980 430712 443090
rect 440332 443012 440384 443018
rect 440332 442954 440384 442960
rect 440344 440980 440372 442954
rect 415400 440360 415452 440366
rect 415400 440302 415452 440308
rect 419448 440360 419500 440366
rect 419448 440302 419500 440308
rect 415412 430681 415440 440302
rect 419460 431361 419488 440302
rect 419446 431352 419502 431361
rect 419446 431287 419502 431296
rect 415398 430672 415454 430681
rect 415398 430607 415454 430616
rect 440528 421682 440556 443090
rect 443644 443080 443696 443086
rect 443644 443022 443696 443028
rect 442264 443012 442316 443018
rect 442264 442954 442316 442960
rect 440358 421654 440556 421682
rect 420932 421110 421038 421138
rect 430698 421110 431080 421138
rect 420932 419354 420960 421110
rect 431052 419354 431080 421110
rect 442276 419354 442304 442954
rect 443000 440292 443052 440298
rect 443000 440234 443052 440240
rect 443012 430681 443040 440234
rect 442998 430672 443054 430681
rect 442998 430607 443054 430616
rect 443656 419490 443684 443022
rect 457272 440994 457300 443090
rect 467012 443012 467064 443018
rect 467012 442954 467064 442960
rect 468484 443012 468536 443018
rect 468484 442954 468536 442960
rect 467024 440994 467052 442954
rect 457272 440966 457654 440994
rect 467024 440966 467314 440994
rect 445668 440292 445720 440298
rect 445668 440234 445720 440240
rect 447244 440286 447994 440314
rect 445680 431361 445708 440234
rect 445666 431352 445722 431361
rect 445666 431287 445722 431296
rect 443644 419484 443696 419490
rect 443644 419426 443696 419432
rect 447244 419354 447272 440286
rect 467656 421728 467708 421734
rect 467406 421676 467656 421682
rect 467406 421670 467708 421676
rect 467406 421654 467696 421670
rect 447704 421110 447994 421138
rect 457746 421110 458128 421138
rect 447704 419490 447732 421110
rect 447692 419484 447744 419490
rect 447692 419426 447744 419432
rect 420920 419348 420972 419354
rect 420920 419290 420972 419296
rect 431040 419348 431092 419354
rect 431040 419290 431092 419296
rect 442264 419348 442316 419354
rect 442264 419290 442316 419296
rect 447232 419348 447284 419354
rect 447232 419290 447284 419296
rect 458100 419286 458128 421110
rect 468496 419286 468524 442954
rect 468588 421734 468616 443090
rect 475016 443080 475068 443086
rect 475016 443022 475068 443028
rect 475028 440980 475056 443022
rect 484688 440980 484716 443090
rect 494336 443012 494388 443018
rect 494336 442954 494388 442960
rect 494348 440980 494376 442954
rect 469220 440360 469272 440366
rect 469220 440302 469272 440308
rect 473268 440360 473320 440366
rect 473268 440302 473320 440308
rect 469232 431225 469260 440302
rect 473280 431633 473308 440302
rect 473266 431624 473322 431633
rect 473266 431559 473322 431568
rect 469218 431216 469274 431225
rect 469218 431151 469274 431160
rect 468576 421728 468628 421734
rect 494532 421682 494560 443090
rect 494704 443080 494756 443086
rect 494704 443022 494756 443028
rect 468576 421670 468628 421676
rect 494362 421654 494560 421682
rect 474752 421110 475042 421138
rect 484702 421110 484992 421138
rect 474752 419354 474780 421110
rect 484964 419354 484992 421110
rect 494716 419490 494744 443022
rect 496084 443012 496136 443018
rect 496084 442954 496136 442960
rect 494704 419484 494756 419490
rect 494704 419426 494756 419432
rect 496096 419354 496124 442954
rect 502076 440980 502104 443158
rect 511632 443148 511684 443154
rect 511632 443090 511684 443096
rect 511644 440980 511672 443090
rect 522304 443080 522356 443086
rect 522304 443022 522356 443028
rect 521292 443012 521344 443018
rect 521292 442954 521344 442960
rect 521304 440980 521332 442954
rect 496820 440292 496872 440298
rect 496820 440234 496872 440240
rect 500868 440292 500920 440298
rect 500868 440234 500920 440240
rect 496832 430681 496860 440234
rect 500880 431361 500908 440234
rect 500866 431352 500922 431361
rect 500866 431287 500922 431296
rect 496818 430672 496874 430681
rect 496818 430607 496874 430616
rect 522316 422294 522344 443022
rect 522396 443012 522448 443018
rect 522396 442954 522448 442960
rect 521856 422266 522344 422294
rect 521856 421682 521884 422266
rect 521410 421654 521884 421682
rect 501616 421110 501998 421138
rect 511750 421110 511948 421138
rect 501616 419490 501644 421110
rect 501604 419484 501656 419490
rect 501604 419426 501656 419432
rect 511920 419354 511948 421110
rect 522408 419354 522436 442954
rect 522500 423094 522528 443158
rect 529032 440980 529060 443634
rect 538680 443080 538732 443086
rect 538680 443022 538732 443028
rect 538692 440980 538720 443022
rect 548340 443012 548392 443018
rect 548340 442954 548392 442960
rect 548352 440980 548380 442954
rect 526444 440904 526496 440910
rect 526444 440846 526496 440852
rect 523040 440360 523092 440366
rect 523040 440302 523092 440308
rect 523052 430681 523080 440302
rect 526456 431361 526484 440846
rect 550640 440292 550692 440298
rect 550640 440234 550692 440240
rect 526442 431352 526498 431361
rect 526442 431287 526498 431296
rect 550652 430681 550680 440234
rect 523038 430672 523094 430681
rect 523038 430607 523094 430616
rect 550638 430672 550694 430681
rect 550638 430607 550694 430616
rect 522488 423088 522540 423094
rect 522488 423030 522540 423036
rect 528652 423088 528704 423094
rect 528652 423030 528704 423036
rect 528664 421682 528692 423030
rect 528664 421654 529046 421682
rect 538416 421110 538706 421138
rect 547984 421110 548366 421138
rect 474740 419348 474792 419354
rect 474740 419290 474792 419296
rect 484952 419348 485004 419354
rect 484952 419290 485004 419296
rect 496084 419348 496136 419354
rect 496084 419290 496136 419296
rect 511908 419348 511960 419354
rect 511908 419290 511960 419296
rect 522396 419348 522448 419354
rect 522396 419290 522448 419296
rect 150716 419280 150768 419286
rect 150716 419222 150768 419228
rect 160560 419280 160612 419286
rect 160560 419222 160612 419228
rect 171784 419280 171836 419286
rect 171784 419222 171836 419228
rect 215024 419280 215076 419286
rect 215024 419222 215076 419228
rect 225604 419280 225656 419286
rect 225604 419222 225656 419228
rect 268936 419280 268988 419286
rect 268936 419222 268988 419228
rect 279424 419280 279476 419286
rect 279424 419222 279476 419228
rect 286140 419280 286192 419286
rect 286140 419222 286192 419228
rect 295984 419280 296036 419286
rect 295984 419222 296036 419228
rect 307024 419280 307076 419286
rect 307024 419222 307076 419228
rect 350080 419280 350132 419286
rect 350080 419222 350132 419228
rect 359556 419280 359608 419286
rect 359556 419222 359608 419228
rect 366732 419280 366784 419286
rect 366732 419222 366784 419228
rect 376576 419280 376628 419286
rect 376576 419222 376628 419228
rect 387064 419280 387116 419286
rect 387064 419222 387116 419228
rect 393412 419280 393464 419286
rect 393412 419222 393464 419228
rect 403992 419280 404044 419286
rect 403992 419222 404044 419228
rect 414664 419280 414716 419286
rect 414664 419222 414716 419228
rect 458088 419280 458140 419286
rect 458088 419222 458140 419228
rect 468484 419280 468536 419286
rect 468484 419222 468536 419228
rect 538416 419218 538444 421110
rect 547984 419422 548012 421110
rect 547972 419416 548024 419422
rect 547972 419358 548024 419364
rect 538404 419212 538456 419218
rect 538404 419154 538456 419160
rect 528744 416084 528796 416090
rect 528744 416026 528796 416032
rect 149704 415744 149756 415750
rect 149704 415686 149756 415692
rect 148966 404288 149022 404297
rect 148966 404223 149022 404232
rect 148980 394670 149008 404223
rect 148968 394664 149020 394670
rect 148968 394606 149020 394612
rect 124036 391876 124088 391882
rect 124036 391818 124088 391824
rect 133696 391876 133748 391882
rect 133696 391818 133748 391824
rect 144184 391876 144236 391882
rect 144184 391818 144236 391824
rect 146944 391876 146996 391882
rect 146944 391818 146996 391824
rect 79692 391808 79744 391814
rect 79692 391750 79744 391756
rect 90364 391808 90416 391814
rect 90364 391750 90416 391756
rect 106648 391808 106700 391814
rect 106648 391750 106700 391756
rect 116584 391808 116636 391814
rect 116584 391750 116636 391756
rect 122932 391808 122984 391814
rect 122932 391750 122984 391756
rect 146944 389496 146996 389502
rect 146944 389438 146996 389444
rect 52460 389428 52512 389434
rect 52460 389370 52512 389376
rect 43352 389360 43404 389366
rect 43352 389302 43404 389308
rect 37924 387116 37976 387122
rect 37924 387058 37976 387064
rect 43364 386866 43392 389302
rect 43102 386838 43392 386866
rect 52472 386866 52500 389370
rect 62764 389360 62816 389366
rect 62764 389302 62816 389308
rect 90456 389360 90508 389366
rect 90456 389302 90508 389308
rect 106372 389360 106424 389366
rect 106372 389302 106424 389308
rect 116492 389360 116544 389366
rect 116492 389302 116544 389308
rect 133420 389360 133472 389366
rect 133420 389302 133472 389308
rect 62120 389292 62172 389298
rect 62120 389234 62172 389240
rect 62132 386866 62160 389234
rect 62488 389224 62540 389230
rect 62488 389166 62540 389172
rect 52472 386838 52670 386866
rect 62132 386838 62330 386866
rect 41326 377224 41382 377233
rect 41326 377159 41382 377168
rect 37922 376000 37978 376009
rect 37922 375935 37978 375944
rect 36820 367056 36872 367062
rect 36820 366998 36872 367004
rect 36728 365560 36780 365566
rect 36728 365502 36780 365508
rect 36636 365424 36688 365430
rect 36636 365366 36688 365372
rect 36820 361820 36872 361826
rect 36820 361762 36872 361768
rect 36636 361684 36688 361690
rect 36636 361626 36688 361632
rect 36648 338094 36676 361626
rect 36728 358828 36780 358834
rect 36728 358770 36780 358776
rect 36636 338088 36688 338094
rect 36636 338030 36688 338036
rect 36544 337816 36596 337822
rect 36544 337758 36596 337764
rect 16028 336048 16080 336054
rect 16028 335990 16080 335996
rect 26056 335640 26108 335646
rect 26056 335582 26108 335588
rect 26068 332874 26096 335582
rect 36544 335572 36596 335578
rect 36544 335514 36596 335520
rect 25714 332846 26096 332874
rect 35374 332586 35664 332602
rect 35374 332580 35676 332586
rect 35374 332574 35624 332580
rect 35624 332522 35676 332528
rect 15212 332302 16054 332330
rect 13726 323232 13782 323241
rect 13726 323167 13782 323176
rect 13740 314634 13768 323167
rect 13728 314628 13780 314634
rect 13728 314570 13780 314576
rect 15212 311778 15240 332302
rect 36556 316034 36584 335514
rect 36636 332580 36688 332586
rect 36636 332522 36688 332528
rect 35912 316006 36584 316034
rect 35912 313834 35940 316006
rect 35728 313806 35940 313834
rect 35728 313698 35756 313806
rect 35374 313670 35756 313698
rect 16054 313126 16344 313154
rect 25714 313126 26004 313154
rect 15200 311772 15252 311778
rect 15200 311714 15252 311720
rect 16316 308446 16344 313126
rect 25976 311710 26004 313126
rect 25964 311704 26016 311710
rect 25964 311646 26016 311652
rect 16304 308440 16356 308446
rect 16304 308382 16356 308388
rect 25688 308100 25740 308106
rect 25688 308042 25740 308048
rect 25700 305932 25728 308042
rect 15212 305238 16054 305266
rect 35374 305238 36032 305266
rect 13726 296304 13782 296313
rect 13726 296239 13782 296248
rect 13740 287026 13768 296239
rect 13728 287020 13780 287026
rect 13728 286962 13780 286968
rect 15212 284238 15240 305238
rect 36004 296714 36032 305238
rect 36004 296686 36584 296714
rect 35624 286952 35676 286958
rect 35624 286894 35676 286900
rect 35636 286770 35664 286894
rect 35374 286742 35664 286770
rect 15200 284232 15252 284238
rect 15200 284174 15252 284180
rect 16040 280838 16068 286076
rect 25700 284170 25728 286076
rect 25688 284164 25740 284170
rect 25688 284106 25740 284112
rect 16028 280832 16080 280838
rect 16028 280774 16080 280780
rect 25964 280492 26016 280498
rect 25964 280434 26016 280440
rect 25976 278882 26004 280434
rect 25714 278854 26004 278882
rect 15212 278310 16054 278338
rect 35374 278310 35664 278338
rect 13728 277432 13780 277438
rect 13728 277374 13780 277380
rect 13740 269385 13768 277374
rect 13726 269376 13782 269385
rect 13726 269311 13782 269320
rect 15212 256630 15240 278310
rect 35636 277506 35664 278310
rect 35624 277500 35676 277506
rect 35624 277442 35676 277448
rect 35374 259418 35664 259434
rect 35374 259412 35676 259418
rect 35374 259406 35624 259412
rect 35624 259354 35676 259360
rect 16054 259134 16344 259162
rect 25714 259134 26096 259162
rect 15200 256624 15252 256630
rect 15200 256566 15252 256572
rect 16316 254590 16344 259134
rect 26068 256698 26096 259134
rect 26056 256692 26108 256698
rect 26056 256634 26108 256640
rect 36556 256426 36584 296686
rect 36648 284034 36676 332522
rect 36740 311574 36768 358770
rect 36832 340814 36860 361762
rect 37936 359514 37964 375935
rect 41340 368422 41368 377159
rect 41328 368416 41380 368422
rect 41328 368358 41380 368364
rect 62500 367690 62528 389166
rect 62422 367662 62528 367690
rect 42812 367118 43010 367146
rect 52762 367118 53144 367146
rect 42812 365634 42840 367118
rect 53116 365702 53144 367118
rect 53104 365696 53156 365702
rect 53104 365638 53156 365644
rect 62776 365634 62804 389302
rect 64144 389292 64196 389298
rect 64144 389234 64196 389240
rect 89076 389292 89128 389298
rect 89076 389234 89128 389240
rect 90364 389292 90416 389298
rect 90364 389234 90416 389240
rect 64156 365702 64184 389234
rect 79324 389224 79376 389230
rect 79324 389166 79376 389172
rect 79336 386866 79364 389166
rect 89088 386866 89116 389234
rect 79336 386838 79718 386866
rect 89088 386838 89378 386866
rect 69676 386294 70058 386322
rect 68926 376816 68982 376825
rect 68926 376751 68982 376760
rect 64878 376544 64934 376553
rect 64878 376479 64934 376488
rect 64892 368490 64920 376479
rect 64880 368484 64932 368490
rect 64880 368426 64932 368432
rect 68940 368354 68968 376751
rect 69676 373994 69704 386294
rect 69124 373966 69704 373994
rect 68928 368348 68980 368354
rect 68928 368290 68980 368296
rect 69124 365702 69152 373966
rect 89720 370592 89772 370598
rect 89720 370534 89772 370540
rect 89732 367690 89760 370534
rect 89378 367662 89760 367690
rect 69768 367118 70058 367146
rect 79718 367118 80008 367146
rect 64144 365696 64196 365702
rect 64144 365638 64196 365644
rect 69112 365696 69164 365702
rect 69112 365638 69164 365644
rect 69768 365634 69796 367118
rect 42800 365628 42852 365634
rect 42800 365570 42852 365576
rect 62764 365628 62816 365634
rect 62764 365570 62816 365576
rect 69756 365628 69808 365634
rect 69756 365570 69808 365576
rect 79980 365566 80008 367118
rect 90376 365566 90404 389234
rect 90468 370598 90496 389302
rect 106384 386866 106412 389302
rect 115940 389292 115992 389298
rect 115940 389234 115992 389240
rect 115952 386866 115980 389234
rect 106384 386838 106674 386866
rect 115952 386838 116334 386866
rect 96724 386294 97014 386322
rect 95146 377224 95202 377233
rect 95146 377159 95202 377168
rect 91098 376544 91154 376553
rect 91098 376479 91154 376488
rect 90456 370592 90508 370598
rect 90456 370534 90508 370540
rect 91112 368422 91140 376479
rect 95160 368490 95188 377159
rect 95148 368484 95200 368490
rect 95148 368426 95200 368432
rect 91100 368416 91152 368422
rect 91100 368358 91152 368364
rect 96724 365702 96752 386294
rect 96816 367118 97014 367146
rect 106568 367118 106674 367146
rect 116228 367118 116334 367146
rect 96712 365696 96764 365702
rect 96712 365638 96764 365644
rect 96816 365634 96844 367118
rect 96804 365628 96856 365634
rect 96804 365570 96856 365576
rect 106568 365566 106596 367118
rect 116228 367010 116256 367118
rect 116504 367010 116532 389302
rect 116584 389292 116636 389298
rect 116584 389234 116636 389240
rect 116228 366982 116532 367010
rect 116596 365566 116624 389234
rect 133432 386866 133460 389302
rect 142988 389292 143040 389298
rect 142988 389234 143040 389240
rect 144276 389292 144328 389298
rect 144276 389234 144328 389240
rect 143000 386866 143028 389234
rect 144184 389224 144236 389230
rect 144184 389166 144236 389172
rect 133432 386838 133722 386866
rect 143000 386838 143382 386866
rect 123588 386294 124062 386322
rect 122746 377224 122802 377233
rect 122746 377159 122802 377168
rect 118698 376544 118754 376553
rect 118698 376479 118754 376488
rect 118712 368354 118740 376479
rect 122760 368422 122788 377159
rect 123588 373994 123616 386294
rect 144196 373994 144224 389166
rect 122944 373966 123616 373994
rect 143736 373966 144224 373994
rect 122748 368416 122800 368422
rect 122748 368358 122800 368364
rect 118700 368348 118752 368354
rect 118700 368290 118752 368296
rect 79968 365560 80020 365566
rect 79968 365502 80020 365508
rect 90364 365560 90416 365566
rect 90364 365502 90416 365508
rect 106556 365560 106608 365566
rect 106556 365502 106608 365508
rect 116584 365560 116636 365566
rect 116584 365502 116636 365508
rect 122944 365498 122972 373966
rect 143736 367690 143764 373966
rect 143382 367662 143764 367690
rect 123680 367118 124062 367146
rect 133722 367118 133828 367146
rect 123680 365634 123708 367118
rect 123668 365628 123720 365634
rect 123668 365570 123720 365576
rect 133800 365566 133828 367118
rect 144288 365566 144316 389234
rect 144826 376000 144882 376009
rect 144826 375935 144882 375944
rect 144840 368490 144868 375935
rect 144828 368484 144880 368490
rect 144828 368426 144880 368432
rect 133788 365560 133840 365566
rect 133788 365502 133840 365508
rect 144276 365560 144328 365566
rect 144276 365502 144328 365508
rect 122932 365492 122984 365498
rect 122932 365434 122984 365440
rect 52644 361820 52696 361826
rect 52644 361762 52696 361768
rect 43076 361616 43128 361622
rect 43076 361558 43128 361564
rect 43088 359924 43116 361558
rect 52656 359924 52684 361762
rect 62488 361752 62540 361758
rect 62488 361694 62540 361700
rect 79692 361752 79744 361758
rect 79692 361694 79744 361700
rect 90364 361752 90416 361758
rect 90364 361694 90416 361700
rect 106648 361752 106700 361758
rect 106648 361694 106700 361700
rect 116492 361752 116544 361758
rect 116492 361694 116544 361700
rect 133696 361752 133748 361758
rect 133696 361694 133748 361700
rect 144276 361752 144328 361758
rect 144276 361694 144328 361700
rect 62304 361684 62356 361690
rect 62304 361626 62356 361632
rect 62316 359924 62344 361626
rect 37924 359508 37976 359514
rect 37924 359450 37976 359456
rect 41326 350296 41382 350305
rect 41326 350231 41382 350240
rect 37922 349208 37978 349217
rect 37922 349143 37978 349152
rect 36820 340808 36872 340814
rect 36820 340750 36872 340756
rect 36820 335436 36872 335442
rect 36820 335378 36872 335384
rect 36832 311710 36860 335378
rect 37936 333266 37964 349143
rect 41340 340814 41368 350231
rect 41328 340808 41380 340814
rect 62500 340762 62528 361694
rect 64144 361684 64196 361690
rect 64144 361626 64196 361632
rect 62764 361616 62816 361622
rect 62764 361558 62816 361564
rect 41328 340750 41380 340756
rect 62422 340734 62528 340762
rect 42996 338026 43024 340068
rect 52748 338094 52776 340068
rect 52736 338088 52788 338094
rect 52736 338030 52788 338036
rect 62776 338026 62804 361558
rect 64156 338094 64184 361626
rect 79704 359924 79732 361694
rect 89352 361684 89404 361690
rect 89352 361626 89404 361632
rect 89364 359924 89392 361626
rect 69124 359230 70058 359258
rect 68926 349752 68982 349761
rect 68926 349687 68982 349696
rect 64878 349616 64934 349625
rect 64878 349551 64934 349560
rect 64892 340882 64920 349551
rect 64880 340876 64932 340882
rect 64880 340818 64932 340824
rect 68940 340746 68968 349687
rect 68928 340740 68980 340746
rect 68928 340682 68980 340688
rect 69124 338094 69152 359230
rect 90376 345014 90404 361694
rect 90456 361684 90508 361690
rect 90456 361626 90508 361632
rect 89824 344986 90404 345014
rect 89824 340762 89852 344986
rect 89378 340734 89852 340762
rect 64144 338088 64196 338094
rect 64144 338030 64196 338036
rect 69112 338088 69164 338094
rect 69112 338030 69164 338036
rect 70044 338026 70072 340068
rect 42984 338020 43036 338026
rect 42984 337962 43036 337968
rect 62764 338020 62816 338026
rect 62764 337962 62816 337968
rect 70032 338020 70084 338026
rect 70032 337962 70084 337968
rect 79704 337958 79732 340068
rect 90468 337958 90496 361626
rect 106660 359924 106688 361694
rect 116308 361684 116360 361690
rect 116308 361626 116360 361632
rect 116320 359924 116348 361626
rect 96724 359230 97014 359258
rect 95146 350296 95202 350305
rect 95146 350231 95202 350240
rect 91098 349616 91154 349625
rect 91098 349551 91154 349560
rect 91112 340814 91140 349551
rect 95160 340882 95188 350231
rect 95148 340876 95200 340882
rect 95148 340818 95200 340824
rect 91100 340808 91152 340814
rect 91100 340750 91152 340756
rect 96724 338094 96752 359230
rect 96712 338088 96764 338094
rect 96712 338030 96764 338036
rect 97000 338026 97028 340068
rect 96988 338020 97040 338026
rect 96988 337962 97040 337968
rect 106660 337958 106688 340068
rect 116320 339946 116348 340068
rect 116504 339946 116532 361694
rect 116584 361684 116636 361690
rect 116584 361626 116636 361632
rect 116320 339918 116532 339946
rect 116596 337958 116624 361626
rect 133708 359924 133736 361694
rect 143356 361684 143408 361690
rect 143356 361626 143408 361632
rect 144184 361684 144236 361690
rect 144184 361626 144236 361632
rect 143368 359924 143396 361626
rect 122944 359230 124062 359258
rect 122746 350296 122802 350305
rect 122746 350231 122802 350240
rect 118698 349616 118754 349625
rect 118698 349551 118754 349560
rect 118712 340746 118740 349551
rect 122760 340814 122788 350231
rect 122748 340808 122800 340814
rect 122748 340750 122800 340756
rect 118700 340740 118752 340746
rect 118700 340682 118752 340688
rect 122944 337958 122972 359230
rect 143632 342576 143684 342582
rect 143632 342518 143684 342524
rect 143644 340762 143672 342518
rect 143382 340734 143672 340762
rect 124048 338026 124076 340068
rect 133708 338026 133736 340068
rect 144196 338026 144224 361626
rect 144288 342582 144316 361694
rect 146298 349208 146354 349217
rect 146298 349143 146354 349152
rect 144276 342576 144328 342582
rect 144276 342518 144328 342524
rect 146312 340882 146340 349143
rect 146300 340876 146352 340882
rect 146300 340818 146352 340824
rect 146956 338094 146984 389438
rect 148966 377224 149022 377233
rect 148966 377159 149022 377168
rect 148980 368490 149008 377159
rect 148968 368484 149020 368490
rect 148968 368426 149020 368432
rect 149716 365634 149744 415686
rect 475384 415676 475436 415682
rect 475384 415618 475436 415624
rect 494704 415676 494756 415682
rect 494704 415618 494756 415624
rect 160284 415608 160336 415614
rect 160284 415550 160336 415556
rect 170496 415608 170548 415614
rect 170496 415550 170548 415556
rect 187792 415608 187844 415614
rect 187792 415550 187844 415556
rect 197544 415608 197596 415614
rect 197544 415550 197596 415556
rect 214380 415608 214432 415614
rect 214380 415550 214432 415556
rect 224500 415608 224552 415614
rect 224500 415550 224552 415556
rect 241520 415608 241572 415614
rect 241520 415550 241572 415556
rect 251456 415608 251508 415614
rect 251456 415550 251508 415556
rect 268292 415608 268344 415614
rect 268292 415550 268344 415556
rect 413468 415608 413520 415614
rect 413468 415550 413520 415556
rect 430580 415608 430632 415614
rect 430580 415550 430632 415556
rect 440516 415608 440568 415614
rect 440516 415550 440568 415556
rect 457260 415608 457312 415614
rect 457260 415550 457312 415556
rect 468576 415608 468628 415614
rect 468576 415550 468628 415556
rect 160296 413930 160324 415550
rect 170036 415540 170088 415546
rect 170036 415482 170088 415488
rect 170048 413930 170076 415482
rect 160296 413902 160678 413930
rect 170048 413902 170338 413930
rect 150544 413222 151018 413250
rect 150544 391814 150572 413222
rect 150532 391808 150584 391814
rect 150532 391750 150584 391756
rect 151004 391746 151032 394060
rect 160664 391746 160692 394060
rect 170324 393938 170352 394060
rect 170508 393938 170536 415550
rect 178408 415540 178460 415546
rect 178408 415482 178460 415488
rect 171784 415472 171836 415478
rect 171784 415414 171836 415420
rect 170324 393910 170536 393938
rect 171796 391746 171824 415414
rect 178420 413930 178448 415482
rect 187804 413930 187832 415550
rect 197452 415472 197504 415478
rect 197452 415414 197504 415420
rect 197464 413930 197492 415414
rect 178066 413902 178448 413930
rect 187726 413902 187832 413930
rect 197386 413902 197492 413930
rect 176566 403744 176622 403753
rect 176566 403679 176622 403688
rect 172518 403608 172574 403617
rect 172518 403543 172574 403552
rect 172532 394602 172560 403543
rect 176580 394602 176608 403679
rect 197556 394754 197584 415550
rect 200764 415540 200816 415546
rect 200764 415482 200816 415488
rect 199384 415472 199436 415478
rect 199384 415414 199436 415420
rect 197386 394726 197584 394754
rect 172520 394596 172572 394602
rect 172520 394538 172572 394544
rect 176568 394596 176620 394602
rect 176568 394538 176620 394544
rect 178052 391814 178080 394060
rect 187712 391814 187740 394060
rect 199396 391814 199424 415414
rect 200118 403608 200174 403617
rect 200118 403543 200174 403552
rect 200132 394670 200160 403543
rect 200120 394664 200172 394670
rect 200120 394606 200172 394612
rect 200776 391950 200804 415482
rect 214392 413930 214420 415550
rect 223948 415472 224000 415478
rect 223948 415414 224000 415420
rect 223960 413930 223988 415414
rect 214392 413902 214682 413930
rect 223960 413902 224342 413930
rect 204364 413222 205022 413250
rect 202786 404288 202842 404297
rect 202786 404223 202842 404232
rect 202800 394670 202828 404223
rect 202788 394664 202840 394670
rect 202788 394606 202840 394612
rect 200764 391944 200816 391950
rect 200764 391886 200816 391892
rect 204364 391814 204392 413222
rect 224512 394754 224540 415550
rect 232320 415540 232372 415546
rect 232320 415482 232372 415488
rect 225604 415472 225656 415478
rect 225604 415414 225656 415420
rect 224342 394726 224540 394754
rect 205008 391950 205036 394060
rect 204996 391944 205048 391950
rect 204996 391886 205048 391892
rect 178040 391808 178092 391814
rect 178040 391750 178092 391756
rect 187700 391808 187752 391814
rect 187700 391750 187752 391756
rect 199384 391808 199436 391814
rect 199384 391750 199436 391756
rect 204352 391808 204404 391814
rect 204352 391750 204404 391756
rect 214668 391746 214696 394060
rect 225616 391746 225644 415414
rect 232332 413930 232360 415482
rect 232070 413902 232360 413930
rect 241532 413930 241560 415550
rect 251180 415472 251232 415478
rect 251180 415414 251232 415420
rect 251192 413930 251220 415414
rect 241532 413902 241730 413930
rect 251192 413902 251390 413930
rect 230386 404288 230442 404297
rect 230386 404223 230442 404232
rect 226338 403608 226394 403617
rect 226338 403543 226394 403552
rect 226352 394602 226380 403543
rect 226340 394596 226392 394602
rect 226340 394538 226392 394544
rect 230400 394534 230428 404223
rect 251468 394754 251496 415550
rect 251824 415540 251876 415546
rect 251824 415482 251876 415488
rect 251390 394726 251496 394754
rect 230388 394528 230440 394534
rect 230388 394470 230440 394476
rect 232056 391814 232084 394060
rect 241716 391814 241744 394060
rect 251836 391950 251864 415482
rect 253204 415472 253256 415478
rect 253204 415414 253256 415420
rect 251824 391944 251876 391950
rect 251824 391886 251876 391892
rect 253216 391814 253244 415414
rect 268304 413930 268332 415550
rect 279516 415540 279568 415546
rect 279516 415482 279568 415488
rect 295800 415540 295852 415546
rect 295800 415482 295852 415488
rect 305644 415540 305696 415546
rect 305644 415482 305696 415488
rect 322388 415540 322440 415546
rect 322388 415482 322440 415488
rect 336004 415540 336056 415546
rect 336004 415482 336056 415488
rect 349804 415540 349856 415546
rect 349804 415482 349856 415488
rect 359648 415540 359700 415546
rect 359648 415482 359700 415488
rect 376300 415540 376352 415546
rect 376300 415482 376352 415488
rect 386512 415540 386564 415546
rect 386512 415482 386564 415488
rect 403348 415540 403400 415546
rect 403348 415482 403400 415488
rect 278044 415472 278096 415478
rect 278044 415414 278096 415420
rect 279424 415472 279476 415478
rect 279424 415414 279476 415420
rect 278056 413930 278084 415414
rect 268304 413902 268686 413930
rect 278056 413902 278346 413930
rect 258184 413222 259026 413250
rect 256606 404288 256662 404297
rect 256606 404223 256662 404232
rect 253938 403336 253994 403345
rect 253938 403271 253994 403280
rect 253952 394670 253980 403271
rect 253940 394664 253992 394670
rect 253940 394606 253992 394612
rect 256620 394602 256648 404223
rect 256608 394596 256660 394602
rect 256608 394538 256660 394544
rect 258184 391814 258212 413222
rect 278688 394664 278740 394670
rect 278346 394612 278688 394618
rect 278346 394606 278740 394612
rect 278346 394590 278728 394606
rect 259012 391950 259040 394060
rect 259000 391944 259052 391950
rect 259000 391886 259052 391892
rect 232044 391808 232096 391814
rect 232044 391750 232096 391756
rect 241704 391808 241756 391814
rect 241704 391750 241756 391756
rect 253204 391808 253256 391814
rect 253204 391750 253256 391756
rect 258172 391808 258224 391814
rect 258172 391750 258224 391756
rect 268672 391746 268700 394060
rect 279436 391746 279464 415414
rect 279528 394670 279556 415482
rect 285784 414038 286180 414066
rect 284206 403744 284262 403753
rect 284206 403679 284262 403688
rect 280158 403608 280214 403617
rect 280158 403543 280214 403552
rect 279516 394664 279568 394670
rect 279516 394606 279568 394612
rect 280172 394534 280200 403543
rect 284220 394670 284248 403679
rect 284208 394664 284260 394670
rect 284208 394606 284260 394612
rect 280160 394528 280212 394534
rect 280160 394470 280212 394476
rect 285784 391814 285812 414038
rect 286152 413930 286180 414038
rect 295812 413930 295840 415482
rect 305552 415472 305604 415478
rect 305552 415414 305604 415420
rect 305564 413930 305592 415414
rect 286074 413902 286180 413930
rect 295734 413902 295840 413930
rect 305394 413902 305592 413930
rect 305656 412634 305684 415482
rect 307024 415472 307076 415478
rect 307024 415414 307076 415420
rect 305472 412606 305684 412634
rect 305472 394754 305500 412606
rect 305394 394726 305500 394754
rect 285772 391808 285824 391814
rect 285772 391750 285824 391756
rect 286060 391746 286088 394060
rect 295720 391746 295748 394060
rect 307036 391746 307064 415414
rect 322400 413930 322428 415482
rect 331956 415472 332008 415478
rect 331956 415414 332008 415420
rect 333244 415472 333296 415478
rect 333244 415414 333296 415420
rect 331968 413930 331996 415414
rect 322400 413902 322690 413930
rect 331968 413902 332350 413930
rect 312004 413222 313030 413250
rect 311806 404288 311862 404297
rect 311806 404223 311862 404232
rect 307758 403608 307814 403617
rect 307758 403543 307814 403552
rect 307772 394602 307800 403543
rect 311820 394602 311848 404223
rect 307760 394596 307812 394602
rect 307760 394538 307812 394544
rect 311808 394596 311860 394602
rect 311808 394538 311860 394544
rect 312004 391746 312032 413222
rect 332600 394528 332652 394534
rect 332350 394476 332600 394482
rect 332350 394470 332652 394476
rect 332350 394454 332640 394470
rect 313016 391814 313044 394060
rect 313004 391808 313056 391814
rect 313004 391750 313056 391756
rect 322676 391746 322704 394060
rect 333256 391746 333284 415414
rect 335358 403608 335414 403617
rect 335358 403543 335414 403552
rect 335372 394670 335400 403543
rect 335360 394664 335412 394670
rect 335360 394606 335412 394612
rect 336016 394534 336044 415482
rect 349816 413930 349844 415482
rect 359464 415472 359516 415478
rect 359464 415414 359516 415420
rect 359476 413930 359504 415414
rect 349738 413902 349844 413930
rect 359398 413902 359504 413930
rect 359660 413658 359688 415482
rect 359740 415472 359792 415478
rect 359740 415414 359792 415420
rect 359476 413630 359688 413658
rect 340078 413370 340184 413386
rect 339592 413364 339644 413370
rect 340078 413364 340196 413370
rect 340078 413358 340144 413364
rect 339592 413306 339644 413312
rect 340144 413306 340196 413312
rect 338026 404288 338082 404297
rect 338026 404223 338082 404232
rect 338040 394670 338068 404223
rect 338028 394664 338080 394670
rect 338028 394606 338080 394612
rect 336004 394528 336056 394534
rect 336004 394470 336056 394476
rect 339604 391746 339632 413306
rect 359476 394754 359504 413630
rect 359752 412706 359780 415414
rect 376312 413930 376340 415482
rect 386052 415472 386104 415478
rect 386052 415414 386104 415420
rect 386064 413930 386092 415414
rect 376312 413902 376694 413930
rect 386064 413902 386354 413930
rect 359398 394726 359504 394754
rect 359568 412678 359780 412706
rect 365824 413222 367034 413250
rect 340064 391814 340092 394060
rect 340052 391808 340104 391814
rect 340052 391750 340104 391756
rect 349724 391746 349752 394060
rect 359568 391746 359596 412678
rect 365626 404288 365682 404297
rect 365626 404223 365682 404232
rect 361578 403336 361634 403345
rect 361578 403271 361634 403280
rect 361592 394602 361620 403271
rect 365640 394602 365668 404223
rect 361580 394596 361632 394602
rect 361580 394538 361632 394544
rect 365628 394596 365680 394602
rect 365628 394538 365680 394544
rect 365824 391746 365852 413222
rect 386524 394754 386552 415482
rect 387064 415472 387116 415478
rect 387064 415414 387116 415420
rect 386354 394726 386552 394754
rect 366744 394046 367034 394074
rect 366744 391814 366772 394046
rect 366732 391808 366784 391814
rect 366732 391750 366784 391756
rect 376680 391746 376708 394060
rect 387076 391746 387104 415414
rect 403360 413930 403388 415482
rect 412916 415472 412968 415478
rect 412916 415414 412968 415420
rect 412928 413930 412956 415414
rect 403360 413902 403650 413930
rect 412928 413902 413310 413930
rect 393424 413222 393990 413250
rect 391846 404288 391902 404297
rect 391846 404223 391902 404232
rect 389178 403608 389234 403617
rect 389178 403543 389234 403552
rect 389192 394670 389220 403543
rect 391860 394670 391888 404223
rect 389180 394664 389232 394670
rect 389180 394606 389232 394612
rect 391848 394664 391900 394670
rect 391848 394606 391900 394612
rect 393424 391746 393452 413222
rect 413480 394754 413508 415550
rect 421288 415540 421340 415546
rect 421288 415482 421340 415488
rect 414664 415472 414716 415478
rect 414664 415414 414716 415420
rect 413402 394726 413508 394754
rect 393976 391814 394004 394060
rect 393964 391808 394016 391814
rect 393964 391750 394016 391756
rect 403728 391746 403756 394060
rect 414676 391746 414704 415414
rect 421300 413930 421328 415482
rect 421038 413902 421328 413930
rect 430592 413930 430620 415550
rect 440240 415472 440292 415478
rect 440240 415414 440292 415420
rect 440252 413930 440280 415414
rect 430592 413902 430698 413930
rect 440252 413902 440358 413930
rect 419446 404288 419502 404297
rect 419446 404223 419502 404232
rect 415398 403608 415454 403617
rect 415398 403543 415454 403552
rect 415412 394602 415440 403543
rect 419460 394602 419488 404223
rect 440528 394754 440556 415550
rect 445024 415540 445076 415546
rect 445024 415482 445076 415488
rect 442264 415472 442316 415478
rect 442264 415414 442316 415420
rect 440358 394726 440556 394754
rect 415400 394596 415452 394602
rect 415400 394538 415452 394544
rect 419448 394596 419500 394602
rect 419448 394538 419500 394544
rect 421024 391814 421052 394060
rect 430684 391814 430712 394060
rect 442276 391814 442304 415414
rect 442998 403608 443054 403617
rect 442998 403543 443054 403552
rect 443012 394670 443040 403543
rect 445036 394738 445064 415482
rect 457272 413930 457300 415550
rect 467012 415472 467064 415478
rect 467012 415414 467064 415420
rect 468484 415472 468536 415478
rect 468484 415414 468536 415420
rect 467024 413930 467052 415414
rect 457272 413902 457654 413930
rect 467024 413902 467314 413930
rect 447244 413222 447994 413250
rect 445666 404288 445722 404297
rect 445666 404223 445722 404232
rect 445024 394732 445076 394738
rect 445024 394674 445076 394680
rect 445680 394670 445708 404223
rect 443000 394664 443052 394670
rect 443000 394606 443052 394612
rect 445668 394664 445720 394670
rect 445668 394606 445720 394612
rect 447244 391814 447272 413222
rect 447692 394732 447744 394738
rect 447692 394674 447744 394680
rect 447704 394618 447732 394674
rect 447704 394590 447994 394618
rect 467406 394602 467696 394618
rect 467406 394596 467708 394602
rect 467406 394590 467656 394596
rect 467656 394538 467708 394544
rect 421012 391808 421064 391814
rect 421012 391750 421064 391756
rect 430672 391808 430724 391814
rect 430672 391750 430724 391756
rect 442264 391808 442316 391814
rect 442264 391750 442316 391756
rect 447232 391808 447284 391814
rect 447232 391750 447284 391756
rect 457732 391746 457760 394060
rect 468496 391746 468524 415414
rect 468588 394602 468616 415550
rect 475396 413930 475424 415618
rect 484400 415608 484452 415614
rect 484400 415550 484452 415556
rect 475042 413902 475424 413930
rect 484412 413930 484440 415550
rect 494520 415540 494572 415546
rect 494520 415482 494572 415488
rect 494060 415472 494112 415478
rect 494060 415414 494112 415420
rect 494072 413930 494100 415414
rect 484412 413902 484702 413930
rect 494072 413902 494362 413930
rect 473266 403744 473322 403753
rect 473266 403679 473322 403688
rect 469218 403336 469274 403345
rect 469218 403271 469274 403280
rect 468576 394596 468628 394602
rect 468576 394538 468628 394544
rect 469232 394534 469260 403271
rect 473280 394602 473308 403679
rect 494532 394754 494560 415482
rect 494362 394726 494560 394754
rect 473268 394596 473320 394602
rect 473268 394538 473320 394544
rect 469220 394528 469272 394534
rect 469220 394470 469272 394476
rect 475028 391814 475056 394060
rect 484688 391814 484716 394060
rect 494716 391950 494744 415618
rect 511356 415540 511408 415546
rect 511356 415482 511408 415488
rect 522304 415540 522356 415546
rect 522304 415482 522356 415488
rect 496084 415472 496136 415478
rect 496084 415414 496136 415420
rect 494704 391944 494756 391950
rect 494704 391886 494756 391892
rect 496096 391814 496124 415414
rect 511368 413930 511396 415482
rect 520924 415472 520976 415478
rect 520924 415414 520976 415420
rect 520936 413930 520964 415414
rect 511368 413902 511658 413930
rect 520936 413902 521318 413930
rect 501064 413222 501998 413250
rect 500866 404288 500922 404297
rect 500866 404223 500922 404232
rect 496818 403608 496874 403617
rect 496818 403543 496874 403552
rect 496832 394670 496860 403543
rect 500880 394670 500908 404223
rect 496820 394664 496872 394670
rect 496820 394606 496872 394612
rect 500868 394664 500920 394670
rect 500868 394606 500920 394612
rect 501064 391814 501092 413222
rect 522316 402974 522344 415482
rect 522396 415472 522448 415478
rect 522396 415414 522448 415420
rect 521856 402946 522344 402974
rect 521856 394618 521884 402946
rect 521410 394590 521884 394618
rect 501984 391950 502012 394060
rect 501972 391944 502024 391950
rect 501972 391886 502024 391892
rect 475016 391808 475068 391814
rect 475016 391750 475068 391756
rect 484676 391808 484728 391814
rect 484676 391750 484728 391756
rect 496084 391808 496136 391814
rect 496084 391750 496136 391756
rect 501052 391808 501104 391814
rect 501052 391750 501104 391756
rect 511736 391746 511764 394060
rect 522408 391746 522436 415414
rect 526444 414724 526496 414730
rect 526444 414666 526496 414672
rect 526456 404297 526484 414666
rect 528756 413930 528784 416026
rect 538404 415540 538456 415546
rect 538404 415482 538456 415488
rect 538416 413930 538444 415482
rect 548064 415472 548116 415478
rect 548064 415414 548116 415420
rect 548076 413930 548104 415414
rect 528756 413902 529046 413930
rect 538416 413902 538706 413930
rect 548076 413902 548366 413930
rect 526442 404288 526498 404297
rect 526442 404223 526498 404232
rect 523038 403608 523094 403617
rect 523038 403543 523094 403552
rect 550638 403608 550694 403617
rect 550638 403543 550694 403552
rect 523052 394602 523080 403543
rect 550652 394670 550680 403543
rect 550640 394664 550692 394670
rect 550640 394606 550692 394612
rect 523040 394596 523092 394602
rect 523040 394538 523092 394544
rect 529032 391814 529060 394060
rect 529020 391808 529072 391814
rect 529020 391750 529072 391756
rect 150992 391740 151044 391746
rect 150992 391682 151044 391688
rect 160652 391740 160704 391746
rect 160652 391682 160704 391688
rect 171784 391740 171836 391746
rect 171784 391682 171836 391688
rect 214656 391740 214708 391746
rect 214656 391682 214708 391688
rect 225604 391740 225656 391746
rect 225604 391682 225656 391688
rect 268660 391740 268712 391746
rect 268660 391682 268712 391688
rect 279424 391740 279476 391746
rect 279424 391682 279476 391688
rect 286048 391740 286100 391746
rect 286048 391682 286100 391688
rect 295708 391740 295760 391746
rect 295708 391682 295760 391688
rect 307024 391740 307076 391746
rect 307024 391682 307076 391688
rect 311992 391740 312044 391746
rect 311992 391682 312044 391688
rect 322664 391740 322716 391746
rect 322664 391682 322716 391688
rect 333244 391740 333296 391746
rect 333244 391682 333296 391688
rect 339592 391740 339644 391746
rect 339592 391682 339644 391688
rect 349712 391740 349764 391746
rect 349712 391682 349764 391688
rect 359556 391740 359608 391746
rect 359556 391682 359608 391688
rect 365812 391740 365864 391746
rect 365812 391682 365864 391688
rect 376668 391740 376720 391746
rect 376668 391682 376720 391688
rect 387064 391740 387116 391746
rect 387064 391682 387116 391688
rect 393412 391740 393464 391746
rect 393412 391682 393464 391688
rect 403716 391740 403768 391746
rect 403716 391682 403768 391688
rect 414664 391740 414716 391746
rect 414664 391682 414716 391688
rect 457720 391740 457772 391746
rect 457720 391682 457772 391688
rect 468484 391740 468536 391746
rect 468484 391682 468536 391688
rect 511724 391740 511776 391746
rect 511724 391682 511776 391688
rect 522396 391740 522448 391746
rect 522396 391682 522448 391688
rect 538692 391678 538720 394060
rect 548352 391882 548380 394060
rect 548340 391876 548392 391882
rect 548340 391818 548392 391824
rect 538680 391672 538732 391678
rect 538680 391614 538732 391620
rect 528744 389836 528796 389842
rect 528744 389778 528796 389784
rect 232320 389428 232372 389434
rect 232320 389370 232372 389376
rect 251824 389428 251876 389434
rect 251824 389370 251876 389376
rect 475384 389428 475436 389434
rect 475384 389370 475436 389376
rect 494704 389428 494756 389434
rect 494704 389370 494756 389376
rect 170496 389360 170548 389366
rect 170496 389302 170548 389308
rect 187792 389360 187844 389366
rect 187792 389302 187844 389308
rect 197544 389360 197596 389366
rect 197544 389302 197596 389308
rect 214380 389360 214432 389366
rect 214380 389302 214432 389308
rect 224500 389360 224552 389366
rect 224500 389302 224552 389308
rect 170036 389292 170088 389298
rect 170036 389234 170088 389240
rect 160284 389224 160336 389230
rect 160284 389166 160336 389172
rect 160296 386866 160324 389166
rect 170048 386866 170076 389234
rect 160296 386838 160678 386866
rect 170048 386838 170338 386866
rect 150636 386294 151018 386322
rect 150636 373994 150664 386294
rect 150544 373966 150664 373994
rect 149704 365628 149756 365634
rect 149704 365570 149756 365576
rect 150544 365566 150572 373966
rect 170232 367674 170338 367690
rect 170508 367674 170536 389302
rect 178408 389292 178460 389298
rect 178408 389234 178460 389240
rect 171784 389224 171836 389230
rect 171784 389166 171836 389172
rect 170220 367668 170338 367674
rect 170272 367662 170338 367668
rect 170496 367668 170548 367674
rect 170220 367610 170272 367616
rect 170496 367610 170548 367616
rect 150728 367118 151018 367146
rect 160572 367118 160678 367146
rect 150532 365560 150584 365566
rect 150532 365502 150584 365508
rect 150728 365498 150756 367118
rect 160572 365498 160600 367118
rect 171796 365498 171824 389166
rect 178420 386866 178448 389234
rect 187804 386866 187832 389302
rect 197452 389224 197504 389230
rect 197452 389166 197504 389172
rect 197464 386866 197492 389166
rect 178066 386838 178448 386866
rect 187726 386838 187832 386866
rect 197386 386838 197492 386866
rect 176566 376816 176622 376825
rect 176566 376751 176622 376760
rect 172518 376544 172574 376553
rect 172518 376479 172574 376488
rect 172532 368422 172560 376479
rect 176580 368422 176608 376751
rect 197556 373994 197584 389302
rect 200764 389292 200816 389298
rect 200764 389234 200816 389240
rect 199384 389224 199436 389230
rect 199384 389166 199436 389172
rect 197464 373966 197584 373994
rect 172520 368416 172572 368422
rect 172520 368358 172572 368364
rect 176568 368416 176620 368422
rect 176568 368358 176620 368364
rect 197464 367690 197492 373966
rect 197386 367662 197492 367690
rect 178066 367118 178172 367146
rect 187726 367118 188016 367146
rect 178144 365566 178172 367118
rect 187988 365566 188016 367118
rect 199396 365566 199424 389166
rect 200118 376544 200174 376553
rect 200118 376479 200174 376488
rect 200132 368490 200160 376479
rect 200120 368484 200172 368490
rect 200120 368426 200172 368432
rect 200776 365702 200804 389234
rect 214392 386866 214420 389302
rect 223948 389224 224000 389230
rect 223948 389166 224000 389172
rect 223960 386866 223988 389166
rect 214392 386838 214682 386866
rect 223960 386838 224342 386866
rect 204548 386294 205022 386322
rect 202786 377224 202842 377233
rect 202786 377159 202842 377168
rect 202800 368490 202828 377159
rect 204548 373994 204576 386294
rect 204364 373966 204576 373994
rect 202788 368484 202840 368490
rect 202788 368426 202840 368432
rect 200764 365696 200816 365702
rect 200764 365638 200816 365644
rect 204364 365566 204392 373966
rect 224512 367690 224540 389302
rect 225604 389224 225656 389230
rect 225604 389166 225656 389172
rect 224342 367662 224540 367690
rect 204640 367118 205022 367146
rect 214682 367118 215064 367146
rect 204640 365702 204668 367118
rect 204628 365696 204680 365702
rect 204628 365638 204680 365644
rect 178132 365560 178184 365566
rect 178132 365502 178184 365508
rect 187976 365560 188028 365566
rect 187976 365502 188028 365508
rect 199384 365560 199436 365566
rect 199384 365502 199436 365508
rect 204352 365560 204404 365566
rect 204352 365502 204404 365508
rect 215036 365498 215064 367118
rect 225616 365498 225644 389166
rect 232332 386866 232360 389370
rect 241520 389360 241572 389366
rect 241520 389302 241572 389308
rect 232070 386838 232360 386866
rect 241532 386866 241560 389302
rect 251456 389292 251508 389298
rect 251456 389234 251508 389240
rect 251180 389224 251232 389230
rect 251180 389166 251232 389172
rect 251192 386866 251220 389166
rect 241532 386838 241730 386866
rect 251192 386838 251390 386866
rect 230386 377224 230442 377233
rect 230386 377159 230442 377168
rect 226338 376544 226394 376553
rect 226338 376479 226394 376488
rect 226352 368422 226380 376479
rect 226340 368416 226392 368422
rect 226340 368358 226392 368364
rect 230400 368354 230428 377159
rect 230388 368348 230440 368354
rect 230388 368290 230440 368296
rect 251468 367690 251496 389234
rect 251390 367662 251496 367690
rect 231872 367118 232070 367146
rect 241730 367118 242112 367146
rect 231872 365566 231900 367118
rect 242084 365566 242112 367118
rect 251836 365702 251864 389370
rect 413468 389360 413520 389366
rect 413468 389302 413520 389308
rect 430580 389360 430632 389366
rect 430580 389302 430632 389308
rect 440516 389360 440568 389366
rect 440516 389302 440568 389308
rect 457260 389360 457312 389366
rect 457260 389302 457312 389308
rect 468576 389360 468628 389366
rect 468576 389302 468628 389308
rect 268292 389292 268344 389298
rect 268292 389234 268344 389240
rect 279424 389292 279476 389298
rect 279424 389234 279476 389240
rect 295800 389292 295852 389298
rect 295800 389234 295852 389240
rect 305644 389292 305696 389298
rect 305644 389234 305696 389240
rect 322388 389292 322440 389298
rect 322388 389234 322440 389240
rect 336004 389292 336056 389298
rect 336004 389234 336056 389240
rect 349804 389292 349856 389298
rect 349804 389234 349856 389240
rect 359556 389292 359608 389298
rect 359556 389234 359608 389240
rect 376300 389292 376352 389298
rect 376300 389234 376352 389240
rect 386512 389292 386564 389298
rect 386512 389234 386564 389240
rect 403348 389292 403400 389298
rect 403348 389234 403400 389240
rect 253204 389224 253256 389230
rect 253204 389166 253256 389172
rect 251824 365696 251876 365702
rect 251824 365638 251876 365644
rect 253216 365566 253244 389166
rect 268304 386866 268332 389234
rect 278044 389224 278096 389230
rect 278044 389166 278096 389172
rect 278056 386866 278084 389166
rect 268304 386838 268686 386866
rect 278056 386838 278346 386866
rect 258644 386294 259026 386322
rect 256606 377224 256662 377233
rect 256606 377159 256662 377168
rect 253938 376000 253994 376009
rect 253938 375935 253994 375944
rect 253952 368490 253980 375935
rect 253940 368484 253992 368490
rect 253940 368426 253992 368432
rect 256620 368422 256648 377159
rect 258644 373994 258672 386294
rect 279436 373994 279464 389234
rect 279516 389224 279568 389230
rect 279516 389166 279568 389172
rect 258184 373966 258672 373994
rect 278792 373966 279464 373994
rect 256608 368416 256660 368422
rect 256608 368358 256660 368364
rect 258184 365566 258212 373966
rect 278792 367690 278820 373966
rect 278346 367662 278820 367690
rect 258736 367118 259026 367146
rect 268686 367118 268976 367146
rect 258736 365702 258764 367118
rect 258724 365696 258776 365702
rect 258724 365638 258776 365644
rect 231860 365560 231912 365566
rect 231860 365502 231912 365508
rect 242072 365560 242124 365566
rect 242072 365502 242124 365508
rect 253204 365560 253256 365566
rect 253204 365502 253256 365508
rect 258172 365560 258224 365566
rect 258172 365502 258224 365508
rect 268948 365498 268976 367118
rect 279528 365498 279556 389166
rect 295812 386866 295840 389234
rect 305552 389224 305604 389230
rect 305552 389166 305604 389172
rect 305564 386866 305592 389166
rect 295734 386838 295840 386866
rect 305394 386838 305592 386866
rect 286074 386306 286180 386322
rect 285772 386300 285824 386306
rect 286074 386300 286192 386306
rect 286074 386294 286140 386300
rect 285772 386242 285824 386248
rect 286140 386242 286192 386248
rect 284206 376816 284262 376825
rect 284206 376751 284262 376760
rect 280158 376544 280214 376553
rect 280158 376479 280214 376488
rect 280172 368354 280200 376479
rect 284220 368490 284248 376751
rect 284208 368484 284260 368490
rect 284208 368426 284260 368432
rect 280160 368348 280212 368354
rect 280160 368290 280212 368296
rect 285784 365498 285812 386242
rect 305656 373994 305684 389234
rect 307024 389224 307076 389230
rect 307024 389166 307076 389172
rect 305472 373966 305684 373994
rect 305472 367690 305500 373966
rect 305394 367662 305500 367690
rect 286074 367118 286180 367146
rect 295734 367118 296024 367146
rect 286152 365566 286180 367118
rect 286140 365560 286192 365566
rect 286140 365502 286192 365508
rect 295996 365498 296024 367118
rect 307036 365498 307064 389166
rect 322400 386866 322428 389234
rect 331956 389224 332008 389230
rect 331956 389166 332008 389172
rect 333244 389224 333296 389230
rect 333244 389166 333296 389172
rect 331968 386866 331996 389166
rect 322400 386838 322690 386866
rect 331968 386838 332350 386866
rect 312556 386294 313030 386322
rect 311806 377224 311862 377233
rect 311806 377159 311862 377168
rect 307758 376544 307814 376553
rect 307758 376479 307814 376488
rect 307772 368422 307800 376479
rect 311820 368422 311848 377159
rect 312556 373994 312584 386294
rect 312004 373966 312584 373994
rect 307760 368416 307812 368422
rect 307760 368358 307812 368364
rect 311808 368416 311860 368422
rect 311808 368358 311860 368364
rect 312004 365498 312032 373966
rect 312648 367118 313030 367146
rect 322690 367118 322888 367146
rect 332350 367118 332548 367146
rect 312648 365566 312676 367118
rect 312636 365560 312688 365566
rect 312636 365502 312688 365508
rect 322860 365498 322888 367118
rect 332520 365702 332548 367118
rect 332508 365696 332560 365702
rect 332508 365638 332560 365644
rect 333256 365498 333284 389166
rect 335358 376544 335414 376553
rect 335358 376479 335414 376488
rect 335372 368490 335400 376479
rect 335360 368484 335412 368490
rect 335360 368426 335412 368432
rect 336016 365702 336044 389234
rect 349816 386866 349844 389234
rect 359464 389224 359516 389230
rect 359464 389166 359516 389172
rect 359476 386866 359504 389166
rect 349738 386838 349844 386866
rect 359398 386838 359504 386866
rect 359568 386594 359596 389234
rect 359740 389224 359792 389230
rect 359740 389166 359792 389172
rect 359476 386566 359596 386594
rect 340078 386306 340184 386322
rect 339592 386300 339644 386306
rect 340078 386300 340196 386306
rect 340078 386294 340144 386300
rect 339592 386242 339644 386248
rect 340144 386242 340196 386248
rect 338026 377224 338082 377233
rect 338026 377159 338082 377168
rect 338040 368490 338068 377159
rect 338028 368484 338080 368490
rect 338028 368426 338080 368432
rect 336004 365696 336056 365702
rect 336004 365638 336056 365644
rect 339604 365498 339632 386242
rect 359476 367690 359504 386566
rect 359752 386322 359780 389166
rect 376312 386866 376340 389234
rect 386052 389224 386104 389230
rect 386052 389166 386104 389172
rect 386064 386866 386092 389166
rect 376312 386838 376694 386866
rect 386064 386838 386354 386866
rect 359398 367662 359504 367690
rect 359568 386294 359780 386322
rect 366652 386294 367034 386322
rect 340078 367118 340184 367146
rect 349738 367118 350120 367146
rect 340156 365566 340184 367118
rect 340144 365560 340196 365566
rect 340144 365502 340196 365508
rect 350092 365498 350120 367118
rect 359568 365498 359596 386294
rect 365626 377224 365682 377233
rect 365626 377159 365682 377168
rect 361578 376000 361634 376009
rect 361578 375935 361634 375944
rect 361592 368422 361620 375935
rect 365640 368422 365668 377159
rect 366652 373994 366680 386294
rect 365824 373966 366680 373994
rect 361580 368416 361632 368422
rect 361580 368358 361632 368364
rect 365628 368416 365680 368422
rect 365628 368358 365680 368364
rect 365824 365498 365852 373966
rect 386524 367690 386552 389234
rect 387064 389224 387116 389230
rect 387064 389166 387116 389172
rect 386354 367662 386552 367690
rect 366744 367118 367034 367146
rect 376588 367118 376694 367146
rect 366744 365566 366772 367118
rect 366732 365560 366784 365566
rect 366732 365502 366784 365508
rect 376588 365498 376616 367118
rect 387076 365498 387104 389166
rect 403360 386866 403388 389234
rect 412916 389224 412968 389230
rect 412916 389166 412968 389172
rect 412928 386866 412956 389166
rect 403360 386838 403650 386866
rect 412928 386838 413310 386866
rect 393424 386294 393990 386322
rect 391846 377224 391902 377233
rect 391846 377159 391902 377168
rect 389178 376544 389234 376553
rect 389178 376479 389234 376488
rect 389192 368490 389220 376479
rect 391860 368490 391888 377159
rect 389180 368484 389232 368490
rect 389180 368426 389232 368432
rect 391848 368484 391900 368490
rect 391848 368426 391900 368432
rect 393424 365498 393452 386294
rect 413480 367690 413508 389302
rect 421288 389292 421340 389298
rect 421288 389234 421340 389240
rect 414664 389224 414716 389230
rect 414664 389166 414716 389172
rect 413402 367662 413508 367690
rect 393608 367118 393990 367146
rect 403742 367118 404032 367146
rect 393608 365566 393636 367118
rect 393596 365560 393648 365566
rect 393596 365502 393648 365508
rect 404004 365498 404032 367118
rect 414676 365498 414704 389166
rect 421300 386866 421328 389234
rect 421038 386838 421328 386866
rect 430592 386866 430620 389302
rect 440240 389224 440292 389230
rect 440240 389166 440292 389172
rect 440252 386866 440280 389166
rect 430592 386838 430698 386866
rect 440252 386838 440358 386866
rect 419446 377224 419502 377233
rect 419446 377159 419502 377168
rect 415398 376544 415454 376553
rect 415398 376479 415454 376488
rect 415412 368422 415440 376479
rect 419460 368422 419488 377159
rect 415400 368416 415452 368422
rect 415400 368358 415452 368364
rect 419448 368416 419500 368422
rect 419448 368358 419500 368364
rect 440528 367690 440556 389302
rect 446404 389292 446456 389298
rect 446404 389234 446456 389240
rect 442264 389224 442316 389230
rect 442264 389166 442316 389172
rect 440358 367662 440556 367690
rect 420932 367118 421038 367146
rect 430698 367118 431080 367146
rect 420932 365566 420960 367118
rect 431052 365566 431080 367118
rect 442276 365566 442304 389166
rect 445666 377224 445722 377233
rect 445666 377159 445722 377168
rect 442998 376544 443054 376553
rect 442998 376479 443054 376488
rect 443012 368490 443040 376479
rect 443000 368484 443052 368490
rect 443000 368426 443052 368432
rect 445680 368354 445708 377159
rect 446416 368490 446444 389234
rect 457272 386866 457300 389302
rect 467012 389224 467064 389230
rect 467012 389166 467064 389172
rect 468484 389224 468536 389230
rect 468484 389166 468536 389172
rect 467024 386866 467052 389166
rect 457272 386838 457654 386866
rect 467024 386838 467314 386866
rect 447244 386294 447994 386322
rect 446404 368484 446456 368490
rect 446404 368426 446456 368432
rect 445668 368348 445720 368354
rect 445668 368290 445720 368296
rect 447244 365566 447272 386294
rect 447692 368484 447744 368490
rect 447692 368426 447744 368432
rect 447704 367690 447732 368426
rect 467656 368348 467708 368354
rect 467656 368290 467708 368296
rect 467668 367690 467696 368290
rect 447704 367662 447994 367690
rect 467406 367662 467696 367690
rect 457746 367118 458128 367146
rect 420920 365560 420972 365566
rect 420920 365502 420972 365508
rect 431040 365560 431092 365566
rect 431040 365502 431092 365508
rect 442264 365560 442316 365566
rect 442264 365502 442316 365508
rect 447232 365560 447284 365566
rect 447232 365502 447284 365508
rect 458100 365498 458128 367118
rect 468496 365498 468524 389166
rect 468588 368354 468616 389302
rect 475396 386866 475424 389370
rect 484400 389360 484452 389366
rect 484400 389302 484452 389308
rect 475042 386838 475424 386866
rect 484412 386866 484440 389302
rect 494520 389292 494572 389298
rect 494520 389234 494572 389240
rect 494060 389224 494112 389230
rect 494060 389166 494112 389172
rect 494072 386866 494100 389166
rect 484412 386838 484702 386866
rect 494072 386838 494362 386866
rect 473266 376816 473322 376825
rect 473266 376751 473322 376760
rect 469218 376000 469274 376009
rect 469218 375935 469274 375944
rect 469232 368422 469260 375935
rect 473280 368422 473308 376751
rect 469220 368416 469272 368422
rect 469220 368358 469272 368364
rect 473268 368416 473320 368422
rect 473268 368358 473320 368364
rect 468576 368348 468628 368354
rect 468576 368290 468628 368296
rect 494532 367690 494560 389234
rect 494362 367662 494560 367690
rect 474752 367118 475042 367146
rect 484702 367118 484992 367146
rect 474752 365566 474780 367118
rect 484964 365566 484992 367118
rect 494716 365702 494744 389370
rect 511356 389292 511408 389298
rect 511356 389234 511408 389240
rect 522304 389292 522356 389298
rect 522304 389234 522356 389240
rect 496084 389224 496136 389230
rect 496084 389166 496136 389172
rect 494704 365696 494756 365702
rect 494704 365638 494756 365644
rect 496096 365566 496124 389166
rect 511368 386866 511396 389234
rect 520924 389224 520976 389230
rect 520924 389166 520976 389172
rect 520936 386866 520964 389166
rect 511368 386838 511658 386866
rect 520936 386838 521318 386866
rect 501064 386294 501998 386322
rect 500866 377224 500922 377233
rect 500866 377159 500922 377168
rect 496818 376544 496874 376553
rect 496818 376479 496874 376488
rect 496832 368490 496860 376479
rect 500880 368490 500908 377159
rect 496820 368484 496872 368490
rect 496820 368426 496872 368432
rect 500868 368484 500920 368490
rect 500868 368426 500920 368432
rect 501064 365566 501092 386294
rect 522316 373994 522344 389234
rect 522396 389224 522448 389230
rect 522396 389166 522448 389172
rect 521856 373966 522344 373994
rect 521856 367690 521884 373966
rect 521410 367662 521884 367690
rect 501616 367118 501998 367146
rect 511750 367118 511948 367146
rect 501616 365702 501644 367118
rect 501604 365696 501656 365702
rect 501604 365638 501656 365644
rect 474740 365560 474792 365566
rect 474740 365502 474792 365508
rect 484952 365560 485004 365566
rect 484952 365502 485004 365508
rect 496084 365560 496136 365566
rect 496084 365502 496136 365508
rect 501052 365560 501104 365566
rect 501052 365502 501104 365508
rect 511920 365498 511948 367118
rect 522408 365498 522436 389166
rect 526444 387116 526496 387122
rect 526444 387058 526496 387064
rect 526456 377369 526484 387058
rect 528756 386866 528784 389778
rect 538404 389292 538456 389298
rect 538404 389234 538456 389240
rect 538416 386866 538444 389234
rect 548064 389224 548116 389230
rect 548064 389166 548116 389172
rect 548076 386866 548104 389166
rect 528756 386838 529046 386866
rect 538416 386838 538706 386866
rect 548076 386838 548366 386866
rect 526442 377360 526498 377369
rect 526442 377295 526498 377304
rect 523038 376544 523094 376553
rect 523038 376479 523094 376488
rect 550638 376544 550694 376553
rect 550638 376479 550694 376488
rect 523052 368422 523080 376479
rect 550652 368490 550680 376479
rect 550640 368484 550692 368490
rect 550640 368426 550692 368432
rect 523040 368416 523092 368422
rect 523040 368358 523092 368364
rect 528664 367118 529046 367146
rect 538416 367118 538706 367146
rect 548076 367118 548366 367146
rect 528664 365566 528692 367118
rect 528652 365560 528704 365566
rect 528652 365502 528704 365508
rect 150716 365492 150768 365498
rect 150716 365434 150768 365440
rect 160560 365492 160612 365498
rect 160560 365434 160612 365440
rect 171784 365492 171836 365498
rect 171784 365434 171836 365440
rect 215024 365492 215076 365498
rect 215024 365434 215076 365440
rect 225604 365492 225656 365498
rect 225604 365434 225656 365440
rect 268936 365492 268988 365498
rect 268936 365434 268988 365440
rect 279516 365492 279568 365498
rect 279516 365434 279568 365440
rect 285772 365492 285824 365498
rect 285772 365434 285824 365440
rect 295984 365492 296036 365498
rect 295984 365434 296036 365440
rect 307024 365492 307076 365498
rect 307024 365434 307076 365440
rect 311992 365492 312044 365498
rect 311992 365434 312044 365440
rect 322848 365492 322900 365498
rect 322848 365434 322900 365440
rect 333244 365492 333296 365498
rect 333244 365434 333296 365440
rect 339592 365492 339644 365498
rect 339592 365434 339644 365440
rect 350080 365492 350132 365498
rect 350080 365434 350132 365440
rect 359556 365492 359608 365498
rect 359556 365434 359608 365440
rect 365812 365492 365864 365498
rect 365812 365434 365864 365440
rect 376576 365492 376628 365498
rect 376576 365434 376628 365440
rect 387064 365492 387116 365498
rect 387064 365434 387116 365440
rect 393412 365492 393464 365498
rect 393412 365434 393464 365440
rect 403992 365492 404044 365498
rect 403992 365434 404044 365440
rect 414664 365492 414716 365498
rect 414664 365434 414716 365440
rect 458088 365492 458140 365498
rect 458088 365434 458140 365440
rect 468484 365492 468536 365498
rect 468484 365434 468536 365440
rect 511908 365492 511960 365498
rect 511908 365434 511960 365440
rect 522396 365492 522448 365498
rect 522396 365434 522448 365440
rect 538416 365430 538444 367118
rect 548076 365634 548104 367118
rect 548064 365628 548116 365634
rect 548064 365570 548116 365576
rect 538404 365424 538456 365430
rect 538404 365366 538456 365372
rect 529020 362228 529072 362234
rect 529020 362170 529072 362176
rect 149704 361888 149756 361894
rect 149704 361830 149756 361836
rect 148966 350296 149022 350305
rect 148966 350231 149022 350240
rect 148980 340882 149008 350231
rect 148968 340876 149020 340882
rect 148968 340818 149020 340824
rect 146944 338088 146996 338094
rect 146944 338030 146996 338036
rect 124036 338020 124088 338026
rect 124036 337962 124088 337968
rect 133696 338020 133748 338026
rect 133696 337962 133748 337968
rect 144184 338020 144236 338026
rect 144184 337962 144236 337968
rect 79692 337952 79744 337958
rect 79692 337894 79744 337900
rect 90456 337952 90508 337958
rect 90456 337894 90508 337900
rect 106648 337952 106700 337958
rect 106648 337894 106700 337900
rect 116584 337952 116636 337958
rect 116584 337894 116636 337900
rect 122932 337952 122984 337958
rect 122932 337894 122984 337900
rect 146944 335640 146996 335646
rect 146944 335582 146996 335588
rect 52460 335572 52512 335578
rect 52460 335514 52512 335520
rect 43352 335368 43404 335374
rect 43352 335310 43404 335316
rect 37924 333260 37976 333266
rect 37924 333202 37976 333208
rect 43364 332874 43392 335310
rect 43102 332846 43392 332874
rect 52472 332874 52500 335514
rect 62488 335504 62540 335510
rect 62488 335446 62540 335452
rect 79324 335504 79376 335510
rect 79324 335446 79376 335452
rect 90456 335504 90508 335510
rect 90456 335446 90508 335452
rect 106464 335504 106516 335510
rect 106464 335446 106516 335452
rect 116492 335504 116544 335510
rect 116492 335446 116544 335452
rect 133420 335504 133472 335510
rect 133420 335446 133472 335452
rect 62120 335436 62172 335442
rect 62120 335378 62172 335384
rect 62132 332874 62160 335378
rect 52472 332846 52670 332874
rect 62132 332846 62330 332874
rect 41326 323232 41382 323241
rect 41326 323167 41382 323176
rect 37922 322008 37978 322017
rect 37922 321943 37978 321952
rect 36820 311704 36872 311710
rect 36820 311646 36872 311652
rect 36728 311568 36780 311574
rect 36728 311510 36780 311516
rect 36820 308032 36872 308038
rect 36820 307974 36872 307980
rect 36728 307896 36780 307902
rect 36728 307838 36780 307844
rect 36740 284170 36768 307838
rect 36832 286958 36860 307974
rect 37936 305658 37964 321943
rect 41340 314566 41368 323167
rect 41328 314560 41380 314566
rect 41328 314502 41380 314508
rect 62500 313698 62528 335446
rect 64144 335436 64196 335442
rect 64144 335378 64196 335384
rect 62764 335368 62816 335374
rect 62764 335310 62816 335316
rect 62422 313670 62528 313698
rect 42812 313126 43010 313154
rect 52762 313126 53144 313154
rect 42812 311778 42840 313126
rect 53116 311778 53144 313126
rect 62776 311846 62804 335310
rect 62764 311840 62816 311846
rect 62764 311782 62816 311788
rect 64156 311778 64184 335378
rect 79336 332874 79364 335446
rect 89076 335436 89128 335442
rect 89076 335378 89128 335384
rect 90364 335436 90416 335442
rect 90364 335378 90416 335384
rect 89088 332874 89116 335378
rect 79336 332846 79718 332874
rect 89088 332846 89378 332874
rect 69124 332302 70058 332330
rect 68926 322960 68982 322969
rect 68926 322895 68982 322904
rect 64878 322552 64934 322561
rect 64878 322487 64934 322496
rect 64892 314634 64920 322487
rect 64880 314628 64932 314634
rect 64880 314570 64932 314576
rect 68940 314498 68968 322895
rect 68928 314492 68980 314498
rect 68928 314434 68980 314440
rect 69124 311778 69152 332302
rect 89720 314628 89772 314634
rect 89720 314570 89772 314576
rect 89732 313698 89760 314570
rect 89378 313670 89760 313698
rect 69768 313126 70058 313154
rect 79718 313126 80008 313154
rect 69768 311846 69796 313126
rect 69756 311840 69808 311846
rect 69756 311782 69808 311788
rect 42800 311772 42852 311778
rect 42800 311714 42852 311720
rect 53104 311772 53156 311778
rect 53104 311714 53156 311720
rect 64144 311772 64196 311778
rect 64144 311714 64196 311720
rect 69112 311772 69164 311778
rect 69112 311714 69164 311720
rect 79980 311710 80008 313126
rect 90376 311710 90404 335378
rect 90468 314634 90496 335446
rect 106476 332874 106504 335446
rect 116124 335436 116176 335442
rect 116124 335378 116176 335384
rect 116136 332874 116164 335378
rect 106476 332846 106674 332874
rect 116136 332846 116334 332874
rect 96724 332302 97014 332330
rect 95146 323232 95202 323241
rect 95146 323167 95202 323176
rect 91098 322552 91154 322561
rect 91098 322487 91154 322496
rect 90456 314628 90508 314634
rect 90456 314570 90508 314576
rect 91112 314566 91140 322487
rect 95160 314634 95188 323167
rect 95148 314628 95200 314634
rect 95148 314570 95200 314576
rect 91100 314560 91152 314566
rect 91100 314502 91152 314508
rect 96724 311846 96752 332302
rect 96816 313126 97014 313154
rect 106568 313126 106674 313154
rect 116228 313126 116334 313154
rect 96712 311840 96764 311846
rect 96712 311782 96764 311788
rect 96816 311778 96844 313126
rect 96804 311772 96856 311778
rect 96804 311714 96856 311720
rect 106568 311710 106596 313126
rect 116228 313018 116256 313126
rect 116504 313018 116532 335446
rect 116584 335436 116636 335442
rect 116584 335378 116636 335384
rect 116228 312990 116532 313018
rect 116596 311710 116624 335378
rect 133432 332874 133460 335446
rect 142988 335436 143040 335442
rect 142988 335378 143040 335384
rect 144276 335436 144328 335442
rect 144276 335378 144328 335384
rect 143000 332874 143028 335378
rect 144184 335368 144236 335374
rect 144184 335310 144236 335316
rect 133432 332846 133722 332874
rect 143000 332846 143382 332874
rect 122944 332302 124062 332330
rect 122746 323232 122802 323241
rect 122746 323167 122802 323176
rect 118698 322552 118754 322561
rect 118698 322487 118754 322496
rect 118712 314498 118740 322487
rect 122760 314566 122788 323167
rect 122748 314560 122800 314566
rect 122748 314502 122800 314508
rect 118700 314492 118752 314498
rect 118700 314434 118752 314440
rect 79968 311704 80020 311710
rect 79968 311646 80020 311652
rect 90364 311704 90416 311710
rect 90364 311646 90416 311652
rect 106556 311704 106608 311710
rect 106556 311646 106608 311652
rect 116584 311704 116636 311710
rect 116584 311646 116636 311652
rect 122944 311642 122972 332302
rect 144196 316034 144224 335310
rect 143736 316006 144224 316034
rect 143736 313698 143764 316006
rect 143382 313670 143764 313698
rect 123680 313126 124062 313154
rect 133722 313126 133828 313154
rect 123680 311778 123708 313126
rect 123668 311772 123720 311778
rect 123668 311714 123720 311720
rect 133800 311710 133828 313126
rect 144288 311710 144316 335378
rect 146298 322008 146354 322017
rect 146298 321943 146354 321952
rect 146312 314634 146340 321943
rect 146300 314628 146352 314634
rect 146300 314570 146352 314576
rect 133788 311704 133840 311710
rect 133788 311646 133840 311652
rect 144276 311704 144328 311710
rect 144276 311646 144328 311652
rect 122932 311636 122984 311642
rect 122932 311578 122984 311584
rect 52644 308032 52696 308038
rect 52644 307974 52696 307980
rect 43076 307828 43128 307834
rect 43076 307770 43128 307776
rect 43088 305932 43116 307770
rect 52656 305932 52684 307974
rect 62488 307964 62540 307970
rect 62488 307906 62540 307912
rect 79692 307964 79744 307970
rect 79692 307906 79744 307912
rect 90364 307964 90416 307970
rect 90364 307906 90416 307912
rect 106648 307964 106700 307970
rect 106648 307906 106700 307912
rect 116492 307964 116544 307970
rect 116492 307906 116544 307912
rect 133696 307964 133748 307970
rect 133696 307906 133748 307912
rect 144184 307964 144236 307970
rect 144184 307906 144236 307912
rect 62304 307896 62356 307902
rect 62304 307838 62356 307844
rect 62316 305932 62344 307838
rect 37924 305652 37976 305658
rect 37924 305594 37976 305600
rect 41326 296304 41382 296313
rect 41326 296239 41382 296248
rect 37922 295352 37978 295361
rect 37922 295287 37978 295296
rect 36820 286952 36872 286958
rect 36820 286894 36872 286900
rect 36728 284164 36780 284170
rect 36728 284106 36780 284112
rect 36636 284028 36688 284034
rect 36636 283970 36688 283976
rect 36820 280424 36872 280430
rect 36820 280366 36872 280372
rect 36728 280288 36780 280294
rect 36728 280230 36780 280236
rect 36636 277500 36688 277506
rect 36636 277442 36688 277448
rect 36544 256420 36596 256426
rect 36544 256362 36596 256368
rect 16304 254584 16356 254590
rect 16304 254526 16356 254532
rect 25688 254244 25740 254250
rect 25688 254186 25740 254192
rect 25700 251940 25728 254186
rect 15212 251246 16054 251274
rect 35374 251246 36032 251274
rect 13726 242176 13782 242185
rect 13726 242111 13782 242120
rect 13740 233238 13768 242111
rect 13728 233232 13780 233238
rect 13728 233174 13780 233180
rect 15212 230382 15240 251246
rect 36004 248414 36032 251246
rect 36004 248386 36584 248414
rect 35374 232762 35664 232778
rect 35374 232756 35676 232762
rect 35374 232750 35624 232756
rect 35624 232698 35676 232704
rect 15304 232070 16054 232098
rect 25714 232070 26096 232098
rect 15200 230376 15252 230382
rect 15200 230318 15252 230324
rect 15304 227050 15332 232070
rect 26068 230450 26096 232070
rect 26056 230444 26108 230450
rect 26056 230386 26108 230392
rect 15292 227044 15344 227050
rect 15292 226986 15344 226992
rect 25964 226636 26016 226642
rect 25964 226578 26016 226584
rect 25976 224890 26004 226578
rect 25714 224862 26004 224890
rect 15212 224318 16054 224346
rect 35374 224318 35664 224346
rect 13726 215248 13782 215257
rect 13726 215183 13782 215192
rect 13740 205630 13768 215183
rect 13728 205624 13780 205630
rect 13728 205566 13780 205572
rect 15212 202774 15240 224318
rect 35636 223650 35664 224318
rect 35624 223644 35676 223650
rect 35624 223586 35676 223592
rect 35374 205562 35664 205578
rect 35374 205556 35676 205562
rect 35374 205550 35624 205556
rect 35624 205498 35676 205504
rect 15200 202768 15252 202774
rect 15200 202710 15252 202716
rect 16040 200802 16068 205020
rect 25700 202706 25728 205020
rect 25688 202700 25740 202706
rect 25688 202642 25740 202648
rect 36556 202570 36584 248386
rect 36648 230178 36676 277442
rect 36740 256698 36768 280230
rect 36832 259418 36860 280366
rect 37936 279478 37964 295287
rect 41340 286958 41368 296239
rect 41328 286952 41380 286958
rect 41328 286894 41380 286900
rect 62500 286770 62528 307906
rect 64144 307896 64196 307902
rect 64144 307838 64196 307844
rect 62764 307828 62816 307834
rect 62764 307770 62816 307776
rect 62422 286742 62528 286770
rect 42996 284238 43024 286076
rect 52748 284238 52776 286076
rect 62776 284306 62804 307770
rect 62764 284300 62816 284306
rect 62764 284242 62816 284248
rect 64156 284238 64184 307838
rect 79704 305932 79732 307906
rect 89352 307896 89404 307902
rect 89352 307838 89404 307844
rect 89364 305932 89392 307838
rect 69124 305238 70058 305266
rect 68926 295760 68982 295769
rect 68926 295695 68982 295704
rect 64878 295624 64934 295633
rect 64878 295559 64934 295568
rect 64892 287026 64920 295559
rect 64880 287020 64932 287026
rect 64880 286962 64932 286968
rect 68940 286890 68968 295695
rect 68928 286884 68980 286890
rect 68928 286826 68980 286832
rect 69124 284238 69152 305238
rect 90376 287054 90404 307906
rect 90456 307896 90508 307902
rect 90456 307838 90508 307844
rect 89824 287026 90404 287054
rect 89824 286770 89852 287026
rect 89378 286742 89852 286770
rect 70044 284306 70072 286076
rect 70032 284300 70084 284306
rect 70032 284242 70084 284248
rect 42984 284232 43036 284238
rect 42984 284174 43036 284180
rect 52736 284232 52788 284238
rect 52736 284174 52788 284180
rect 64144 284232 64196 284238
rect 64144 284174 64196 284180
rect 69112 284232 69164 284238
rect 69112 284174 69164 284180
rect 79704 284170 79732 286076
rect 90468 284170 90496 307838
rect 106660 305932 106688 307906
rect 116308 307896 116360 307902
rect 116308 307838 116360 307844
rect 116320 305932 116348 307838
rect 96724 305238 97014 305266
rect 95146 296304 95202 296313
rect 95146 296239 95202 296248
rect 91098 295624 91154 295633
rect 91098 295559 91154 295568
rect 91112 286958 91140 295559
rect 95160 287026 95188 296239
rect 95148 287020 95200 287026
rect 95148 286962 95200 286968
rect 91100 286952 91152 286958
rect 91100 286894 91152 286900
rect 96724 284306 96752 305238
rect 96712 284300 96764 284306
rect 96712 284242 96764 284248
rect 97000 284238 97028 286076
rect 96988 284232 97040 284238
rect 96988 284174 97040 284180
rect 106660 284170 106688 286076
rect 116320 285954 116348 286076
rect 116504 285954 116532 307906
rect 116584 307896 116636 307902
rect 116584 307838 116636 307844
rect 116320 285926 116532 285954
rect 116596 284170 116624 307838
rect 133708 305932 133736 307906
rect 143356 307896 143408 307902
rect 143356 307838 143408 307844
rect 143368 305932 143396 307838
rect 122944 305238 124062 305266
rect 122746 296304 122802 296313
rect 122746 296239 122802 296248
rect 118698 295624 118754 295633
rect 118698 295559 118754 295568
rect 118712 286890 118740 295559
rect 122760 286958 122788 296239
rect 122748 286952 122800 286958
rect 122748 286894 122800 286900
rect 118700 286884 118752 286890
rect 118700 286826 118752 286832
rect 122944 284170 122972 305238
rect 144196 287054 144224 307906
rect 144276 307896 144328 307902
rect 144276 307838 144328 307844
rect 143736 287026 144224 287054
rect 143736 286770 143764 287026
rect 143382 286742 143764 286770
rect 124048 284238 124076 286076
rect 133708 284238 133736 286076
rect 144288 284238 144316 307838
rect 146298 295352 146354 295361
rect 146298 295287 146354 295296
rect 146312 287026 146340 295287
rect 146300 287020 146352 287026
rect 146300 286962 146352 286968
rect 146956 284306 146984 335582
rect 148966 323232 149022 323241
rect 148966 323167 149022 323176
rect 148980 314634 149008 323167
rect 148968 314628 149020 314634
rect 148968 314570 149020 314576
rect 149716 311778 149744 361830
rect 232044 361820 232096 361826
rect 232044 361762 232096 361768
rect 251824 361820 251876 361826
rect 251824 361762 251876 361768
rect 475016 361820 475068 361826
rect 475016 361762 475068 361768
rect 494704 361820 494756 361826
rect 494704 361762 494756 361768
rect 160652 361752 160704 361758
rect 160652 361694 160704 361700
rect 170496 361752 170548 361758
rect 170496 361694 170548 361700
rect 187700 361752 187752 361758
rect 187700 361694 187752 361700
rect 197452 361752 197504 361758
rect 197452 361694 197504 361700
rect 214656 361752 214708 361758
rect 214656 361694 214708 361700
rect 224500 361752 224552 361758
rect 224500 361694 224552 361700
rect 160664 359924 160692 361694
rect 170312 361684 170364 361690
rect 170312 361626 170364 361632
rect 170324 359924 170352 361626
rect 150544 359230 151018 359258
rect 150544 338026 150572 359230
rect 150532 338020 150584 338026
rect 150532 337962 150584 337968
rect 151004 337958 151032 340068
rect 150992 337952 151044 337958
rect 150992 337894 151044 337900
rect 160664 337890 160692 340068
rect 170324 339946 170352 340068
rect 170508 339946 170536 361694
rect 178040 361684 178092 361690
rect 178040 361626 178092 361632
rect 171784 361616 171836 361622
rect 171784 361558 171836 361564
rect 170324 339918 170536 339946
rect 171796 337890 171824 361558
rect 178052 359924 178080 361626
rect 187712 359924 187740 361694
rect 197360 361616 197412 361622
rect 197360 361558 197412 361564
rect 197372 359924 197400 361558
rect 176566 349752 176622 349761
rect 176566 349687 176622 349696
rect 172518 349616 172574 349625
rect 172518 349551 172574 349560
rect 172532 340814 172560 349551
rect 176580 340814 176608 349687
rect 172520 340808 172572 340814
rect 172520 340750 172572 340756
rect 176568 340808 176620 340814
rect 197464 340762 197492 361694
rect 200764 361684 200816 361690
rect 200764 361626 200816 361632
rect 199384 361616 199436 361622
rect 199384 361558 199436 361564
rect 176568 340750 176620 340756
rect 197386 340734 197492 340762
rect 178052 337958 178080 340068
rect 187712 337958 187740 340068
rect 199396 337958 199424 361558
rect 200118 349616 200174 349625
rect 200118 349551 200174 349560
rect 200132 340882 200160 349551
rect 200120 340876 200172 340882
rect 200120 340818 200172 340824
rect 200776 340746 200804 361626
rect 214668 359924 214696 361694
rect 224316 361616 224368 361622
rect 224316 361558 224368 361564
rect 224328 359924 224356 361558
rect 204364 359230 205022 359258
rect 202786 350296 202842 350305
rect 202786 350231 202842 350240
rect 202800 340882 202828 350231
rect 202788 340876 202840 340882
rect 202788 340818 202840 340824
rect 200764 340740 200816 340746
rect 200764 340682 200816 340688
rect 204364 337958 204392 359230
rect 224512 340762 224540 361694
rect 225604 361616 225656 361622
rect 225604 361558 225656 361564
rect 204640 340746 205022 340762
rect 204628 340740 205022 340746
rect 204680 340734 205022 340740
rect 224342 340734 224540 340762
rect 204628 340682 204680 340688
rect 178040 337952 178092 337958
rect 178040 337894 178092 337900
rect 187700 337952 187752 337958
rect 187700 337894 187752 337900
rect 199384 337952 199436 337958
rect 199384 337894 199436 337900
rect 204352 337952 204404 337958
rect 204352 337894 204404 337900
rect 214668 337890 214696 340068
rect 225616 337890 225644 361558
rect 232056 359924 232084 361762
rect 241704 361752 241756 361758
rect 241704 361694 241756 361700
rect 241716 359924 241744 361694
rect 251456 361684 251508 361690
rect 251456 361626 251508 361632
rect 251364 361616 251416 361622
rect 251364 361558 251416 361564
rect 251376 359924 251404 361558
rect 230386 350296 230442 350305
rect 230386 350231 230442 350240
rect 226338 349616 226394 349625
rect 226338 349551 226394 349560
rect 226352 340814 226380 349551
rect 230400 340814 230428 350231
rect 226340 340808 226392 340814
rect 226340 340750 226392 340756
rect 230388 340808 230440 340814
rect 251468 340762 251496 361626
rect 230388 340750 230440 340756
rect 251390 340734 251496 340762
rect 232056 337958 232084 340068
rect 241716 337958 241744 340068
rect 251836 338094 251864 361762
rect 413468 361752 413520 361758
rect 413468 361694 413520 361700
rect 430672 361752 430724 361758
rect 430672 361694 430724 361700
rect 440516 361752 440568 361758
rect 440516 361694 440568 361700
rect 457628 361752 457680 361758
rect 457628 361694 457680 361700
rect 468576 361752 468628 361758
rect 468576 361694 468628 361700
rect 268660 361684 268712 361690
rect 268660 361626 268712 361632
rect 279516 361684 279568 361690
rect 279516 361626 279568 361632
rect 295708 361684 295760 361690
rect 295708 361626 295760 361632
rect 305460 361684 305512 361690
rect 305460 361626 305512 361632
rect 322664 361684 322716 361690
rect 322664 361626 322716 361632
rect 334624 361684 334676 361690
rect 334624 361626 334676 361632
rect 349712 361684 349764 361690
rect 349712 361626 349764 361632
rect 359464 361684 359516 361690
rect 359464 361626 359516 361632
rect 376668 361684 376720 361690
rect 376668 361626 376720 361632
rect 386512 361684 386564 361690
rect 386512 361626 386564 361632
rect 403624 361684 403676 361690
rect 403624 361626 403676 361632
rect 253204 361616 253256 361622
rect 253204 361558 253256 361564
rect 251824 338088 251876 338094
rect 251824 338030 251876 338036
rect 253216 337958 253244 361558
rect 268672 359924 268700 361626
rect 278320 361616 278372 361622
rect 278320 361558 278372 361564
rect 279424 361616 279476 361622
rect 279424 361558 279476 361564
rect 278332 359924 278360 361558
rect 258184 359230 259026 359258
rect 256606 350296 256662 350305
rect 256606 350231 256662 350240
rect 253938 349208 253994 349217
rect 253938 349143 253994 349152
rect 253952 340882 253980 349143
rect 256620 340882 256648 350231
rect 253940 340876 253992 340882
rect 253940 340818 253992 340824
rect 256608 340876 256660 340882
rect 256608 340818 256660 340824
rect 258184 337958 258212 359230
rect 278346 340746 278728 340762
rect 278346 340740 278740 340746
rect 278346 340734 278688 340740
rect 278688 340682 278740 340688
rect 259012 338094 259040 340068
rect 259000 338088 259052 338094
rect 259000 338030 259052 338036
rect 232044 337952 232096 337958
rect 232044 337894 232096 337900
rect 241704 337952 241756 337958
rect 241704 337894 241756 337900
rect 253204 337952 253256 337958
rect 253204 337894 253256 337900
rect 258172 337952 258224 337958
rect 258172 337894 258224 337900
rect 268672 337890 268700 340068
rect 279436 337890 279464 361558
rect 279528 340746 279556 361626
rect 285784 360046 286088 360074
rect 284206 349752 284262 349761
rect 284206 349687 284262 349696
rect 280158 349616 280214 349625
rect 280158 349551 280214 349560
rect 280172 340814 280200 349551
rect 284220 340814 284248 349687
rect 280160 340808 280212 340814
rect 280160 340750 280212 340756
rect 284208 340808 284260 340814
rect 284208 340750 284260 340756
rect 279516 340740 279568 340746
rect 279516 340682 279568 340688
rect 285784 337890 285812 360046
rect 286060 359924 286088 360046
rect 295720 359924 295748 361626
rect 305368 361616 305420 361622
rect 305368 361558 305420 361564
rect 305380 359924 305408 361558
rect 305472 340762 305500 361626
rect 307024 361616 307076 361622
rect 307024 361558 307076 361564
rect 305394 340734 305500 340762
rect 286060 337958 286088 340068
rect 286048 337952 286100 337958
rect 286048 337894 286100 337900
rect 295720 337890 295748 340068
rect 307036 337890 307064 361558
rect 322676 359924 322704 361626
rect 332324 361616 332376 361622
rect 332324 361558 332376 361564
rect 333244 361616 333296 361622
rect 333244 361558 333296 361564
rect 332336 359924 332364 361558
rect 312004 359230 313030 359258
rect 311806 350296 311862 350305
rect 311806 350231 311862 350240
rect 307758 349616 307814 349625
rect 307758 349551 307814 349560
rect 307772 340882 307800 349551
rect 307760 340876 307812 340882
rect 307760 340818 307812 340824
rect 311820 340746 311848 350231
rect 311808 340740 311860 340746
rect 311808 340682 311860 340688
rect 312004 337890 312032 359230
rect 332508 340876 332560 340882
rect 332508 340818 332560 340824
rect 332520 340762 332548 340818
rect 332350 340734 332548 340762
rect 313016 337958 313044 340068
rect 313004 337952 313056 337958
rect 313004 337894 313056 337900
rect 322676 337890 322704 340068
rect 333256 337890 333284 361558
rect 334636 340882 334664 361626
rect 339604 360046 340092 360074
rect 338026 350296 338082 350305
rect 338026 350231 338082 350240
rect 335358 349616 335414 349625
rect 335358 349551 335414 349560
rect 334624 340876 334676 340882
rect 334624 340818 334676 340824
rect 335372 340814 335400 349551
rect 338040 340882 338068 350231
rect 338028 340876 338080 340882
rect 338028 340818 338080 340824
rect 335360 340808 335412 340814
rect 335360 340750 335412 340756
rect 339604 337890 339632 360046
rect 340064 359924 340092 360046
rect 349724 359924 349752 361626
rect 359372 361616 359424 361622
rect 359372 361558 359424 361564
rect 359384 359924 359412 361558
rect 359476 340762 359504 361626
rect 359556 361616 359608 361622
rect 359556 361558 359608 361564
rect 359398 340734 359504 340762
rect 340064 337958 340092 340068
rect 340052 337952 340104 337958
rect 340052 337894 340104 337900
rect 349724 337890 349752 340068
rect 359568 337890 359596 361558
rect 376680 359924 376708 361626
rect 386328 361616 386380 361622
rect 386328 361558 386380 361564
rect 386340 359924 386368 361558
rect 365824 359230 367034 359258
rect 365626 350296 365682 350305
rect 365626 350231 365682 350240
rect 361578 349208 361634 349217
rect 361578 349143 361634 349152
rect 361592 340746 361620 349143
rect 365640 340814 365668 350231
rect 365628 340808 365680 340814
rect 365628 340750 365680 340756
rect 361580 340740 361632 340746
rect 361580 340682 361632 340688
rect 365824 337890 365852 359230
rect 386524 340762 386552 361626
rect 387064 361616 387116 361622
rect 387064 361558 387116 361564
rect 386354 340734 386552 340762
rect 367020 337958 367048 340068
rect 367008 337952 367060 337958
rect 367008 337894 367060 337900
rect 376680 337890 376708 340068
rect 387076 337890 387104 361558
rect 403636 359924 403664 361626
rect 413284 361616 413336 361622
rect 413284 361558 413336 361564
rect 413296 359924 413324 361558
rect 393424 359230 393990 359258
rect 391846 350296 391902 350305
rect 391846 350231 391902 350240
rect 389178 349616 389234 349625
rect 389178 349551 389234 349560
rect 389192 340882 389220 349551
rect 391860 340882 391888 350231
rect 389180 340876 389232 340882
rect 389180 340818 389232 340824
rect 391848 340876 391900 340882
rect 391848 340818 391900 340824
rect 393424 337890 393452 359230
rect 413480 340762 413508 361694
rect 421012 361684 421064 361690
rect 421012 361626 421064 361632
rect 414664 361616 414716 361622
rect 414664 361558 414716 361564
rect 413402 340734 413508 340762
rect 393976 337958 394004 340068
rect 393964 337952 394016 337958
rect 393964 337894 394016 337900
rect 403728 337890 403756 340068
rect 414676 337890 414704 361558
rect 421024 359924 421052 361626
rect 430684 359924 430712 361694
rect 440332 361616 440384 361622
rect 440332 361558 440384 361564
rect 440344 359924 440372 361558
rect 419446 350296 419502 350305
rect 419446 350231 419502 350240
rect 415398 349616 415454 349625
rect 415398 349551 415454 349560
rect 415412 340814 415440 349551
rect 419460 340814 419488 350231
rect 415400 340808 415452 340814
rect 415400 340750 415452 340756
rect 419448 340808 419500 340814
rect 440528 340762 440556 361694
rect 443644 361684 443696 361690
rect 443644 361626 443696 361632
rect 442264 361616 442316 361622
rect 442264 361558 442316 361564
rect 419448 340750 419500 340756
rect 440358 340734 440556 340762
rect 421024 337958 421052 340068
rect 430684 337958 430712 340068
rect 442276 337958 442304 361558
rect 442998 349616 443054 349625
rect 442998 349551 443054 349560
rect 443012 340882 443040 349551
rect 443656 340950 443684 361626
rect 457640 359924 457668 361694
rect 467288 361616 467340 361622
rect 467288 361558 467340 361564
rect 468484 361616 468536 361622
rect 468484 361558 468536 361564
rect 467300 359924 467328 361558
rect 447244 359230 447994 359258
rect 445666 350296 445722 350305
rect 445666 350231 445722 350240
rect 443644 340944 443696 340950
rect 443644 340886 443696 340892
rect 445680 340882 445708 350231
rect 443000 340876 443052 340882
rect 443000 340818 443052 340824
rect 445668 340876 445720 340882
rect 445668 340818 445720 340824
rect 447244 337958 447272 359230
rect 447692 340944 447744 340950
rect 447692 340886 447744 340892
rect 447704 340762 447732 340886
rect 447704 340734 447994 340762
rect 467406 340746 467696 340762
rect 467406 340740 467708 340746
rect 467406 340734 467656 340740
rect 467656 340682 467708 340688
rect 421012 337952 421064 337958
rect 421012 337894 421064 337900
rect 430672 337952 430724 337958
rect 430672 337894 430724 337900
rect 442264 337952 442316 337958
rect 442264 337894 442316 337900
rect 447232 337952 447284 337958
rect 447232 337894 447284 337900
rect 457732 337890 457760 340068
rect 468496 337890 468524 361558
rect 468588 340746 468616 361694
rect 475028 359924 475056 361762
rect 484676 361752 484728 361758
rect 484676 361694 484728 361700
rect 484688 359924 484716 361694
rect 494520 361684 494572 361690
rect 494520 361626 494572 361632
rect 494336 361616 494388 361622
rect 494336 361558 494388 361564
rect 494348 359924 494376 361558
rect 473266 349752 473322 349761
rect 473266 349687 473322 349696
rect 469218 349208 469274 349217
rect 469218 349143 469274 349152
rect 469232 340814 469260 349143
rect 473280 340814 473308 349687
rect 469220 340808 469272 340814
rect 469220 340750 469272 340756
rect 473268 340808 473320 340814
rect 494532 340762 494560 361626
rect 473268 340750 473320 340756
rect 468576 340740 468628 340746
rect 494362 340734 494560 340762
rect 468576 340682 468628 340688
rect 475028 337958 475056 340068
rect 484688 337958 484716 340068
rect 494716 338094 494744 361762
rect 511632 361684 511684 361690
rect 511632 361626 511684 361632
rect 522304 361684 522356 361690
rect 522304 361626 522356 361632
rect 496084 361616 496136 361622
rect 496084 361558 496136 361564
rect 494704 338088 494756 338094
rect 494704 338030 494756 338036
rect 496096 337958 496124 361558
rect 511644 359924 511672 361626
rect 521292 361616 521344 361622
rect 521292 361558 521344 361564
rect 521304 359924 521332 361558
rect 501064 359230 501998 359258
rect 500866 350296 500922 350305
rect 500866 350231 500922 350240
rect 496818 349616 496874 349625
rect 496818 349551 496874 349560
rect 496832 340882 496860 349551
rect 500880 340882 500908 350231
rect 496820 340876 496872 340882
rect 496820 340818 496872 340824
rect 500868 340876 500920 340882
rect 500868 340818 500920 340824
rect 501064 337958 501092 359230
rect 522316 345014 522344 361626
rect 522396 361616 522448 361622
rect 522396 361558 522448 361564
rect 521856 344986 522344 345014
rect 521856 340762 521884 344986
rect 521410 340734 521884 340762
rect 501984 338094 502012 340068
rect 501972 338088 502024 338094
rect 501972 338030 502024 338036
rect 475016 337952 475068 337958
rect 475016 337894 475068 337900
rect 484676 337952 484728 337958
rect 484676 337894 484728 337900
rect 496084 337952 496136 337958
rect 496084 337894 496136 337900
rect 501052 337952 501104 337958
rect 501052 337894 501104 337900
rect 511736 337890 511764 340068
rect 522408 337890 522436 361558
rect 529032 359924 529060 362170
rect 538680 361684 538732 361690
rect 538680 361626 538732 361632
rect 538692 359924 538720 361626
rect 548340 361616 548392 361622
rect 548340 361558 548392 361564
rect 548352 359924 548380 361558
rect 526444 359508 526496 359514
rect 526444 359450 526496 359456
rect 526456 350305 526484 359450
rect 526442 350296 526498 350305
rect 526442 350231 526498 350240
rect 523038 349616 523094 349625
rect 523038 349551 523094 349560
rect 550638 349616 550694 349625
rect 550638 349551 550694 349560
rect 523052 340814 523080 349551
rect 550652 340882 550680 349551
rect 550640 340876 550692 340882
rect 550640 340818 550692 340824
rect 523040 340808 523092 340814
rect 523040 340750 523092 340756
rect 529032 337958 529060 340068
rect 529020 337952 529072 337958
rect 529020 337894 529072 337900
rect 160652 337884 160704 337890
rect 160652 337826 160704 337832
rect 171784 337884 171836 337890
rect 171784 337826 171836 337832
rect 214656 337884 214708 337890
rect 214656 337826 214708 337832
rect 225604 337884 225656 337890
rect 225604 337826 225656 337832
rect 268660 337884 268712 337890
rect 268660 337826 268712 337832
rect 279424 337884 279476 337890
rect 279424 337826 279476 337832
rect 285772 337884 285824 337890
rect 285772 337826 285824 337832
rect 295708 337884 295760 337890
rect 295708 337826 295760 337832
rect 307024 337884 307076 337890
rect 307024 337826 307076 337832
rect 311992 337884 312044 337890
rect 311992 337826 312044 337832
rect 322664 337884 322716 337890
rect 322664 337826 322716 337832
rect 333244 337884 333296 337890
rect 333244 337826 333296 337832
rect 339592 337884 339644 337890
rect 339592 337826 339644 337832
rect 349712 337884 349764 337890
rect 349712 337826 349764 337832
rect 359556 337884 359608 337890
rect 359556 337826 359608 337832
rect 365812 337884 365864 337890
rect 365812 337826 365864 337832
rect 376668 337884 376720 337890
rect 376668 337826 376720 337832
rect 387064 337884 387116 337890
rect 387064 337826 387116 337832
rect 393412 337884 393464 337890
rect 393412 337826 393464 337832
rect 403716 337884 403768 337890
rect 403716 337826 403768 337832
rect 414664 337884 414716 337890
rect 414664 337826 414716 337832
rect 457720 337884 457772 337890
rect 457720 337826 457772 337832
rect 468484 337884 468536 337890
rect 468484 337826 468536 337832
rect 511724 337884 511776 337890
rect 511724 337826 511776 337832
rect 522396 337884 522448 337890
rect 522396 337826 522448 337832
rect 538692 337822 538720 340068
rect 548352 338026 548380 340068
rect 548340 338020 548392 338026
rect 548340 337962 548392 337968
rect 538680 337816 538732 337822
rect 538680 337758 538732 337764
rect 528652 336048 528704 336054
rect 528652 335990 528704 335996
rect 232320 335572 232372 335578
rect 232320 335514 232372 335520
rect 251824 335572 251876 335578
rect 251824 335514 251876 335520
rect 475384 335572 475436 335578
rect 475384 335514 475436 335520
rect 494704 335572 494756 335578
rect 494704 335514 494756 335520
rect 170496 335504 170548 335510
rect 170496 335446 170548 335452
rect 187792 335504 187844 335510
rect 187792 335446 187844 335452
rect 197544 335504 197596 335510
rect 197544 335446 197596 335452
rect 214380 335504 214432 335510
rect 214380 335446 214432 335452
rect 224500 335504 224552 335510
rect 224500 335446 224552 335452
rect 170036 335436 170088 335442
rect 170036 335378 170088 335384
rect 160284 335368 160336 335374
rect 160284 335310 160336 335316
rect 160296 332874 160324 335310
rect 170048 332874 170076 335378
rect 160296 332846 160678 332874
rect 170048 332846 170338 332874
rect 150544 332302 151018 332330
rect 149704 311772 149756 311778
rect 149704 311714 149756 311720
rect 150544 311710 150572 332302
rect 170232 313682 170338 313698
rect 170508 313682 170536 335446
rect 178408 335436 178460 335442
rect 178408 335378 178460 335384
rect 171784 335368 171836 335374
rect 171784 335310 171836 335316
rect 170220 313676 170338 313682
rect 170272 313670 170338 313676
rect 170496 313676 170548 313682
rect 170220 313618 170272 313624
rect 170496 313618 170548 313624
rect 150728 313126 151018 313154
rect 160572 313126 160678 313154
rect 150532 311704 150584 311710
rect 150532 311646 150584 311652
rect 150728 311642 150756 313126
rect 160572 311642 160600 313126
rect 171796 311642 171824 335310
rect 178420 332874 178448 335378
rect 187804 332874 187832 335446
rect 197452 335368 197504 335374
rect 197452 335310 197504 335316
rect 197464 332874 197492 335310
rect 178066 332846 178448 332874
rect 187726 332846 187832 332874
rect 197386 332846 197492 332874
rect 176566 322960 176622 322969
rect 176566 322895 176622 322904
rect 172518 322552 172574 322561
rect 172518 322487 172574 322496
rect 172532 314566 172560 322487
rect 176580 314566 176608 322895
rect 197556 316034 197584 335446
rect 200764 335436 200816 335442
rect 200764 335378 200816 335384
rect 199384 335368 199436 335374
rect 199384 335310 199436 335316
rect 197464 316006 197584 316034
rect 172520 314560 172572 314566
rect 172520 314502 172572 314508
rect 176568 314560 176620 314566
rect 176568 314502 176620 314508
rect 197464 313698 197492 316006
rect 197386 313670 197492 313698
rect 178066 313126 178172 313154
rect 187726 313126 188016 313154
rect 178144 311710 178172 313126
rect 187988 311710 188016 313126
rect 199396 311710 199424 335310
rect 200118 322552 200174 322561
rect 200118 322487 200174 322496
rect 200132 314634 200160 322487
rect 200120 314628 200172 314634
rect 200120 314570 200172 314576
rect 200776 311846 200804 335378
rect 214392 332874 214420 335446
rect 223948 335368 224000 335374
rect 223948 335310 224000 335316
rect 223960 332874 223988 335310
rect 214392 332846 214682 332874
rect 223960 332846 224342 332874
rect 204364 332302 205022 332330
rect 202786 323232 202842 323241
rect 202786 323167 202842 323176
rect 202800 314634 202828 323167
rect 202788 314628 202840 314634
rect 202788 314570 202840 314576
rect 200764 311840 200816 311846
rect 200764 311782 200816 311788
rect 204364 311710 204392 332302
rect 224512 313698 224540 335446
rect 225604 335368 225656 335374
rect 225604 335310 225656 335316
rect 224342 313670 224540 313698
rect 204640 313126 205022 313154
rect 214682 313126 215064 313154
rect 204640 311846 204668 313126
rect 204628 311840 204680 311846
rect 204628 311782 204680 311788
rect 178132 311704 178184 311710
rect 178132 311646 178184 311652
rect 187976 311704 188028 311710
rect 187976 311646 188028 311652
rect 199384 311704 199436 311710
rect 199384 311646 199436 311652
rect 204352 311704 204404 311710
rect 204352 311646 204404 311652
rect 215036 311642 215064 313126
rect 225616 311642 225644 335310
rect 232332 332874 232360 335514
rect 241612 335504 241664 335510
rect 241612 335446 241664 335452
rect 232070 332846 232360 332874
rect 241624 332874 241652 335446
rect 251456 335436 251508 335442
rect 251456 335378 251508 335384
rect 251272 335368 251324 335374
rect 251272 335310 251324 335316
rect 251284 332874 251312 335310
rect 241624 332846 241730 332874
rect 251284 332846 251390 332874
rect 230386 323232 230442 323241
rect 230386 323167 230442 323176
rect 226338 322552 226394 322561
rect 226338 322487 226394 322496
rect 226352 314566 226380 322487
rect 230400 314566 230428 323167
rect 226340 314560 226392 314566
rect 226340 314502 226392 314508
rect 230388 314560 230440 314566
rect 230388 314502 230440 314508
rect 251468 313698 251496 335378
rect 251390 313670 251496 313698
rect 231872 313126 232070 313154
rect 241730 313126 242112 313154
rect 231872 311710 231900 313126
rect 242084 311710 242112 313126
rect 251836 311846 251864 335514
rect 413468 335504 413520 335510
rect 413468 335446 413520 335452
rect 430580 335504 430632 335510
rect 430580 335446 430632 335452
rect 440516 335504 440568 335510
rect 440516 335446 440568 335452
rect 457260 335504 457312 335510
rect 457260 335446 457312 335452
rect 468484 335504 468536 335510
rect 468484 335446 468536 335452
rect 268292 335436 268344 335442
rect 268292 335378 268344 335384
rect 279516 335436 279568 335442
rect 279516 335378 279568 335384
rect 295800 335436 295852 335442
rect 295800 335378 295852 335384
rect 305552 335436 305604 335442
rect 305552 335378 305604 335384
rect 322388 335436 322440 335442
rect 322388 335378 322440 335384
rect 336004 335436 336056 335442
rect 336004 335378 336056 335384
rect 349804 335436 349856 335442
rect 349804 335378 349856 335384
rect 359648 335436 359700 335442
rect 359648 335378 359700 335384
rect 376300 335436 376352 335442
rect 376300 335378 376352 335384
rect 386512 335436 386564 335442
rect 386512 335378 386564 335384
rect 403348 335436 403400 335442
rect 403348 335378 403400 335384
rect 253204 335368 253256 335374
rect 253204 335310 253256 335316
rect 251824 311840 251876 311846
rect 251824 311782 251876 311788
rect 253216 311710 253244 335310
rect 268304 332874 268332 335378
rect 278044 335368 278096 335374
rect 278044 335310 278096 335316
rect 279424 335368 279476 335374
rect 279424 335310 279476 335316
rect 278056 332874 278084 335310
rect 268304 332846 268686 332874
rect 278056 332846 278346 332874
rect 258184 332302 259026 332330
rect 256606 323232 256662 323241
rect 256606 323167 256662 323176
rect 253938 322008 253994 322017
rect 253938 321943 253994 321952
rect 253952 314634 253980 321943
rect 256620 314634 256648 323167
rect 253940 314628 253992 314634
rect 253940 314570 253992 314576
rect 256608 314628 256660 314634
rect 256608 314570 256660 314576
rect 258184 311710 258212 332302
rect 278688 314492 278740 314498
rect 278688 314434 278740 314440
rect 278700 313698 278728 314434
rect 278346 313670 278728 313698
rect 258736 313126 259026 313154
rect 268686 313126 268976 313154
rect 258736 311846 258764 313126
rect 258724 311840 258776 311846
rect 258724 311782 258776 311788
rect 231860 311704 231912 311710
rect 231860 311646 231912 311652
rect 242072 311704 242124 311710
rect 242072 311646 242124 311652
rect 253204 311704 253256 311710
rect 253204 311646 253256 311652
rect 258172 311704 258224 311710
rect 258172 311646 258224 311652
rect 268948 311642 268976 313126
rect 279436 311642 279464 335310
rect 279528 314498 279556 335378
rect 295812 332874 295840 335378
rect 305460 335368 305512 335374
rect 305460 335310 305512 335316
rect 305472 332874 305500 335310
rect 295734 332846 295840 332874
rect 305394 332846 305500 332874
rect 286074 332314 286180 332330
rect 285772 332308 285824 332314
rect 286074 332308 286192 332314
rect 286074 332302 286140 332308
rect 285772 332250 285824 332256
rect 286140 332250 286192 332256
rect 284206 322960 284262 322969
rect 284206 322895 284262 322904
rect 280158 322552 280214 322561
rect 280158 322487 280214 322496
rect 280172 314566 280200 322487
rect 284220 314566 284248 322895
rect 280160 314560 280212 314566
rect 280160 314502 280212 314508
rect 284208 314560 284260 314566
rect 284208 314502 284260 314508
rect 279516 314492 279568 314498
rect 279516 314434 279568 314440
rect 285784 311642 285812 332250
rect 305564 316034 305592 335378
rect 307024 335368 307076 335374
rect 307024 335310 307076 335316
rect 305472 316006 305592 316034
rect 305472 313698 305500 316006
rect 305394 313670 305500 313698
rect 286074 313126 286180 313154
rect 295734 313126 296024 313154
rect 286152 311710 286180 313126
rect 286140 311704 286192 311710
rect 286140 311646 286192 311652
rect 295996 311642 296024 313126
rect 307036 311642 307064 335310
rect 322400 332874 322428 335378
rect 331956 335368 332008 335374
rect 331956 335310 332008 335316
rect 333244 335368 333296 335374
rect 333244 335310 333296 335316
rect 331968 332874 331996 335310
rect 322400 332846 322690 332874
rect 331968 332846 332350 332874
rect 312004 332302 313030 332330
rect 311806 323232 311862 323241
rect 311806 323167 311862 323176
rect 307758 322552 307814 322561
rect 307758 322487 307814 322496
rect 307772 314634 307800 322487
rect 307760 314628 307812 314634
rect 307760 314570 307812 314576
rect 311820 314498 311848 323167
rect 311808 314492 311860 314498
rect 311808 314434 311860 314440
rect 312004 311642 312032 332302
rect 312648 313126 313030 313154
rect 322690 313126 322888 313154
rect 332350 313126 332548 313154
rect 312648 311710 312676 313126
rect 312636 311704 312688 311710
rect 312636 311646 312688 311652
rect 322860 311642 322888 313126
rect 332520 311846 332548 313126
rect 332508 311840 332560 311846
rect 332508 311782 332560 311788
rect 333256 311642 333284 335310
rect 335358 322552 335414 322561
rect 335358 322487 335414 322496
rect 335372 314566 335400 322487
rect 335360 314560 335412 314566
rect 335360 314502 335412 314508
rect 336016 311846 336044 335378
rect 349816 332874 349844 335378
rect 359464 335368 359516 335374
rect 359464 335310 359516 335316
rect 359556 335368 359608 335374
rect 359556 335310 359608 335316
rect 359476 332874 359504 335310
rect 349738 332846 349844 332874
rect 359398 332846 359504 332874
rect 340078 332314 340184 332330
rect 339592 332308 339644 332314
rect 340078 332308 340196 332314
rect 340078 332302 340144 332308
rect 339592 332250 339644 332256
rect 340144 332250 340196 332256
rect 338026 323232 338082 323241
rect 338026 323167 338082 323176
rect 338040 314634 338068 323167
rect 338028 314628 338080 314634
rect 338028 314570 338080 314576
rect 336004 311840 336056 311846
rect 336004 311782 336056 311788
rect 339604 311642 339632 332250
rect 359568 330682 359596 335310
rect 359556 330676 359608 330682
rect 359556 330618 359608 330624
rect 359660 330562 359688 335378
rect 376312 332874 376340 335378
rect 386052 335368 386104 335374
rect 386052 335310 386104 335316
rect 386064 332874 386092 335310
rect 376312 332846 376694 332874
rect 386064 332846 386354 332874
rect 359476 330534 359688 330562
rect 365824 332302 367034 332330
rect 359476 313698 359504 330534
rect 359556 330472 359608 330478
rect 359556 330414 359608 330420
rect 359398 313670 359504 313698
rect 340078 313126 340184 313154
rect 349738 313126 350120 313154
rect 340156 311710 340184 313126
rect 340144 311704 340196 311710
rect 340144 311646 340196 311652
rect 350092 311642 350120 313126
rect 359568 311642 359596 330414
rect 365626 323232 365682 323241
rect 365626 323167 365682 323176
rect 361578 322008 361634 322017
rect 361578 321943 361634 321952
rect 361592 314498 361620 321943
rect 365640 314566 365668 323167
rect 365628 314560 365680 314566
rect 365628 314502 365680 314508
rect 361580 314492 361632 314498
rect 361580 314434 361632 314440
rect 365824 311642 365852 332302
rect 386524 313698 386552 335378
rect 387064 335368 387116 335374
rect 387064 335310 387116 335316
rect 386354 313670 386552 313698
rect 366744 313126 367034 313154
rect 376588 313126 376694 313154
rect 366744 311710 366772 313126
rect 366732 311704 366784 311710
rect 366732 311646 366784 311652
rect 376588 311642 376616 313126
rect 387076 311642 387104 335310
rect 403360 332874 403388 335378
rect 412916 335368 412968 335374
rect 412916 335310 412968 335316
rect 412928 332874 412956 335310
rect 403360 332846 403650 332874
rect 412928 332846 413310 332874
rect 393424 332302 393990 332330
rect 391846 323232 391902 323241
rect 391846 323167 391902 323176
rect 389178 322552 389234 322561
rect 389178 322487 389234 322496
rect 389192 314634 389220 322487
rect 391860 314634 391888 323167
rect 389180 314628 389232 314634
rect 389180 314570 389232 314576
rect 391848 314628 391900 314634
rect 391848 314570 391900 314576
rect 393424 311642 393452 332302
rect 413480 313698 413508 335446
rect 421288 335436 421340 335442
rect 421288 335378 421340 335384
rect 414664 335368 414716 335374
rect 414664 335310 414716 335316
rect 413402 313670 413508 313698
rect 393608 313126 393990 313154
rect 403742 313126 404032 313154
rect 393608 311710 393636 313126
rect 393596 311704 393648 311710
rect 393596 311646 393648 311652
rect 404004 311642 404032 313126
rect 414676 311642 414704 335310
rect 421300 332874 421328 335378
rect 421038 332846 421328 332874
rect 430592 332874 430620 335446
rect 440240 335368 440292 335374
rect 440240 335310 440292 335316
rect 440252 332874 440280 335310
rect 430592 332846 430698 332874
rect 440252 332846 440358 332874
rect 419446 323232 419502 323241
rect 419446 323167 419502 323176
rect 415398 322552 415454 322561
rect 415398 322487 415454 322496
rect 415412 314566 415440 322487
rect 419460 314566 419488 323167
rect 415400 314560 415452 314566
rect 415400 314502 415452 314508
rect 419448 314560 419500 314566
rect 419448 314502 419500 314508
rect 440528 313698 440556 335446
rect 446404 335436 446456 335442
rect 446404 335378 446456 335384
rect 442264 335368 442316 335374
rect 442264 335310 442316 335316
rect 440358 313670 440556 313698
rect 420932 313126 421038 313154
rect 430698 313126 431080 313154
rect 420932 311710 420960 313126
rect 431052 311710 431080 313126
rect 442276 311710 442304 335310
rect 445666 323232 445722 323241
rect 445666 323167 445722 323176
rect 442998 322552 443054 322561
rect 442998 322487 443054 322496
rect 443012 314634 443040 322487
rect 445680 314702 445708 323167
rect 445668 314696 445720 314702
rect 445668 314638 445720 314644
rect 446416 314634 446444 335378
rect 457272 332874 457300 335446
rect 467012 335368 467064 335374
rect 467012 335310 467064 335316
rect 467024 332874 467052 335310
rect 457272 332846 457654 332874
rect 467024 332846 467314 332874
rect 447244 332302 447994 332330
rect 443000 314628 443052 314634
rect 443000 314570 443052 314576
rect 446404 314628 446456 314634
rect 446404 314570 446456 314576
rect 447244 311710 447272 332302
rect 468496 316034 468524 335446
rect 468576 335368 468628 335374
rect 468576 335310 468628 335316
rect 467852 316006 468524 316034
rect 447692 314628 447744 314634
rect 447692 314570 447744 314576
rect 447704 313698 447732 314570
rect 467852 313698 467880 316006
rect 447704 313670 447994 313698
rect 467406 313670 467880 313698
rect 457746 313126 458128 313154
rect 420920 311704 420972 311710
rect 420920 311646 420972 311652
rect 431040 311704 431092 311710
rect 431040 311646 431092 311652
rect 442264 311704 442316 311710
rect 442264 311646 442316 311652
rect 447232 311704 447284 311710
rect 447232 311646 447284 311652
rect 458100 311642 458128 313126
rect 468588 311642 468616 335310
rect 475396 332874 475424 335514
rect 484400 335504 484452 335510
rect 484400 335446 484452 335452
rect 475042 332846 475424 332874
rect 484412 332874 484440 335446
rect 494520 335436 494572 335442
rect 494520 335378 494572 335384
rect 494060 335368 494112 335374
rect 494060 335310 494112 335316
rect 494072 332874 494100 335310
rect 484412 332846 484702 332874
rect 494072 332846 494362 332874
rect 473266 322960 473322 322969
rect 473266 322895 473322 322904
rect 469218 322008 469274 322017
rect 469218 321943 469274 321952
rect 469232 314566 469260 321943
rect 473280 314566 473308 322895
rect 469220 314560 469272 314566
rect 469220 314502 469272 314508
rect 473268 314560 473320 314566
rect 473268 314502 473320 314508
rect 494532 313698 494560 335378
rect 494362 313670 494560 313698
rect 474752 313126 475042 313154
rect 484702 313126 484992 313154
rect 474752 311710 474780 313126
rect 484964 311710 484992 313126
rect 494716 311846 494744 335514
rect 511356 335436 511408 335442
rect 511356 335378 511408 335384
rect 522304 335436 522356 335442
rect 522304 335378 522356 335384
rect 496084 335368 496136 335374
rect 496084 335310 496136 335316
rect 494704 311840 494756 311846
rect 494704 311782 494756 311788
rect 496096 311710 496124 335310
rect 511368 332874 511396 335378
rect 520924 335368 520976 335374
rect 520924 335310 520976 335316
rect 520936 332874 520964 335310
rect 511368 332846 511658 332874
rect 520936 332846 521318 332874
rect 501064 332302 501998 332330
rect 500866 323232 500922 323241
rect 500866 323167 500922 323176
rect 496818 322552 496874 322561
rect 496818 322487 496874 322496
rect 496832 314634 496860 322487
rect 500880 314634 500908 323167
rect 496820 314628 496872 314634
rect 496820 314570 496872 314576
rect 500868 314628 500920 314634
rect 500868 314570 500920 314576
rect 501064 311710 501092 332302
rect 522316 316034 522344 335378
rect 522396 335368 522448 335374
rect 522396 335310 522448 335316
rect 521856 316006 522344 316034
rect 521856 313698 521884 316006
rect 521410 313670 521884 313698
rect 501616 313126 501998 313154
rect 511750 313126 511948 313154
rect 501616 311846 501644 313126
rect 501604 311840 501656 311846
rect 501604 311782 501656 311788
rect 474740 311704 474792 311710
rect 474740 311646 474792 311652
rect 484952 311704 485004 311710
rect 484952 311646 485004 311652
rect 496084 311704 496136 311710
rect 496084 311646 496136 311652
rect 501052 311704 501104 311710
rect 501052 311646 501104 311652
rect 511920 311642 511948 313126
rect 522408 311642 522436 335310
rect 526444 333260 526496 333266
rect 526444 333202 526496 333208
rect 526456 323377 526484 333202
rect 528664 332874 528692 335990
rect 538404 335436 538456 335442
rect 538404 335378 538456 335384
rect 538416 332874 538444 335378
rect 547972 335368 548024 335374
rect 547972 335310 548024 335316
rect 547984 332874 548012 335310
rect 528664 332846 529046 332874
rect 538416 332846 538706 332874
rect 547984 332846 548366 332874
rect 526442 323368 526498 323377
rect 526442 323303 526498 323312
rect 523038 322552 523094 322561
rect 523038 322487 523094 322496
rect 550638 322552 550694 322561
rect 550638 322487 550694 322496
rect 523052 314566 523080 322487
rect 550652 314634 550680 322487
rect 550640 314628 550692 314634
rect 550640 314570 550692 314576
rect 523040 314560 523092 314566
rect 523040 314502 523092 314508
rect 528756 313126 529046 313154
rect 538416 313126 538706 313154
rect 548076 313126 548366 313154
rect 528756 311710 528784 313126
rect 528744 311704 528796 311710
rect 528744 311646 528796 311652
rect 150716 311636 150768 311642
rect 150716 311578 150768 311584
rect 160560 311636 160612 311642
rect 160560 311578 160612 311584
rect 171784 311636 171836 311642
rect 171784 311578 171836 311584
rect 215024 311636 215076 311642
rect 215024 311578 215076 311584
rect 225604 311636 225656 311642
rect 225604 311578 225656 311584
rect 268936 311636 268988 311642
rect 268936 311578 268988 311584
rect 279424 311636 279476 311642
rect 279424 311578 279476 311584
rect 285772 311636 285824 311642
rect 285772 311578 285824 311584
rect 295984 311636 296036 311642
rect 295984 311578 296036 311584
rect 307024 311636 307076 311642
rect 307024 311578 307076 311584
rect 311992 311636 312044 311642
rect 311992 311578 312044 311584
rect 322848 311636 322900 311642
rect 322848 311578 322900 311584
rect 333244 311636 333296 311642
rect 333244 311578 333296 311584
rect 339592 311636 339644 311642
rect 339592 311578 339644 311584
rect 350080 311636 350132 311642
rect 350080 311578 350132 311584
rect 359556 311636 359608 311642
rect 359556 311578 359608 311584
rect 365812 311636 365864 311642
rect 365812 311578 365864 311584
rect 376576 311636 376628 311642
rect 376576 311578 376628 311584
rect 387064 311636 387116 311642
rect 387064 311578 387116 311584
rect 393412 311636 393464 311642
rect 393412 311578 393464 311584
rect 403992 311636 404044 311642
rect 403992 311578 404044 311584
rect 414664 311636 414716 311642
rect 414664 311578 414716 311584
rect 458088 311636 458140 311642
rect 458088 311578 458140 311584
rect 468576 311636 468628 311642
rect 468576 311578 468628 311584
rect 511908 311636 511960 311642
rect 511908 311578 511960 311584
rect 522396 311636 522448 311642
rect 522396 311578 522448 311584
rect 538416 311574 538444 313126
rect 548076 311778 548104 313126
rect 548064 311772 548116 311778
rect 548064 311714 548116 311720
rect 538404 311568 538456 311574
rect 538404 311510 538456 311516
rect 529020 308440 529072 308446
rect 529020 308382 529072 308388
rect 149704 308100 149756 308106
rect 149704 308042 149756 308048
rect 148966 296304 149022 296313
rect 148966 296239 149022 296248
rect 148980 287026 149008 296239
rect 148968 287020 149020 287026
rect 148968 286962 149020 286968
rect 146944 284300 146996 284306
rect 146944 284242 146996 284248
rect 124036 284232 124088 284238
rect 124036 284174 124088 284180
rect 133696 284232 133748 284238
rect 133696 284174 133748 284180
rect 144276 284232 144328 284238
rect 144276 284174 144328 284180
rect 79692 284164 79744 284170
rect 79692 284106 79744 284112
rect 90456 284164 90508 284170
rect 90456 284106 90508 284112
rect 106648 284164 106700 284170
rect 106648 284106 106700 284112
rect 116584 284164 116636 284170
rect 116584 284106 116636 284112
rect 122932 284164 122984 284170
rect 122932 284106 122984 284112
rect 146944 280492 146996 280498
rect 146944 280434 146996 280440
rect 52460 280424 52512 280430
rect 52460 280366 52512 280372
rect 43352 280220 43404 280226
rect 43352 280162 43404 280168
rect 37924 279472 37976 279478
rect 37924 279414 37976 279420
rect 43364 278882 43392 280162
rect 43102 278854 43392 278882
rect 52472 278882 52500 280366
rect 62488 280356 62540 280362
rect 62488 280298 62540 280304
rect 79324 280356 79376 280362
rect 79324 280298 79376 280304
rect 90364 280356 90416 280362
rect 90364 280298 90416 280304
rect 106372 280356 106424 280362
rect 106372 280298 106424 280304
rect 116492 280356 116544 280362
rect 116492 280298 116544 280304
rect 133420 280356 133472 280362
rect 133420 280298 133472 280304
rect 62120 280288 62172 280294
rect 62120 280230 62172 280236
rect 62132 278882 62160 280230
rect 52472 278854 52670 278882
rect 62132 278854 62330 278882
rect 41328 277500 41380 277506
rect 41328 277442 41380 277448
rect 41340 269385 41368 277442
rect 41326 269376 41382 269385
rect 41326 269311 41382 269320
rect 37922 268016 37978 268025
rect 37922 267951 37978 267960
rect 36820 259412 36872 259418
rect 36820 259354 36872 259360
rect 36728 256692 36780 256698
rect 36728 256634 36780 256640
rect 36820 254176 36872 254182
rect 36820 254118 36872 254124
rect 36728 254040 36780 254046
rect 36728 253982 36780 253988
rect 36740 230450 36768 253982
rect 36832 232762 36860 254118
rect 37936 251870 37964 267951
rect 62500 259706 62528 280298
rect 64144 280288 64196 280294
rect 64144 280230 64196 280236
rect 62764 280220 62816 280226
rect 62764 280162 62816 280168
rect 62422 259678 62528 259706
rect 42812 259134 43010 259162
rect 52762 259134 53144 259162
rect 42812 256630 42840 259134
rect 53116 256630 53144 259134
rect 62776 256698 62804 280162
rect 62764 256692 62816 256698
rect 62764 256634 62816 256640
rect 64156 256630 64184 280230
rect 79336 278882 79364 280298
rect 89076 280288 89128 280294
rect 89076 280230 89128 280236
rect 89088 278882 89116 280230
rect 79336 278854 79718 278882
rect 89088 278854 89378 278882
rect 69124 278310 70058 278338
rect 68928 277568 68980 277574
rect 68928 277510 68980 277516
rect 64880 277432 64932 277438
rect 64880 277374 64932 277380
rect 64892 268705 64920 277374
rect 68940 269929 68968 277510
rect 68926 269920 68982 269929
rect 68926 269855 68982 269864
rect 64878 268696 64934 268705
rect 64878 268631 64934 268640
rect 69124 256630 69152 278310
rect 90376 267734 90404 280298
rect 90456 280288 90508 280294
rect 90456 280230 90508 280236
rect 89824 267706 90404 267734
rect 89824 259434 89852 267706
rect 89378 259406 89852 259434
rect 69768 259134 70058 259162
rect 79718 259134 80008 259162
rect 69768 256698 69796 259134
rect 69756 256692 69808 256698
rect 69756 256634 69808 256640
rect 42800 256624 42852 256630
rect 42800 256566 42852 256572
rect 53104 256624 53156 256630
rect 53104 256566 53156 256572
rect 64144 256624 64196 256630
rect 64144 256566 64196 256572
rect 69112 256624 69164 256630
rect 69112 256566 69164 256572
rect 79980 256562 80008 259134
rect 90468 256562 90496 280230
rect 106384 278882 106412 280298
rect 115940 280288 115992 280294
rect 115940 280230 115992 280236
rect 115952 278882 115980 280230
rect 106384 278854 106674 278882
rect 115952 278854 116334 278882
rect 96724 278310 97014 278338
rect 91100 277500 91152 277506
rect 91100 277442 91152 277448
rect 91112 268705 91140 277442
rect 95148 277432 95200 277438
rect 95148 277374 95200 277380
rect 95160 269385 95188 277374
rect 95146 269376 95202 269385
rect 95146 269311 95202 269320
rect 91098 268696 91154 268705
rect 91098 268631 91154 268640
rect 96724 267734 96752 278310
rect 96632 267706 96752 267734
rect 96632 256698 96660 267706
rect 96724 259134 97014 259162
rect 106568 259134 106674 259162
rect 116228 259134 116334 259162
rect 96620 256692 96672 256698
rect 96620 256634 96672 256640
rect 96724 256630 96752 259134
rect 96712 256624 96764 256630
rect 96712 256566 96764 256572
rect 106568 256562 106596 259134
rect 116228 259026 116256 259134
rect 116504 259026 116532 280298
rect 116584 280288 116636 280294
rect 116584 280230 116636 280236
rect 116228 258998 116532 259026
rect 116596 256562 116624 280230
rect 133432 278882 133460 280298
rect 142988 280288 143040 280294
rect 142988 280230 143040 280236
rect 144276 280288 144328 280294
rect 144276 280230 144328 280236
rect 143000 278882 143028 280230
rect 144184 280220 144236 280226
rect 144184 280162 144236 280168
rect 133432 278854 133722 278882
rect 143000 278854 143382 278882
rect 122944 278310 124062 278338
rect 118700 277568 118752 277574
rect 118700 277510 118752 277516
rect 118712 268705 118740 277510
rect 122748 277500 122800 277506
rect 122748 277442 122800 277448
rect 122760 269385 122788 277442
rect 122746 269376 122802 269385
rect 122746 269311 122802 269320
rect 118698 268696 118754 268705
rect 118698 268631 118754 268640
rect 79968 256556 80020 256562
rect 79968 256498 80020 256504
rect 90456 256556 90508 256562
rect 90456 256498 90508 256504
rect 106556 256556 106608 256562
rect 106556 256498 106608 256504
rect 116584 256556 116636 256562
rect 116584 256498 116636 256504
rect 122944 256494 122972 278310
rect 144196 267734 144224 280162
rect 143736 267706 144224 267734
rect 143736 259706 143764 267706
rect 143382 259678 143764 259706
rect 123680 259134 124062 259162
rect 133722 259134 133828 259162
rect 123680 256630 123708 259134
rect 123668 256624 123720 256630
rect 123668 256566 123720 256572
rect 133800 256562 133828 259134
rect 144288 256562 144316 280230
rect 146300 277432 146352 277438
rect 146300 277374 146352 277380
rect 146312 269113 146340 277374
rect 146298 269104 146354 269113
rect 146298 269039 146354 269048
rect 133788 256556 133840 256562
rect 133788 256498 133840 256504
rect 144276 256556 144328 256562
rect 144276 256498 144328 256504
rect 122932 256488 122984 256494
rect 122932 256430 122984 256436
rect 52644 254176 52696 254182
rect 52644 254118 52696 254124
rect 43076 253972 43128 253978
rect 43076 253914 43128 253920
rect 43088 251940 43116 253914
rect 52656 251940 52684 254118
rect 62488 254108 62540 254114
rect 62488 254050 62540 254056
rect 79692 254108 79744 254114
rect 79692 254050 79744 254056
rect 90364 254108 90416 254114
rect 90364 254050 90416 254056
rect 106648 254108 106700 254114
rect 106648 254050 106700 254056
rect 116492 254108 116544 254114
rect 116492 254050 116544 254056
rect 133696 254108 133748 254114
rect 133696 254050 133748 254056
rect 62304 254040 62356 254046
rect 62304 253982 62356 253988
rect 62316 251940 62344 253982
rect 37924 251864 37976 251870
rect 37924 251806 37976 251812
rect 41328 251252 41380 251258
rect 41328 251194 41380 251200
rect 41340 242321 41368 251194
rect 41326 242312 41382 242321
rect 41326 242247 41382 242256
rect 37922 241904 37978 241913
rect 37922 241839 37978 241848
rect 36820 232756 36872 232762
rect 36820 232698 36872 232704
rect 36728 230444 36780 230450
rect 36728 230386 36780 230392
rect 36636 230172 36688 230178
rect 36636 230114 36688 230120
rect 36820 226568 36872 226574
rect 36820 226510 36872 226516
rect 36728 226432 36780 226438
rect 36728 226374 36780 226380
rect 36636 223644 36688 223650
rect 36636 223586 36688 223592
rect 36544 202564 36596 202570
rect 36544 202506 36596 202512
rect 16028 200796 16080 200802
rect 16028 200738 16080 200744
rect 25688 200456 25740 200462
rect 25688 200398 25740 200404
rect 25700 197948 25728 200398
rect 35374 197390 35940 197418
rect 15212 197254 16054 197282
rect 13726 188184 13782 188193
rect 13726 188119 13782 188128
rect 13740 179382 13768 188119
rect 13728 179376 13780 179382
rect 13728 179318 13780 179324
rect 15212 176594 15240 197254
rect 35912 190454 35940 197390
rect 35912 190426 36584 190454
rect 35624 179308 35676 179314
rect 35624 179250 35676 179256
rect 35636 178786 35664 179250
rect 35374 178758 35664 178786
rect 16054 178078 16344 178106
rect 25714 178078 26096 178106
rect 15200 176588 15252 176594
rect 15200 176530 15252 176536
rect 16316 173194 16344 178078
rect 26068 176526 26096 178078
rect 26056 176520 26108 176526
rect 26056 176462 26108 176468
rect 16304 173188 16356 173194
rect 16304 173130 16356 173136
rect 26056 172848 26108 172854
rect 26056 172790 26108 172796
rect 26068 170898 26096 172790
rect 25714 170870 26096 170898
rect 15212 170326 16054 170354
rect 35374 170326 35664 170354
rect 13726 161256 13782 161265
rect 13726 161191 13782 161200
rect 13740 151774 13768 161191
rect 13728 151768 13780 151774
rect 13728 151710 13780 151716
rect 15212 148986 15240 170326
rect 35636 169794 35664 170326
rect 35624 169788 35676 169794
rect 35624 169730 35676 169736
rect 35374 151706 35664 151722
rect 35374 151700 35676 151706
rect 35374 151694 35624 151700
rect 35624 151642 35676 151648
rect 15200 148980 15252 148986
rect 15200 148922 15252 148928
rect 16040 146946 16068 151028
rect 25700 148918 25728 151028
rect 25688 148912 25740 148918
rect 25688 148854 25740 148860
rect 36556 148782 36584 190426
rect 36648 176390 36676 223586
rect 36740 202706 36768 226374
rect 36832 205562 36860 226510
rect 37936 225622 37964 241839
rect 62500 232778 62528 254050
rect 64144 254040 64196 254046
rect 64144 253982 64196 253988
rect 62764 253972 62816 253978
rect 62764 253914 62816 253920
rect 62422 232750 62528 232778
rect 42812 232070 43010 232098
rect 52762 232070 53144 232098
rect 42812 230382 42840 232070
rect 53116 230382 53144 232070
rect 62776 230450 62804 253914
rect 62764 230444 62816 230450
rect 62764 230386 62816 230392
rect 64156 230382 64184 253982
rect 79704 251940 79732 254050
rect 89352 254040 89404 254046
rect 89352 253982 89404 253988
rect 89364 251940 89392 253982
rect 68928 251320 68980 251326
rect 68928 251262 68980 251268
rect 68940 242865 68968 251262
rect 69124 251246 70058 251274
rect 68926 242856 68982 242865
rect 68926 242791 68982 242800
rect 64878 241632 64934 241641
rect 64878 241567 64934 241576
rect 64892 233238 64920 241567
rect 64880 233232 64932 233238
rect 64880 233174 64932 233180
rect 69124 230382 69152 251246
rect 90376 238754 90404 254050
rect 90456 254040 90508 254046
rect 90456 253982 90508 253988
rect 89824 238726 90404 238754
rect 89824 232778 89852 238726
rect 89378 232750 89852 232778
rect 69768 232070 70058 232098
rect 79718 232070 80008 232098
rect 69768 230450 69796 232070
rect 69756 230444 69808 230450
rect 69756 230386 69808 230392
rect 42800 230376 42852 230382
rect 42800 230318 42852 230324
rect 53104 230376 53156 230382
rect 53104 230318 53156 230324
rect 64144 230376 64196 230382
rect 64144 230318 64196 230324
rect 69112 230376 69164 230382
rect 69112 230318 69164 230324
rect 79980 230314 80008 232070
rect 90468 230314 90496 253982
rect 106660 251940 106688 254050
rect 116308 254040 116360 254046
rect 116308 253982 116360 253988
rect 116320 251940 116348 253982
rect 91100 251252 91152 251258
rect 91100 251194 91152 251200
rect 96724 251246 97014 251274
rect 91112 241641 91140 251194
rect 95146 242176 95202 242185
rect 95146 242111 95202 242120
rect 91098 241632 91154 241641
rect 91098 241567 91154 241576
rect 95160 233238 95188 242111
rect 95148 233232 95200 233238
rect 95148 233174 95200 233180
rect 96724 230450 96752 251246
rect 96816 232070 97014 232098
rect 106568 232070 106674 232098
rect 116228 232070 116334 232098
rect 96712 230444 96764 230450
rect 96712 230386 96764 230392
rect 96816 230382 96844 232070
rect 96804 230376 96856 230382
rect 96804 230318 96856 230324
rect 106568 230314 106596 232070
rect 116228 231962 116256 232070
rect 116504 231962 116532 254050
rect 116584 254040 116636 254046
rect 116584 253982 116636 253988
rect 116228 231934 116532 231962
rect 116596 230314 116624 253982
rect 133708 251940 133736 254050
rect 143356 254040 143408 254046
rect 143356 253982 143408 253988
rect 144276 254040 144328 254046
rect 144276 253982 144328 253988
rect 143368 251940 143396 253982
rect 144184 253972 144236 253978
rect 144184 253914 144236 253920
rect 118700 251320 118752 251326
rect 118700 251262 118752 251268
rect 122748 251320 122800 251326
rect 122748 251262 122800 251268
rect 118712 241641 118740 251262
rect 122760 242321 122788 251262
rect 122944 251246 124062 251274
rect 122746 242312 122802 242321
rect 122746 242247 122802 242256
rect 118698 241632 118754 241641
rect 118698 241567 118754 241576
rect 122944 230314 122972 251246
rect 144196 238754 144224 253914
rect 143736 238726 144224 238754
rect 143736 232778 143764 238726
rect 143382 232750 143764 232778
rect 123680 232070 124062 232098
rect 133722 232070 133828 232098
rect 123680 230382 123708 232070
rect 133800 230382 133828 232070
rect 144288 230382 144316 253982
rect 146298 241904 146354 241913
rect 146298 241839 146354 241848
rect 146312 233238 146340 241839
rect 146300 233232 146352 233238
rect 146300 233174 146352 233180
rect 146956 230450 146984 280434
rect 148968 277432 149020 277438
rect 148968 277374 149020 277380
rect 148980 269385 149008 277374
rect 148966 269376 149022 269385
rect 148966 269311 149022 269320
rect 149716 256630 149744 308042
rect 232044 308032 232096 308038
rect 232044 307974 232096 307980
rect 251824 308032 251876 308038
rect 251824 307974 251876 307980
rect 475016 308032 475068 308038
rect 475016 307974 475068 307980
rect 494704 308032 494756 308038
rect 494704 307974 494756 307980
rect 160652 307964 160704 307970
rect 160652 307906 160704 307912
rect 170496 307964 170548 307970
rect 170496 307906 170548 307912
rect 187700 307964 187752 307970
rect 187700 307906 187752 307912
rect 197452 307964 197504 307970
rect 197452 307906 197504 307912
rect 214656 307964 214708 307970
rect 214656 307906 214708 307912
rect 224500 307964 224552 307970
rect 224500 307906 224552 307912
rect 160664 305932 160692 307906
rect 170312 307896 170364 307902
rect 170312 307838 170364 307844
rect 170324 305932 170352 307838
rect 150544 305238 151018 305266
rect 150544 284238 150572 305238
rect 150532 284232 150584 284238
rect 150532 284174 150584 284180
rect 151004 284170 151032 286076
rect 150992 284164 151044 284170
rect 150992 284106 151044 284112
rect 160664 284102 160692 286076
rect 170324 285954 170352 286076
rect 170508 285954 170536 307906
rect 178040 307896 178092 307902
rect 178040 307838 178092 307844
rect 171784 307828 171836 307834
rect 171784 307770 171836 307776
rect 170324 285926 170536 285954
rect 171796 284102 171824 307770
rect 178052 305932 178080 307838
rect 187712 305932 187740 307906
rect 197360 307828 197412 307834
rect 197360 307770 197412 307776
rect 197372 305932 197400 307770
rect 176566 295760 176622 295769
rect 176566 295695 176622 295704
rect 172518 295624 172574 295633
rect 172518 295559 172574 295568
rect 172532 286958 172560 295559
rect 176580 286958 176608 295695
rect 172520 286952 172572 286958
rect 172520 286894 172572 286900
rect 176568 286952 176620 286958
rect 176568 286894 176620 286900
rect 197464 286770 197492 307906
rect 200764 307896 200816 307902
rect 200764 307838 200816 307844
rect 199384 307828 199436 307834
rect 199384 307770 199436 307776
rect 197386 286742 197492 286770
rect 178052 284170 178080 286076
rect 187712 284170 187740 286076
rect 199396 284170 199424 307770
rect 200118 295624 200174 295633
rect 200118 295559 200174 295568
rect 200132 287026 200160 295559
rect 200120 287020 200172 287026
rect 200120 286962 200172 286968
rect 200776 286822 200804 307838
rect 214668 305932 214696 307906
rect 224316 307828 224368 307834
rect 224316 307770 224368 307776
rect 224328 305932 224356 307770
rect 204364 305238 205022 305266
rect 202786 296304 202842 296313
rect 202786 296239 202842 296248
rect 202800 287026 202828 296239
rect 202788 287020 202840 287026
rect 202788 286962 202840 286968
rect 200764 286816 200816 286822
rect 200764 286758 200816 286764
rect 204364 284170 204392 305238
rect 204628 286816 204680 286822
rect 224512 286770 224540 307906
rect 225604 307828 225656 307834
rect 225604 307770 225656 307776
rect 204680 286764 205022 286770
rect 204628 286758 205022 286764
rect 204640 286742 205022 286758
rect 224342 286742 224540 286770
rect 178040 284164 178092 284170
rect 178040 284106 178092 284112
rect 187700 284164 187752 284170
rect 187700 284106 187752 284112
rect 199384 284164 199436 284170
rect 199384 284106 199436 284112
rect 204352 284164 204404 284170
rect 204352 284106 204404 284112
rect 214668 284102 214696 286076
rect 225616 284102 225644 307770
rect 232056 305932 232084 307974
rect 241704 307964 241756 307970
rect 241704 307906 241756 307912
rect 241716 305932 241744 307906
rect 251456 307896 251508 307902
rect 251456 307838 251508 307844
rect 251364 307828 251416 307834
rect 251364 307770 251416 307776
rect 251376 305932 251404 307770
rect 230386 296304 230442 296313
rect 230386 296239 230442 296248
rect 226338 295624 226394 295633
rect 226338 295559 226394 295568
rect 226352 286958 226380 295559
rect 230400 286958 230428 296239
rect 226340 286952 226392 286958
rect 226340 286894 226392 286900
rect 230388 286952 230440 286958
rect 230388 286894 230440 286900
rect 251468 286770 251496 307838
rect 251390 286742 251496 286770
rect 232056 284170 232084 286076
rect 241716 284170 241744 286076
rect 251836 284306 251864 307974
rect 413468 307964 413520 307970
rect 413468 307906 413520 307912
rect 430672 307964 430724 307970
rect 430672 307906 430724 307912
rect 440516 307964 440568 307970
rect 440516 307906 440568 307912
rect 457628 307964 457680 307970
rect 457628 307906 457680 307912
rect 468576 307964 468628 307970
rect 468576 307906 468628 307912
rect 268660 307896 268712 307902
rect 268660 307838 268712 307844
rect 279516 307896 279568 307902
rect 279516 307838 279568 307844
rect 295708 307896 295760 307902
rect 295708 307838 295760 307844
rect 305460 307896 305512 307902
rect 305460 307838 305512 307844
rect 322664 307896 322716 307902
rect 322664 307838 322716 307844
rect 334624 307896 334676 307902
rect 334624 307838 334676 307844
rect 349712 307896 349764 307902
rect 349712 307838 349764 307844
rect 359464 307896 359516 307902
rect 359464 307838 359516 307844
rect 376668 307896 376720 307902
rect 376668 307838 376720 307844
rect 386512 307896 386564 307902
rect 386512 307838 386564 307844
rect 403624 307896 403676 307902
rect 403624 307838 403676 307844
rect 253204 307828 253256 307834
rect 253204 307770 253256 307776
rect 251824 284300 251876 284306
rect 251824 284242 251876 284248
rect 253216 284170 253244 307770
rect 268672 305932 268700 307838
rect 278320 307828 278372 307834
rect 278320 307770 278372 307776
rect 279424 307828 279476 307834
rect 279424 307770 279476 307776
rect 278332 305932 278360 307770
rect 258184 305238 259026 305266
rect 256606 296304 256662 296313
rect 256606 296239 256662 296248
rect 253938 295352 253994 295361
rect 253938 295287 253994 295296
rect 253952 287026 253980 295287
rect 256620 287026 256648 296239
rect 253940 287020 253992 287026
rect 253940 286962 253992 286968
rect 256608 287020 256660 287026
rect 256608 286962 256660 286968
rect 258184 284170 258212 305238
rect 278688 286816 278740 286822
rect 278346 286764 278688 286770
rect 278346 286758 278740 286764
rect 278346 286742 278728 286758
rect 259012 284306 259040 286076
rect 259000 284300 259052 284306
rect 259000 284242 259052 284248
rect 232044 284164 232096 284170
rect 232044 284106 232096 284112
rect 241704 284164 241756 284170
rect 241704 284106 241756 284112
rect 253204 284164 253256 284170
rect 253204 284106 253256 284112
rect 258172 284164 258224 284170
rect 258172 284106 258224 284112
rect 268672 284102 268700 286076
rect 279436 284102 279464 307770
rect 279528 286822 279556 307838
rect 285784 306054 286088 306082
rect 284206 295760 284262 295769
rect 284206 295695 284262 295704
rect 280158 295624 280214 295633
rect 280158 295559 280214 295568
rect 280172 286958 280200 295559
rect 284220 286958 284248 295695
rect 280160 286952 280212 286958
rect 280160 286894 280212 286900
rect 284208 286952 284260 286958
rect 284208 286894 284260 286900
rect 279516 286816 279568 286822
rect 279516 286758 279568 286764
rect 285784 284102 285812 306054
rect 286060 305932 286088 306054
rect 295720 305932 295748 307838
rect 305368 307828 305420 307834
rect 305368 307770 305420 307776
rect 305380 305932 305408 307770
rect 305472 286770 305500 307838
rect 307024 307828 307076 307834
rect 307024 307770 307076 307776
rect 305394 286742 305500 286770
rect 286060 284170 286088 286076
rect 286048 284164 286100 284170
rect 286048 284106 286100 284112
rect 295720 284102 295748 286076
rect 307036 284102 307064 307770
rect 322676 305932 322704 307838
rect 332324 307828 332376 307834
rect 332324 307770 332376 307776
rect 333244 307828 333296 307834
rect 333244 307770 333296 307776
rect 332336 305932 332364 307770
rect 312004 305238 313030 305266
rect 311806 296304 311862 296313
rect 311806 296239 311862 296248
rect 307758 295624 307814 295633
rect 307758 295559 307814 295568
rect 307772 287026 307800 295559
rect 307760 287020 307812 287026
rect 307760 286962 307812 286968
rect 311820 286890 311848 296239
rect 311808 286884 311860 286890
rect 311808 286826 311860 286832
rect 312004 284102 312032 305238
rect 332508 286816 332560 286822
rect 332350 286764 332508 286770
rect 332350 286758 332560 286764
rect 332350 286742 332548 286758
rect 313016 284170 313044 286076
rect 313004 284164 313056 284170
rect 313004 284106 313056 284112
rect 322676 284102 322704 286076
rect 333256 284102 333284 307770
rect 334636 286822 334664 307838
rect 339604 306054 340092 306082
rect 338026 296304 338082 296313
rect 338026 296239 338082 296248
rect 335358 295624 335414 295633
rect 335358 295559 335414 295568
rect 335372 286958 335400 295559
rect 338040 287026 338068 296239
rect 338028 287020 338080 287026
rect 338028 286962 338080 286968
rect 335360 286952 335412 286958
rect 335360 286894 335412 286900
rect 334624 286816 334676 286822
rect 334624 286758 334676 286764
rect 339604 284102 339632 306054
rect 340064 305932 340092 306054
rect 349724 305932 349752 307838
rect 359372 307828 359424 307834
rect 359372 307770 359424 307776
rect 359384 305932 359412 307770
rect 359476 286770 359504 307838
rect 359556 307828 359608 307834
rect 359556 307770 359608 307776
rect 359398 286742 359504 286770
rect 340064 284170 340092 286076
rect 340052 284164 340104 284170
rect 340052 284106 340104 284112
rect 349724 284102 349752 286076
rect 359568 284102 359596 307770
rect 376680 305932 376708 307838
rect 386328 307828 386380 307834
rect 386328 307770 386380 307776
rect 386340 305932 386368 307770
rect 365824 305238 367034 305266
rect 365626 296304 365682 296313
rect 365626 296239 365682 296248
rect 361578 295352 361634 295361
rect 361578 295287 361634 295296
rect 361592 286890 361620 295287
rect 365640 286958 365668 296239
rect 365628 286952 365680 286958
rect 365628 286894 365680 286900
rect 361580 286884 361632 286890
rect 361580 286826 361632 286832
rect 365824 284102 365852 305238
rect 386524 286770 386552 307838
rect 387064 307828 387116 307834
rect 387064 307770 387116 307776
rect 386354 286742 386552 286770
rect 367020 284170 367048 286076
rect 367008 284164 367060 284170
rect 367008 284106 367060 284112
rect 376680 284102 376708 286076
rect 387076 284102 387104 307770
rect 403636 305932 403664 307838
rect 413284 307828 413336 307834
rect 413284 307770 413336 307776
rect 413296 305932 413324 307770
rect 393424 305238 393990 305266
rect 391846 296304 391902 296313
rect 391846 296239 391902 296248
rect 389178 295624 389234 295633
rect 389178 295559 389234 295568
rect 389192 287026 389220 295559
rect 391860 287026 391888 296239
rect 389180 287020 389232 287026
rect 389180 286962 389232 286968
rect 391848 287020 391900 287026
rect 391848 286962 391900 286968
rect 393424 284102 393452 305238
rect 413480 286770 413508 307906
rect 421012 307896 421064 307902
rect 421012 307838 421064 307844
rect 414664 307828 414716 307834
rect 414664 307770 414716 307776
rect 413402 286742 413508 286770
rect 393976 284170 394004 286076
rect 393964 284164 394016 284170
rect 393964 284106 394016 284112
rect 403728 284102 403756 286076
rect 414676 284102 414704 307770
rect 421024 305932 421052 307838
rect 430684 305932 430712 307906
rect 440332 307828 440384 307834
rect 440332 307770 440384 307776
rect 440344 305932 440372 307770
rect 419446 296304 419502 296313
rect 419446 296239 419502 296248
rect 415398 295624 415454 295633
rect 415398 295559 415454 295568
rect 415412 286958 415440 295559
rect 419460 286958 419488 296239
rect 415400 286952 415452 286958
rect 415400 286894 415452 286900
rect 419448 286952 419500 286958
rect 419448 286894 419500 286900
rect 440528 286770 440556 307906
rect 443644 307896 443696 307902
rect 443644 307838 443696 307844
rect 442264 307828 442316 307834
rect 442264 307770 442316 307776
rect 440358 286742 440556 286770
rect 421024 284170 421052 286076
rect 430684 284170 430712 286076
rect 442276 284170 442304 307770
rect 442998 295624 443054 295633
rect 442998 295559 443054 295568
rect 443012 287026 443040 295559
rect 443000 287020 443052 287026
rect 443000 286962 443052 286968
rect 443656 284306 443684 307838
rect 457640 305932 457668 307906
rect 467288 307828 467340 307834
rect 467288 307770 467340 307776
rect 468484 307828 468536 307834
rect 468484 307770 468536 307776
rect 467300 305932 467328 307770
rect 447244 305238 447994 305266
rect 445666 296304 445722 296313
rect 445666 296239 445722 296248
rect 445680 287026 445708 296239
rect 445668 287020 445720 287026
rect 445668 286962 445720 286968
rect 443644 284300 443696 284306
rect 443644 284242 443696 284248
rect 447244 284170 447272 305238
rect 467656 286816 467708 286822
rect 467406 286764 467656 286770
rect 467406 286758 467708 286764
rect 467406 286742 467696 286758
rect 447980 284306 448008 286076
rect 447968 284300 448020 284306
rect 447968 284242 448020 284248
rect 421012 284164 421064 284170
rect 421012 284106 421064 284112
rect 430672 284164 430724 284170
rect 430672 284106 430724 284112
rect 442264 284164 442316 284170
rect 442264 284106 442316 284112
rect 447232 284164 447284 284170
rect 447232 284106 447284 284112
rect 457732 284102 457760 286076
rect 468496 284102 468524 307770
rect 468588 286822 468616 307906
rect 475028 305932 475056 307974
rect 484676 307964 484728 307970
rect 484676 307906 484728 307912
rect 484688 305932 484716 307906
rect 494520 307896 494572 307902
rect 494520 307838 494572 307844
rect 494336 307828 494388 307834
rect 494336 307770 494388 307776
rect 494348 305932 494376 307770
rect 473266 295760 473322 295769
rect 473266 295695 473322 295704
rect 469218 295352 469274 295361
rect 469218 295287 469274 295296
rect 469232 286958 469260 295287
rect 473280 286958 473308 295695
rect 469220 286952 469272 286958
rect 469220 286894 469272 286900
rect 473268 286952 473320 286958
rect 473268 286894 473320 286900
rect 468576 286816 468628 286822
rect 494532 286770 494560 307838
rect 468576 286758 468628 286764
rect 494362 286742 494560 286770
rect 475028 284170 475056 286076
rect 484688 284170 484716 286076
rect 494716 284306 494744 307974
rect 511632 307896 511684 307902
rect 511632 307838 511684 307844
rect 522304 307896 522356 307902
rect 522304 307838 522356 307844
rect 496084 307828 496136 307834
rect 496084 307770 496136 307776
rect 494704 284300 494756 284306
rect 494704 284242 494756 284248
rect 496096 284170 496124 307770
rect 511644 305932 511672 307838
rect 521292 307828 521344 307834
rect 521292 307770 521344 307776
rect 521304 305932 521332 307770
rect 501064 305238 501998 305266
rect 500866 296304 500922 296313
rect 500866 296239 500922 296248
rect 496818 295624 496874 295633
rect 496818 295559 496874 295568
rect 496832 287026 496860 295559
rect 500880 287026 500908 296239
rect 496820 287020 496872 287026
rect 496820 286962 496872 286968
rect 500868 287020 500920 287026
rect 500868 286962 500920 286968
rect 501064 284170 501092 305238
rect 522316 287054 522344 307838
rect 522396 307828 522448 307834
rect 522396 307770 522448 307776
rect 521856 287026 522344 287054
rect 521856 286770 521884 287026
rect 521410 286742 521884 286770
rect 501984 284306 502012 286076
rect 501972 284300 502024 284306
rect 501972 284242 502024 284248
rect 475016 284164 475068 284170
rect 475016 284106 475068 284112
rect 484676 284164 484728 284170
rect 484676 284106 484728 284112
rect 496084 284164 496136 284170
rect 496084 284106 496136 284112
rect 501052 284164 501104 284170
rect 501052 284106 501104 284112
rect 511736 284102 511764 286076
rect 522408 284102 522436 307770
rect 529032 305932 529060 308382
rect 538680 307896 538732 307902
rect 538680 307838 538732 307844
rect 538692 305932 538720 307838
rect 548340 307828 548392 307834
rect 548340 307770 548392 307776
rect 548352 305932 548380 307770
rect 526444 305652 526496 305658
rect 526444 305594 526496 305600
rect 526456 296313 526484 305594
rect 526442 296304 526498 296313
rect 526442 296239 526498 296248
rect 523038 295624 523094 295633
rect 523038 295559 523094 295568
rect 550638 295624 550694 295633
rect 550638 295559 550694 295568
rect 523052 286958 523080 295559
rect 550652 287026 550680 295559
rect 550640 287020 550692 287026
rect 550640 286962 550692 286968
rect 523040 286952 523092 286958
rect 523040 286894 523092 286900
rect 529032 284170 529060 286076
rect 529020 284164 529072 284170
rect 529020 284106 529072 284112
rect 160652 284096 160704 284102
rect 160652 284038 160704 284044
rect 171784 284096 171836 284102
rect 171784 284038 171836 284044
rect 214656 284096 214708 284102
rect 214656 284038 214708 284044
rect 225604 284096 225656 284102
rect 225604 284038 225656 284044
rect 268660 284096 268712 284102
rect 268660 284038 268712 284044
rect 279424 284096 279476 284102
rect 279424 284038 279476 284044
rect 285772 284096 285824 284102
rect 285772 284038 285824 284044
rect 295708 284096 295760 284102
rect 295708 284038 295760 284044
rect 307024 284096 307076 284102
rect 307024 284038 307076 284044
rect 311992 284096 312044 284102
rect 311992 284038 312044 284044
rect 322664 284096 322716 284102
rect 322664 284038 322716 284044
rect 333244 284096 333296 284102
rect 333244 284038 333296 284044
rect 339592 284096 339644 284102
rect 339592 284038 339644 284044
rect 349712 284096 349764 284102
rect 349712 284038 349764 284044
rect 359556 284096 359608 284102
rect 359556 284038 359608 284044
rect 365812 284096 365864 284102
rect 365812 284038 365864 284044
rect 376668 284096 376720 284102
rect 376668 284038 376720 284044
rect 387064 284096 387116 284102
rect 387064 284038 387116 284044
rect 393412 284096 393464 284102
rect 393412 284038 393464 284044
rect 403716 284096 403768 284102
rect 403716 284038 403768 284044
rect 414664 284096 414716 284102
rect 414664 284038 414716 284044
rect 457720 284096 457772 284102
rect 457720 284038 457772 284044
rect 468484 284096 468536 284102
rect 468484 284038 468536 284044
rect 511724 284096 511776 284102
rect 511724 284038 511776 284044
rect 522396 284096 522448 284102
rect 522396 284038 522448 284044
rect 538692 284034 538720 286076
rect 548352 284238 548380 286076
rect 548340 284232 548392 284238
rect 548340 284174 548392 284180
rect 538680 284028 538732 284034
rect 538680 283970 538732 283976
rect 528744 280832 528796 280838
rect 528744 280774 528796 280780
rect 232320 280424 232372 280430
rect 232320 280366 232372 280372
rect 251824 280424 251876 280430
rect 251824 280366 251876 280372
rect 475384 280424 475436 280430
rect 475384 280366 475436 280372
rect 494704 280424 494756 280430
rect 494704 280366 494756 280372
rect 170496 280356 170548 280362
rect 170496 280298 170548 280304
rect 187792 280356 187844 280362
rect 187792 280298 187844 280304
rect 197544 280356 197596 280362
rect 197544 280298 197596 280304
rect 214380 280356 214432 280362
rect 214380 280298 214432 280304
rect 224500 280356 224552 280362
rect 224500 280298 224552 280304
rect 170036 280288 170088 280294
rect 170036 280230 170088 280236
rect 160284 280220 160336 280226
rect 160284 280162 160336 280168
rect 160296 278882 160324 280162
rect 170048 278882 170076 280230
rect 160296 278854 160678 278882
rect 170048 278854 170338 278882
rect 150544 278310 151018 278338
rect 149704 256624 149756 256630
rect 149704 256566 149756 256572
rect 150544 256562 150572 278310
rect 170232 259690 170338 259706
rect 170508 259690 170536 280298
rect 178408 280288 178460 280294
rect 178408 280230 178460 280236
rect 171784 280220 171836 280226
rect 171784 280162 171836 280168
rect 170220 259684 170338 259690
rect 170272 259678 170338 259684
rect 170496 259684 170548 259690
rect 170220 259626 170272 259632
rect 170496 259626 170548 259632
rect 150728 259134 151018 259162
rect 160572 259134 160678 259162
rect 150532 256556 150584 256562
rect 150532 256498 150584 256504
rect 150728 256494 150756 259134
rect 160572 256494 160600 259134
rect 171796 256494 171824 280162
rect 178420 278882 178448 280230
rect 187804 278882 187832 280298
rect 197452 280220 197504 280226
rect 197452 280162 197504 280168
rect 197464 278882 197492 280162
rect 178066 278854 178448 278882
rect 187726 278854 187832 278882
rect 197386 278854 197492 278882
rect 172520 277500 172572 277506
rect 172520 277442 172572 277448
rect 176568 277500 176620 277506
rect 176568 277442 176620 277448
rect 172532 268705 172560 277442
rect 176580 269929 176608 277442
rect 176566 269920 176622 269929
rect 176566 269855 176622 269864
rect 172518 268696 172574 268705
rect 172518 268631 172574 268640
rect 197556 259706 197584 280298
rect 200764 280288 200816 280294
rect 200764 280230 200816 280236
rect 199384 280220 199436 280226
rect 199384 280162 199436 280168
rect 197386 259678 197584 259706
rect 178066 259134 178172 259162
rect 187726 259134 188016 259162
rect 178144 256562 178172 259134
rect 187988 256562 188016 259134
rect 199396 256562 199424 280162
rect 200120 277432 200172 277438
rect 200120 277374 200172 277380
rect 200132 268705 200160 277374
rect 200118 268696 200174 268705
rect 200118 268631 200174 268640
rect 200776 256698 200804 280230
rect 214392 278882 214420 280298
rect 223948 280220 224000 280226
rect 223948 280162 224000 280168
rect 223960 278882 223988 280162
rect 214392 278854 214682 278882
rect 223960 278854 224342 278882
rect 204364 278310 205022 278338
rect 202788 277432 202840 277438
rect 202788 277374 202840 277380
rect 202800 269385 202828 277374
rect 202786 269376 202842 269385
rect 202786 269311 202842 269320
rect 200764 256692 200816 256698
rect 200764 256634 200816 256640
rect 204364 256562 204392 278310
rect 224512 259706 224540 280298
rect 225604 280220 225656 280226
rect 225604 280162 225656 280168
rect 224342 259678 224540 259706
rect 204640 259134 205022 259162
rect 214682 259134 215064 259162
rect 204640 256698 204668 259134
rect 204628 256692 204680 256698
rect 204628 256634 204680 256640
rect 178132 256556 178184 256562
rect 178132 256498 178184 256504
rect 187976 256556 188028 256562
rect 187976 256498 188028 256504
rect 199384 256556 199436 256562
rect 199384 256498 199436 256504
rect 204352 256556 204404 256562
rect 204352 256498 204404 256504
rect 215036 256494 215064 259134
rect 225616 256494 225644 280162
rect 232332 278882 232360 280366
rect 241520 280356 241572 280362
rect 241520 280298 241572 280304
rect 232070 278854 232360 278882
rect 241532 278882 241560 280298
rect 251456 280288 251508 280294
rect 251456 280230 251508 280236
rect 251180 280220 251232 280226
rect 251180 280162 251232 280168
rect 251192 278882 251220 280162
rect 241532 278854 241730 278882
rect 251192 278854 251390 278882
rect 226340 277500 226392 277506
rect 226340 277442 226392 277448
rect 230388 277500 230440 277506
rect 230388 277442 230440 277448
rect 226352 268705 226380 277442
rect 230400 269385 230428 277442
rect 230386 269376 230442 269385
rect 230386 269311 230442 269320
rect 226338 268696 226394 268705
rect 226338 268631 226394 268640
rect 251468 259706 251496 280230
rect 251390 259678 251496 259706
rect 231964 259134 232070 259162
rect 241730 259134 242112 259162
rect 231964 256562 231992 259134
rect 242084 256562 242112 259134
rect 251836 256698 251864 280366
rect 413468 280356 413520 280362
rect 413468 280298 413520 280304
rect 430580 280356 430632 280362
rect 430580 280298 430632 280304
rect 440516 280356 440568 280362
rect 440516 280298 440568 280304
rect 457260 280356 457312 280362
rect 457260 280298 457312 280304
rect 468576 280356 468628 280362
rect 468576 280298 468628 280304
rect 268292 280288 268344 280294
rect 268292 280230 268344 280236
rect 279516 280288 279568 280294
rect 279516 280230 279568 280236
rect 295800 280288 295852 280294
rect 295800 280230 295852 280236
rect 305552 280288 305604 280294
rect 305552 280230 305604 280236
rect 322388 280288 322440 280294
rect 322388 280230 322440 280236
rect 336004 280288 336056 280294
rect 336004 280230 336056 280236
rect 349804 280288 349856 280294
rect 349804 280230 349856 280236
rect 359648 280288 359700 280294
rect 359648 280230 359700 280236
rect 376300 280288 376352 280294
rect 376300 280230 376352 280236
rect 386512 280288 386564 280294
rect 386512 280230 386564 280236
rect 403348 280288 403400 280294
rect 403348 280230 403400 280236
rect 253204 280220 253256 280226
rect 253204 280162 253256 280168
rect 251824 256692 251876 256698
rect 251824 256634 251876 256640
rect 253216 256562 253244 280162
rect 268304 278882 268332 280230
rect 278044 280220 278096 280226
rect 278044 280162 278096 280168
rect 279424 280220 279476 280226
rect 279424 280162 279476 280168
rect 278056 278882 278084 280162
rect 268304 278854 268686 278882
rect 278056 278854 278346 278882
rect 258184 278310 259026 278338
rect 253940 277432 253992 277438
rect 253940 277374 253992 277380
rect 256608 277432 256660 277438
rect 256608 277374 256660 277380
rect 253952 269113 253980 277374
rect 256620 269385 256648 277374
rect 256606 269376 256662 269385
rect 256606 269311 256662 269320
rect 253938 269104 253994 269113
rect 253938 269039 253994 269048
rect 258184 256562 258212 278310
rect 278346 259418 278728 259434
rect 278346 259412 278740 259418
rect 278346 259406 278688 259412
rect 278688 259354 278740 259360
rect 258736 259134 259026 259162
rect 268686 259134 268976 259162
rect 258736 256698 258764 259134
rect 258724 256692 258776 256698
rect 258724 256634 258776 256640
rect 231952 256556 232004 256562
rect 231952 256498 232004 256504
rect 242072 256556 242124 256562
rect 242072 256498 242124 256504
rect 253204 256556 253256 256562
rect 253204 256498 253256 256504
rect 258172 256556 258224 256562
rect 258172 256498 258224 256504
rect 268948 256494 268976 259134
rect 279436 256494 279464 280162
rect 279528 259418 279556 280230
rect 295812 278882 295840 280230
rect 305460 280220 305512 280226
rect 305460 280162 305512 280168
rect 305472 278882 305500 280162
rect 295734 278854 295840 278882
rect 305394 278854 305500 278882
rect 286074 278322 286180 278338
rect 285772 278316 285824 278322
rect 286074 278316 286192 278322
rect 286074 278310 286140 278316
rect 285772 278258 285824 278264
rect 286140 278258 286192 278264
rect 280160 277500 280212 277506
rect 280160 277442 280212 277448
rect 284208 277500 284260 277506
rect 284208 277442 284260 277448
rect 280172 268705 280200 277442
rect 284220 269929 284248 277442
rect 284206 269920 284262 269929
rect 284206 269855 284262 269864
rect 280158 268696 280214 268705
rect 280158 268631 280214 268640
rect 279516 259412 279568 259418
rect 279516 259354 279568 259360
rect 285784 256562 285812 278258
rect 305564 277394 305592 280230
rect 307024 280220 307076 280226
rect 307024 280162 307076 280168
rect 305472 277366 305592 277394
rect 305472 259706 305500 277366
rect 305394 259678 305500 259706
rect 286074 259134 286180 259162
rect 295734 259134 296024 259162
rect 285772 256556 285824 256562
rect 285772 256498 285824 256504
rect 286152 256494 286180 259134
rect 295996 256494 296024 259134
rect 307036 256494 307064 280162
rect 322400 278882 322428 280230
rect 331956 280220 332008 280226
rect 331956 280162 332008 280168
rect 333244 280220 333296 280226
rect 333244 280162 333296 280168
rect 331968 278882 331996 280162
rect 322400 278854 322690 278882
rect 331968 278854 332350 278882
rect 312004 278310 313030 278338
rect 311808 277568 311860 277574
rect 311808 277510 311860 277516
rect 307760 277432 307812 277438
rect 307760 277374 307812 277380
rect 307772 268705 307800 277374
rect 311820 269385 311848 277510
rect 311806 269376 311862 269385
rect 311806 269311 311862 269320
rect 307758 268696 307814 268705
rect 307758 268631 307814 268640
rect 312004 256494 312032 278310
rect 332350 259418 332640 259434
rect 332350 259412 332652 259418
rect 332350 259406 332600 259412
rect 332600 259354 332652 259360
rect 312648 259134 313030 259162
rect 322690 259134 322888 259162
rect 312648 256562 312676 259134
rect 312636 256556 312688 256562
rect 312636 256498 312688 256504
rect 322860 256494 322888 259134
rect 333256 256494 333284 280162
rect 335360 277500 335412 277506
rect 335360 277442 335412 277448
rect 335372 268705 335400 277442
rect 335358 268696 335414 268705
rect 335358 268631 335414 268640
rect 336016 259418 336044 280230
rect 349816 278882 349844 280230
rect 359464 280220 359516 280226
rect 359464 280162 359516 280168
rect 359476 278882 359504 280162
rect 349738 278854 349844 278882
rect 359398 278854 359504 278882
rect 359660 278610 359688 280230
rect 359740 280220 359792 280226
rect 359740 280162 359792 280168
rect 359476 278582 359688 278610
rect 340078 278322 340184 278338
rect 339592 278316 339644 278322
rect 340078 278316 340196 278322
rect 340078 278310 340144 278316
rect 339592 278258 339644 278264
rect 340144 278258 340196 278264
rect 338028 277432 338080 277438
rect 338028 277374 338080 277380
rect 338040 269385 338068 277374
rect 338026 269376 338082 269385
rect 338026 269311 338082 269320
rect 336004 259412 336056 259418
rect 336004 259354 336056 259360
rect 339604 256494 339632 278258
rect 359476 259706 359504 278582
rect 359752 277394 359780 280162
rect 376312 278882 376340 280230
rect 386052 280220 386104 280226
rect 386052 280162 386104 280168
rect 386064 278882 386092 280162
rect 376312 278854 376694 278882
rect 386064 278854 386354 278882
rect 365824 278310 367034 278338
rect 361580 277568 361632 277574
rect 361580 277510 361632 277516
rect 359398 259678 359504 259706
rect 359568 277366 359780 277394
rect 340078 259134 340184 259162
rect 349738 259134 350120 259162
rect 340156 256562 340184 259134
rect 340144 256556 340196 256562
rect 340144 256498 340196 256504
rect 350092 256494 350120 259134
rect 359568 256494 359596 277366
rect 361592 269113 361620 277510
rect 365628 277500 365680 277506
rect 365628 277442 365680 277448
rect 365640 269385 365668 277442
rect 365626 269376 365682 269385
rect 365626 269311 365682 269320
rect 361578 269104 361634 269113
rect 361578 269039 361634 269048
rect 365824 256562 365852 278310
rect 386524 259706 386552 280230
rect 387064 280220 387116 280226
rect 387064 280162 387116 280168
rect 386354 259678 386552 259706
rect 366744 259134 367034 259162
rect 376588 259134 376694 259162
rect 365812 256556 365864 256562
rect 365812 256498 365864 256504
rect 366744 256494 366772 259134
rect 376588 256494 376616 259134
rect 387076 256494 387104 280162
rect 403360 278882 403388 280230
rect 412916 280220 412968 280226
rect 412916 280162 412968 280168
rect 412928 278882 412956 280162
rect 403360 278854 403650 278882
rect 412928 278854 413310 278882
rect 393424 278310 393990 278338
rect 389180 277432 389232 277438
rect 389180 277374 389232 277380
rect 391848 277432 391900 277438
rect 391848 277374 391900 277380
rect 389192 268705 389220 277374
rect 391860 269385 391888 277374
rect 391846 269376 391902 269385
rect 391846 269311 391902 269320
rect 389178 268696 389234 268705
rect 389178 268631 389234 268640
rect 393424 256494 393452 278310
rect 413480 259706 413508 280298
rect 421288 280288 421340 280294
rect 421288 280230 421340 280236
rect 414664 280220 414716 280226
rect 414664 280162 414716 280168
rect 413402 259678 413508 259706
rect 393608 259134 393990 259162
rect 403742 259134 404032 259162
rect 393608 256562 393636 259134
rect 393596 256556 393648 256562
rect 393596 256498 393648 256504
rect 404004 256494 404032 259134
rect 414676 256494 414704 280162
rect 421300 278882 421328 280230
rect 421038 278854 421328 278882
rect 430592 278882 430620 280298
rect 440240 280220 440292 280226
rect 440240 280162 440292 280168
rect 440252 278882 440280 280162
rect 430592 278854 430698 278882
rect 440252 278854 440358 278882
rect 415400 277500 415452 277506
rect 415400 277442 415452 277448
rect 419448 277500 419500 277506
rect 419448 277442 419500 277448
rect 415412 268705 415440 277442
rect 419460 269385 419488 277442
rect 419446 269376 419502 269385
rect 419446 269311 419502 269320
rect 415398 268696 415454 268705
rect 415398 268631 415454 268640
rect 440528 259706 440556 280298
rect 446404 280288 446456 280294
rect 446404 280230 446456 280236
rect 442264 280220 442316 280226
rect 442264 280162 442316 280168
rect 440358 259678 440556 259706
rect 420932 259134 421038 259162
rect 430698 259134 431080 259162
rect 420932 256562 420960 259134
rect 431052 256562 431080 259134
rect 442276 256562 442304 280162
rect 443000 277432 443052 277438
rect 443000 277374 443052 277380
rect 445668 277432 445720 277438
rect 445668 277374 445720 277380
rect 443012 268705 443040 277374
rect 445680 269385 445708 277374
rect 445666 269376 445722 269385
rect 445666 269311 445722 269320
rect 442998 268696 443054 268705
rect 442998 268631 443054 268640
rect 446416 259486 446444 280230
rect 457272 278882 457300 280298
rect 467012 280220 467064 280226
rect 467012 280162 467064 280168
rect 468484 280220 468536 280226
rect 468484 280162 468536 280168
rect 467024 278882 467052 280162
rect 457272 278854 457654 278882
rect 467024 278854 467314 278882
rect 447244 278310 447994 278338
rect 446404 259480 446456 259486
rect 446404 259422 446456 259428
rect 447244 256562 447272 278310
rect 447692 259480 447744 259486
rect 447744 259428 447994 259434
rect 447692 259422 447994 259428
rect 447704 259406 447994 259422
rect 467406 259418 467696 259434
rect 467406 259412 467708 259418
rect 467406 259406 467656 259412
rect 467656 259354 467708 259360
rect 457746 259134 458128 259162
rect 420920 256556 420972 256562
rect 420920 256498 420972 256504
rect 431040 256556 431092 256562
rect 431040 256498 431092 256504
rect 442264 256556 442316 256562
rect 442264 256498 442316 256504
rect 447232 256556 447284 256562
rect 447232 256498 447284 256504
rect 458100 256494 458128 259134
rect 468496 256494 468524 280162
rect 468588 259418 468616 280298
rect 475396 278882 475424 280366
rect 484400 280356 484452 280362
rect 484400 280298 484452 280304
rect 475042 278854 475424 278882
rect 484412 278882 484440 280298
rect 494520 280288 494572 280294
rect 494520 280230 494572 280236
rect 494060 280220 494112 280226
rect 494060 280162 494112 280168
rect 494072 278882 494100 280162
rect 484412 278854 484702 278882
rect 494072 278854 494362 278882
rect 469220 277500 469272 277506
rect 469220 277442 469272 277448
rect 473268 277500 473320 277506
rect 473268 277442 473320 277448
rect 469232 269113 469260 277442
rect 473280 269929 473308 277442
rect 473266 269920 473322 269929
rect 473266 269855 473322 269864
rect 469218 269104 469274 269113
rect 469218 269039 469274 269048
rect 494532 259706 494560 280230
rect 494362 259678 494560 259706
rect 468576 259412 468628 259418
rect 468576 259354 468628 259360
rect 474752 259134 475042 259162
rect 484702 259134 484992 259162
rect 474752 256562 474780 259134
rect 484964 256562 484992 259134
rect 494716 256698 494744 280366
rect 511356 280288 511408 280294
rect 511356 280230 511408 280236
rect 522304 280288 522356 280294
rect 522304 280230 522356 280236
rect 496084 280220 496136 280226
rect 496084 280162 496136 280168
rect 494704 256692 494756 256698
rect 494704 256634 494756 256640
rect 496096 256562 496124 280162
rect 511368 278882 511396 280230
rect 520924 280220 520976 280226
rect 520924 280162 520976 280168
rect 520936 278882 520964 280162
rect 511368 278854 511658 278882
rect 520936 278854 521318 278882
rect 501064 278310 501998 278338
rect 496820 277432 496872 277438
rect 496820 277374 496872 277380
rect 500868 277432 500920 277438
rect 500868 277374 500920 277380
rect 496832 268705 496860 277374
rect 500880 269385 500908 277374
rect 500866 269376 500922 269385
rect 500866 269311 500922 269320
rect 496818 268696 496874 268705
rect 496818 268631 496874 268640
rect 501064 256562 501092 278310
rect 522316 267734 522344 280230
rect 522396 280220 522448 280226
rect 522396 280162 522448 280168
rect 521856 267706 522344 267734
rect 521856 259434 521884 267706
rect 521410 259406 521884 259434
rect 501616 259134 501998 259162
rect 511750 259134 511856 259162
rect 501616 256698 501644 259134
rect 501604 256692 501656 256698
rect 501604 256634 501656 256640
rect 474740 256556 474792 256562
rect 474740 256498 474792 256504
rect 484952 256556 485004 256562
rect 484952 256498 485004 256504
rect 496084 256556 496136 256562
rect 496084 256498 496136 256504
rect 501052 256556 501104 256562
rect 501052 256498 501104 256504
rect 511828 256494 511856 259134
rect 522408 256494 522436 280162
rect 526444 279472 526496 279478
rect 526444 279414 526496 279420
rect 523040 277500 523092 277506
rect 523040 277442 523092 277448
rect 523052 268705 523080 277442
rect 526456 269385 526484 279414
rect 528756 278882 528784 280774
rect 538404 280288 538456 280294
rect 538404 280230 538456 280236
rect 538416 278882 538444 280230
rect 548064 280220 548116 280226
rect 548064 280162 548116 280168
rect 548076 278882 548104 280162
rect 528756 278854 529046 278882
rect 538416 278854 538706 278882
rect 548076 278854 548366 278882
rect 550640 277432 550692 277438
rect 550640 277374 550692 277380
rect 526442 269376 526498 269385
rect 526442 269311 526498 269320
rect 550652 268705 550680 277374
rect 523038 268696 523094 268705
rect 523038 268631 523094 268640
rect 550638 268696 550694 268705
rect 550638 268631 550694 268640
rect 528664 259134 529046 259162
rect 538416 259134 538706 259162
rect 547984 259134 548366 259162
rect 528664 256562 528692 259134
rect 528652 256556 528704 256562
rect 528652 256498 528704 256504
rect 150716 256488 150768 256494
rect 150716 256430 150768 256436
rect 160560 256488 160612 256494
rect 160560 256430 160612 256436
rect 171784 256488 171836 256494
rect 171784 256430 171836 256436
rect 215024 256488 215076 256494
rect 215024 256430 215076 256436
rect 225604 256488 225656 256494
rect 225604 256430 225656 256436
rect 268936 256488 268988 256494
rect 268936 256430 268988 256436
rect 279424 256488 279476 256494
rect 279424 256430 279476 256436
rect 286140 256488 286192 256494
rect 286140 256430 286192 256436
rect 295984 256488 296036 256494
rect 295984 256430 296036 256436
rect 307024 256488 307076 256494
rect 307024 256430 307076 256436
rect 311992 256488 312044 256494
rect 311992 256430 312044 256436
rect 322848 256488 322900 256494
rect 322848 256430 322900 256436
rect 333244 256488 333296 256494
rect 333244 256430 333296 256436
rect 339592 256488 339644 256494
rect 339592 256430 339644 256436
rect 350080 256488 350132 256494
rect 350080 256430 350132 256436
rect 359556 256488 359608 256494
rect 359556 256430 359608 256436
rect 366732 256488 366784 256494
rect 366732 256430 366784 256436
rect 376576 256488 376628 256494
rect 376576 256430 376628 256436
rect 387064 256488 387116 256494
rect 387064 256430 387116 256436
rect 393412 256488 393464 256494
rect 393412 256430 393464 256436
rect 403992 256488 404044 256494
rect 403992 256430 404044 256436
rect 414664 256488 414716 256494
rect 414664 256430 414716 256436
rect 458088 256488 458140 256494
rect 458088 256430 458140 256436
rect 468484 256488 468536 256494
rect 468484 256430 468536 256436
rect 511816 256488 511868 256494
rect 511816 256430 511868 256436
rect 522396 256488 522448 256494
rect 522396 256430 522448 256436
rect 538416 256426 538444 259134
rect 547984 256630 548012 259134
rect 547972 256624 548024 256630
rect 547972 256566 548024 256572
rect 538404 256420 538456 256426
rect 538404 256362 538456 256368
rect 529020 254584 529072 254590
rect 529020 254526 529072 254532
rect 148324 254244 148376 254250
rect 148324 254186 148376 254192
rect 146944 230444 146996 230450
rect 146944 230386 146996 230392
rect 123668 230376 123720 230382
rect 123668 230318 123720 230324
rect 133788 230376 133840 230382
rect 133788 230318 133840 230324
rect 144276 230376 144328 230382
rect 144276 230318 144328 230324
rect 79968 230308 80020 230314
rect 79968 230250 80020 230256
rect 90456 230308 90508 230314
rect 90456 230250 90508 230256
rect 106556 230308 106608 230314
rect 106556 230250 106608 230256
rect 116584 230308 116636 230314
rect 116584 230250 116636 230256
rect 122932 230308 122984 230314
rect 122932 230250 122984 230256
rect 146944 226636 146996 226642
rect 146944 226578 146996 226584
rect 52460 226568 52512 226574
rect 52460 226510 52512 226516
rect 62488 226568 62540 226574
rect 62488 226510 62540 226516
rect 79324 226568 79376 226574
rect 79324 226510 79376 226516
rect 43352 226500 43404 226506
rect 43352 226442 43404 226448
rect 37924 225616 37976 225622
rect 37924 225558 37976 225564
rect 43364 224890 43392 226442
rect 43102 224862 43392 224890
rect 52472 224890 52500 226510
rect 62120 226432 62172 226438
rect 62120 226374 62172 226380
rect 62132 224890 62160 226374
rect 52472 224862 52670 224890
rect 62132 224862 62330 224890
rect 41326 215248 41382 215257
rect 41326 215183 41382 215192
rect 37922 214024 37978 214033
rect 37922 213959 37978 213968
rect 36820 205556 36872 205562
rect 36820 205498 36872 205504
rect 36728 202700 36780 202706
rect 36728 202642 36780 202648
rect 36728 200388 36780 200394
rect 36728 200330 36780 200336
rect 36740 179314 36768 200330
rect 36820 200252 36872 200258
rect 36820 200194 36872 200200
rect 36728 179308 36780 179314
rect 36728 179250 36780 179256
rect 36832 176526 36860 200194
rect 37936 198014 37964 213959
rect 41340 205562 41368 215183
rect 62500 205714 62528 226510
rect 62764 226500 62816 226506
rect 62764 226442 62816 226448
rect 62422 205686 62528 205714
rect 41328 205556 41380 205562
rect 41328 205498 41380 205504
rect 42996 202774 43024 205020
rect 52762 205006 53144 205034
rect 53116 202842 53144 205006
rect 53104 202836 53156 202842
rect 53104 202778 53156 202784
rect 62776 202774 62804 226442
rect 64144 226432 64196 226438
rect 64144 226374 64196 226380
rect 64156 202842 64184 226374
rect 70308 226364 70360 226370
rect 70308 226306 70360 226312
rect 70320 224890 70348 226306
rect 70058 224862 70348 224890
rect 79336 224890 79364 226510
rect 90364 226500 90416 226506
rect 90364 226442 90416 226448
rect 106372 226500 106424 226506
rect 106372 226442 106424 226448
rect 116492 226500 116544 226506
rect 116492 226442 116544 226448
rect 133420 226500 133472 226506
rect 133420 226442 133472 226448
rect 89076 226432 89128 226438
rect 89076 226374 89128 226380
rect 89088 224890 89116 226374
rect 79336 224862 79718 224890
rect 89088 224862 89378 224890
rect 68926 214704 68982 214713
rect 68926 214639 68982 214648
rect 64878 214568 64934 214577
rect 64878 214503 64934 214512
rect 64892 205630 64920 214503
rect 64880 205624 64932 205630
rect 64880 205566 64932 205572
rect 68940 205494 68968 214639
rect 90376 209774 90404 226442
rect 90456 226432 90508 226438
rect 90456 226374 90508 226380
rect 89824 209746 90404 209774
rect 89824 205578 89852 209746
rect 89378 205550 89852 205578
rect 68928 205488 68980 205494
rect 68928 205430 68980 205436
rect 64144 202836 64196 202842
rect 64144 202778 64196 202784
rect 70044 202774 70072 205020
rect 79704 202774 79732 205020
rect 90468 202774 90496 226374
rect 90548 226364 90600 226370
rect 90548 226306 90600 226312
rect 90560 206310 90588 226306
rect 106384 224890 106412 226442
rect 115940 226432 115992 226438
rect 115940 226374 115992 226380
rect 115952 224890 115980 226374
rect 106384 224862 106674 224890
rect 115952 224862 116334 224890
rect 96724 224318 97014 224346
rect 95146 215248 95202 215257
rect 95146 215183 95202 215192
rect 91098 214568 91154 214577
rect 91098 214503 91154 214512
rect 90548 206304 90600 206310
rect 90548 206246 90600 206252
rect 91112 205562 91140 214503
rect 95160 205630 95188 215183
rect 95148 205624 95200 205630
rect 95148 205566 95200 205572
rect 91100 205556 91152 205562
rect 91100 205498 91152 205504
rect 96724 202774 96752 224318
rect 96804 206304 96856 206310
rect 96804 206246 96856 206252
rect 96816 205714 96844 206246
rect 96816 205686 97014 205714
rect 42984 202768 43036 202774
rect 42984 202710 43036 202716
rect 62764 202768 62816 202774
rect 62764 202710 62816 202716
rect 70032 202768 70084 202774
rect 70032 202710 70084 202716
rect 79692 202768 79744 202774
rect 79692 202710 79744 202716
rect 90456 202768 90508 202774
rect 90456 202710 90508 202716
rect 96712 202768 96764 202774
rect 96712 202710 96764 202716
rect 106660 202706 106688 205020
rect 116320 204898 116348 205020
rect 116504 204898 116532 226442
rect 116584 226432 116636 226438
rect 116584 226374 116636 226380
rect 116320 204870 116532 204898
rect 116596 202706 116624 226374
rect 133432 224890 133460 226442
rect 142988 226432 143040 226438
rect 142988 226374 143040 226380
rect 144276 226432 144328 226438
rect 144276 226374 144328 226380
rect 143000 224890 143028 226374
rect 144184 226364 144236 226370
rect 144184 226306 144236 226312
rect 133432 224862 133722 224890
rect 143000 224862 143382 224890
rect 122944 224318 124062 224346
rect 122746 215248 122802 215257
rect 122746 215183 122802 215192
rect 118698 214568 118754 214577
rect 118698 214503 118754 214512
rect 118712 205494 118740 214503
rect 122760 205562 122788 215183
rect 122748 205556 122800 205562
rect 122748 205498 122800 205504
rect 118700 205488 118752 205494
rect 118700 205430 118752 205436
rect 106648 202700 106700 202706
rect 106648 202642 106700 202648
rect 116584 202700 116636 202706
rect 116584 202642 116636 202648
rect 122944 202638 122972 224318
rect 144196 209774 144224 226306
rect 143736 209746 144224 209774
rect 143736 205578 143764 209746
rect 143382 205550 143764 205578
rect 124048 202774 124076 205020
rect 124036 202768 124088 202774
rect 124036 202710 124088 202716
rect 133708 202706 133736 205020
rect 144288 202706 144316 226374
rect 146298 214024 146354 214033
rect 146298 213959 146354 213968
rect 146312 205630 146340 213959
rect 146300 205624 146352 205630
rect 146300 205566 146352 205572
rect 133696 202700 133748 202706
rect 133696 202642 133748 202648
rect 144276 202700 144328 202706
rect 144276 202642 144328 202648
rect 122932 202632 122984 202638
rect 122932 202574 122984 202580
rect 52644 200388 52696 200394
rect 52644 200330 52696 200336
rect 43076 200320 43128 200326
rect 43076 200262 43128 200268
rect 37924 198008 37976 198014
rect 37924 197950 37976 197956
rect 43088 197948 43116 200262
rect 52656 197948 52684 200330
rect 62764 200320 62816 200326
rect 62764 200262 62816 200268
rect 90364 200320 90416 200326
rect 90364 200262 90416 200268
rect 106648 200320 106700 200326
rect 106648 200262 106700 200268
rect 116492 200320 116544 200326
rect 116492 200262 116544 200268
rect 133696 200320 133748 200326
rect 133696 200262 133748 200268
rect 144184 200320 144236 200326
rect 144184 200262 144236 200268
rect 62304 200252 62356 200258
rect 62304 200194 62356 200200
rect 62316 197948 62344 200194
rect 62488 200184 62540 200190
rect 62488 200126 62540 200132
rect 41326 188184 41382 188193
rect 41326 188119 41382 188128
rect 37922 186960 37978 186969
rect 37922 186895 37978 186904
rect 36820 176520 36872 176526
rect 36820 176462 36872 176468
rect 36636 176384 36688 176390
rect 36636 176326 36688 176332
rect 36728 172780 36780 172786
rect 36728 172722 36780 172728
rect 36636 169788 36688 169794
rect 36636 169730 36688 169736
rect 36544 148776 36596 148782
rect 36544 148718 36596 148724
rect 16028 146940 16080 146946
rect 16028 146882 16080 146888
rect 25688 146600 25740 146606
rect 25688 146542 25740 146548
rect 25700 143956 25728 146542
rect 35374 143534 35940 143562
rect 15212 143262 16054 143290
rect 13726 134192 13782 134201
rect 13726 134127 13782 134136
rect 13740 125594 13768 134127
rect 13728 125588 13780 125594
rect 13728 125530 13780 125536
rect 15212 122738 15240 143262
rect 35912 142154 35940 143534
rect 35912 142126 36584 142154
rect 35624 124840 35676 124846
rect 35374 124788 35624 124794
rect 35374 124782 35676 124788
rect 35374 124766 35664 124782
rect 16054 124086 16344 124114
rect 25714 124086 26096 124114
rect 15200 122732 15252 122738
rect 15200 122674 15252 122680
rect 16316 119406 16344 124086
rect 26068 122670 26096 124086
rect 26056 122664 26108 122670
rect 26056 122606 26108 122612
rect 16304 119400 16356 119406
rect 16304 119342 16356 119348
rect 25964 118992 26016 118998
rect 25964 118934 26016 118940
rect 25976 116906 26004 118934
rect 25714 116878 26004 116906
rect 15212 116334 16054 116362
rect 35374 116334 35664 116362
rect 13726 107264 13782 107273
rect 13726 107199 13782 107208
rect 13740 97986 13768 107199
rect 13728 97980 13780 97986
rect 13728 97922 13780 97928
rect 15212 95130 15240 116334
rect 35636 116142 35664 116334
rect 35624 116136 35676 116142
rect 35624 116078 35676 116084
rect 35374 97714 35664 97730
rect 35374 97708 35676 97714
rect 35374 97702 35624 97708
rect 35624 97650 35676 97656
rect 15304 97022 16054 97050
rect 15200 95124 15252 95130
rect 15200 95066 15252 95072
rect 15304 91798 15332 97022
rect 25700 95062 25728 97036
rect 25688 95056 25740 95062
rect 25688 94998 25740 95004
rect 36556 94926 36584 142126
rect 36648 122534 36676 169730
rect 36740 151706 36768 172722
rect 36820 172644 36872 172650
rect 36820 172586 36872 172592
rect 36728 151700 36780 151706
rect 36728 151642 36780 151648
rect 36832 148918 36860 172586
rect 37936 170406 37964 186895
rect 41340 179314 41368 188119
rect 41328 179308 41380 179314
rect 41328 179250 41380 179256
rect 62500 178786 62528 200126
rect 62422 178758 62528 178786
rect 42812 178078 43010 178106
rect 52762 178078 53144 178106
rect 42812 176594 42840 178078
rect 53116 176594 53144 178078
rect 62776 176662 62804 200262
rect 64144 200252 64196 200258
rect 64144 200194 64196 200200
rect 89352 200252 89404 200258
rect 89352 200194 89404 200200
rect 62764 176656 62816 176662
rect 62764 176598 62816 176604
rect 64156 176594 64184 200194
rect 79692 200184 79744 200190
rect 79692 200126 79744 200132
rect 79704 197948 79732 200126
rect 89364 197948 89392 200194
rect 69124 197254 70058 197282
rect 68926 187776 68982 187785
rect 68926 187711 68982 187720
rect 64878 187504 64934 187513
rect 64878 187439 64934 187448
rect 64892 179382 64920 187439
rect 64880 179376 64932 179382
rect 64880 179318 64932 179324
rect 68940 179246 68968 187711
rect 68928 179240 68980 179246
rect 68928 179182 68980 179188
rect 69124 176594 69152 197254
rect 90376 180794 90404 200262
rect 90456 200252 90508 200258
rect 90456 200194 90508 200200
rect 89824 180766 90404 180794
rect 89824 178786 89852 180766
rect 89378 178758 89852 178786
rect 69768 178078 70058 178106
rect 79718 178078 80008 178106
rect 69768 176662 69796 178078
rect 69756 176656 69808 176662
rect 69756 176598 69808 176604
rect 42800 176588 42852 176594
rect 42800 176530 42852 176536
rect 53104 176588 53156 176594
rect 53104 176530 53156 176536
rect 64144 176588 64196 176594
rect 64144 176530 64196 176536
rect 69112 176588 69164 176594
rect 69112 176530 69164 176536
rect 79980 176526 80008 178078
rect 90468 176526 90496 200194
rect 106660 197948 106688 200262
rect 116308 200252 116360 200258
rect 116308 200194 116360 200200
rect 116320 197948 116348 200194
rect 96724 197254 97014 197282
rect 95146 188184 95202 188193
rect 95146 188119 95202 188128
rect 91098 187504 91154 187513
rect 91098 187439 91154 187448
rect 91112 179314 91140 187439
rect 95160 179382 95188 188119
rect 95148 179376 95200 179382
rect 95148 179318 95200 179324
rect 91100 179308 91152 179314
rect 91100 179250 91152 179256
rect 96724 176662 96752 197254
rect 96816 178078 97014 178106
rect 106568 178078 106674 178106
rect 116228 178078 116334 178106
rect 96712 176656 96764 176662
rect 96712 176598 96764 176604
rect 96816 176594 96844 178078
rect 96804 176588 96856 176594
rect 96804 176530 96856 176536
rect 106568 176526 106596 178078
rect 116228 177970 116256 178078
rect 116504 177970 116532 200262
rect 116584 200252 116636 200258
rect 116584 200194 116636 200200
rect 116228 177942 116532 177970
rect 116596 176526 116624 200194
rect 133708 197948 133736 200262
rect 143356 200252 143408 200258
rect 143356 200194 143408 200200
rect 143368 197948 143396 200194
rect 122944 197254 124062 197282
rect 122746 188184 122802 188193
rect 122746 188119 122802 188128
rect 118698 187504 118754 187513
rect 118698 187439 118754 187448
rect 118712 179246 118740 187439
rect 122760 179314 122788 188119
rect 122748 179308 122800 179314
rect 122748 179250 122800 179256
rect 118700 179240 118752 179246
rect 118700 179182 118752 179188
rect 122944 176526 122972 197254
rect 144196 180794 144224 200262
rect 144276 200252 144328 200258
rect 144276 200194 144328 200200
rect 143736 180766 144224 180794
rect 143736 178786 143764 180766
rect 143382 178758 143764 178786
rect 123680 178078 124062 178106
rect 133722 178078 133828 178106
rect 123680 176594 123708 178078
rect 133800 176594 133828 178078
rect 144288 176594 144316 200194
rect 146298 186960 146354 186969
rect 146298 186895 146354 186904
rect 146312 179382 146340 186895
rect 146300 179376 146352 179382
rect 146300 179318 146352 179324
rect 146956 176662 146984 226578
rect 148336 202774 148364 254186
rect 232044 254176 232096 254182
rect 232044 254118 232096 254124
rect 251824 254176 251876 254182
rect 251824 254118 251876 254124
rect 475016 254176 475068 254182
rect 475016 254118 475068 254124
rect 494704 254176 494756 254182
rect 494704 254118 494756 254124
rect 170496 254108 170548 254114
rect 170496 254050 170548 254056
rect 187700 254108 187752 254114
rect 187700 254050 187752 254056
rect 197452 254108 197504 254114
rect 197452 254050 197504 254056
rect 214656 254108 214708 254114
rect 214656 254050 214708 254056
rect 224500 254108 224552 254114
rect 224500 254050 224552 254056
rect 170312 254040 170364 254046
rect 170312 253982 170364 253988
rect 160652 253972 160704 253978
rect 160652 253914 160704 253920
rect 160664 251940 160692 253914
rect 170324 251940 170352 253982
rect 148968 251252 149020 251258
rect 148968 251194 149020 251200
rect 150544 251246 151018 251274
rect 148980 242321 149008 251194
rect 148966 242312 149022 242321
rect 148966 242247 149022 242256
rect 150544 230314 150572 251246
rect 150728 232070 151018 232098
rect 160572 232070 160678 232098
rect 170232 232070 170338 232098
rect 150728 230382 150756 232070
rect 150716 230376 150768 230382
rect 150716 230318 150768 230324
rect 150532 230308 150584 230314
rect 150532 230250 150584 230256
rect 160572 230246 160600 232070
rect 170232 231962 170260 232070
rect 170508 231962 170536 254050
rect 178040 254040 178092 254046
rect 178040 253982 178092 253988
rect 171784 253972 171836 253978
rect 171784 253914 171836 253920
rect 170232 231934 170536 231962
rect 171796 230246 171824 253914
rect 178052 251940 178080 253982
rect 187712 251940 187740 254050
rect 197360 253972 197412 253978
rect 197360 253914 197412 253920
rect 197372 251940 197400 253914
rect 172520 251320 172572 251326
rect 172520 251262 172572 251268
rect 172532 241641 172560 251262
rect 172518 241632 172574 241641
rect 172518 241567 172574 241576
rect 176566 241632 176622 241641
rect 176566 241567 176622 241576
rect 176580 233238 176608 241567
rect 176568 233232 176620 233238
rect 176568 233174 176620 233180
rect 197464 232778 197492 254050
rect 200764 254040 200816 254046
rect 200764 253982 200816 253988
rect 199384 253972 199436 253978
rect 199384 253914 199436 253920
rect 197386 232750 197492 232778
rect 178066 232070 178172 232098
rect 187726 232070 188016 232098
rect 178144 230314 178172 232070
rect 187988 230314 188016 232070
rect 199396 230314 199424 253914
rect 200120 251252 200172 251258
rect 200120 251194 200172 251200
rect 200132 241641 200160 251194
rect 200118 241632 200174 241641
rect 200118 241567 200174 241576
rect 200776 230450 200804 253982
rect 214668 251940 214696 254050
rect 224316 253972 224368 253978
rect 224316 253914 224368 253920
rect 224328 251940 224356 253914
rect 202788 251252 202840 251258
rect 202788 251194 202840 251200
rect 204364 251246 205022 251274
rect 202800 242321 202828 251194
rect 202786 242312 202842 242321
rect 202786 242247 202842 242256
rect 200764 230444 200816 230450
rect 200764 230386 200816 230392
rect 204364 230314 204392 251246
rect 224512 232778 224540 254050
rect 225604 253972 225656 253978
rect 225604 253914 225656 253920
rect 224342 232750 224540 232778
rect 204640 232070 205022 232098
rect 214682 232070 215064 232098
rect 204640 230450 204668 232070
rect 204628 230444 204680 230450
rect 204628 230386 204680 230392
rect 178132 230308 178184 230314
rect 178132 230250 178184 230256
rect 187976 230308 188028 230314
rect 187976 230250 188028 230256
rect 199384 230308 199436 230314
rect 199384 230250 199436 230256
rect 204352 230308 204404 230314
rect 204352 230250 204404 230256
rect 215036 230246 215064 232070
rect 225616 230246 225644 253914
rect 232056 251940 232084 254118
rect 241704 254108 241756 254114
rect 241704 254050 241756 254056
rect 241716 251940 241744 254050
rect 251456 254040 251508 254046
rect 251456 253982 251508 253988
rect 251364 253972 251416 253978
rect 251364 253914 251416 253920
rect 251376 251940 251404 253914
rect 230388 251320 230440 251326
rect 230388 251262 230440 251268
rect 230400 242321 230428 251262
rect 230386 242312 230442 242321
rect 230386 242247 230442 242256
rect 226338 241632 226394 241641
rect 226338 241567 226394 241576
rect 226352 233238 226380 241567
rect 226340 233232 226392 233238
rect 226340 233174 226392 233180
rect 251468 232778 251496 253982
rect 251390 232750 251496 232778
rect 231872 232070 232070 232098
rect 241730 232070 242112 232098
rect 231872 230314 231900 232070
rect 242084 230314 242112 232070
rect 251836 230450 251864 254118
rect 413468 254108 413520 254114
rect 413468 254050 413520 254056
rect 430672 254108 430724 254114
rect 430672 254050 430724 254056
rect 440516 254108 440568 254114
rect 440516 254050 440568 254056
rect 457628 254108 457680 254114
rect 457628 254050 457680 254056
rect 468576 254108 468628 254114
rect 468576 254050 468628 254056
rect 268660 254040 268712 254046
rect 268660 253982 268712 253988
rect 279424 254040 279476 254046
rect 279424 253982 279476 253988
rect 295708 254040 295760 254046
rect 295708 253982 295760 253988
rect 305460 254040 305512 254046
rect 305460 253982 305512 253988
rect 322664 254040 322716 254046
rect 322664 253982 322716 253988
rect 334624 254040 334676 254046
rect 334624 253982 334676 253988
rect 349712 254040 349764 254046
rect 349712 253982 349764 253988
rect 359464 254040 359516 254046
rect 359464 253982 359516 253988
rect 376668 254040 376720 254046
rect 376668 253982 376720 253988
rect 386512 254040 386564 254046
rect 386512 253982 386564 253988
rect 403624 254040 403676 254046
rect 403624 253982 403676 253988
rect 253204 253972 253256 253978
rect 253204 253914 253256 253920
rect 251824 230444 251876 230450
rect 251824 230386 251876 230392
rect 253216 230314 253244 253914
rect 268672 251940 268700 253982
rect 278320 253972 278372 253978
rect 278320 253914 278372 253920
rect 278332 251940 278360 253914
rect 253940 251252 253992 251258
rect 253940 251194 253992 251200
rect 258184 251246 259026 251274
rect 253952 242185 253980 251194
rect 253938 242176 253994 242185
rect 253938 242111 253994 242120
rect 256606 242176 256662 242185
rect 256606 242111 256662 242120
rect 256620 233238 256648 242111
rect 256608 233232 256660 233238
rect 256608 233174 256660 233180
rect 257988 231872 258040 231878
rect 257988 231814 258040 231820
rect 258000 230450 258028 231814
rect 257988 230444 258040 230450
rect 257988 230386 258040 230392
rect 258184 230314 258212 251246
rect 279436 238754 279464 253982
rect 279516 253972 279568 253978
rect 279516 253914 279568 253920
rect 278792 238726 279464 238754
rect 278792 232778 278820 238726
rect 278346 232750 278820 232778
rect 258736 232070 259026 232098
rect 268686 232070 268976 232098
rect 258736 231878 258764 232070
rect 258724 231872 258776 231878
rect 258724 231814 258776 231820
rect 231860 230308 231912 230314
rect 231860 230250 231912 230256
rect 242072 230308 242124 230314
rect 242072 230250 242124 230256
rect 253204 230308 253256 230314
rect 253204 230250 253256 230256
rect 258172 230308 258224 230314
rect 258172 230250 258224 230256
rect 268948 230246 268976 232070
rect 279528 230246 279556 253914
rect 285784 252062 286088 252090
rect 280160 251320 280212 251326
rect 280160 251262 280212 251268
rect 280172 241641 280200 251262
rect 284208 251252 284260 251258
rect 284208 251194 284260 251200
rect 284220 242865 284248 251194
rect 284206 242856 284262 242865
rect 284206 242791 284262 242800
rect 280158 241632 280214 241641
rect 280158 241567 280214 241576
rect 285784 230246 285812 252062
rect 286060 251940 286088 252062
rect 295720 251940 295748 253982
rect 305368 253972 305420 253978
rect 305368 253914 305420 253920
rect 305380 251940 305408 253914
rect 305472 232778 305500 253982
rect 307024 253972 307076 253978
rect 307024 253914 307076 253920
rect 305394 232750 305500 232778
rect 286074 232070 286180 232098
rect 295734 232070 296024 232098
rect 286152 230314 286180 232070
rect 286140 230308 286192 230314
rect 286140 230250 286192 230256
rect 295996 230246 296024 232070
rect 307036 230246 307064 253914
rect 322676 251940 322704 253982
rect 332324 253972 332376 253978
rect 332324 253914 332376 253920
rect 333244 253972 333296 253978
rect 333244 253914 333296 253920
rect 332336 251940 332364 253914
rect 311808 251320 311860 251326
rect 311808 251262 311860 251268
rect 311820 242321 311848 251262
rect 312004 251246 313030 251274
rect 311806 242312 311862 242321
rect 311806 242247 311862 242256
rect 307758 241632 307814 241641
rect 307758 241567 307814 241576
rect 307772 233238 307800 241567
rect 307760 233232 307812 233238
rect 307760 233174 307812 233180
rect 312004 230246 312032 251246
rect 332508 233232 332560 233238
rect 332508 233174 332560 233180
rect 332520 232778 332548 233174
rect 332350 232750 332548 232778
rect 312648 232070 313030 232098
rect 322690 232070 322888 232098
rect 312648 230314 312676 232070
rect 312636 230308 312688 230314
rect 312636 230250 312688 230256
rect 322860 230246 322888 232070
rect 333256 230246 333284 253914
rect 334636 233238 334664 253982
rect 339604 252062 340092 252090
rect 335360 251252 335412 251258
rect 335360 251194 335412 251200
rect 335372 241641 335400 251194
rect 338026 242176 338082 242185
rect 338026 242111 338082 242120
rect 335358 241632 335414 241641
rect 335358 241567 335414 241576
rect 338040 233238 338068 242111
rect 334624 233232 334676 233238
rect 334624 233174 334676 233180
rect 338028 233232 338080 233238
rect 338028 233174 338080 233180
rect 339604 230246 339632 252062
rect 340064 251940 340092 252062
rect 349724 251940 349752 253982
rect 359372 253972 359424 253978
rect 359372 253914 359424 253920
rect 359384 251940 359412 253914
rect 359476 232778 359504 253982
rect 359556 253972 359608 253978
rect 359556 253914 359608 253920
rect 359398 232750 359504 232778
rect 340078 232070 340184 232098
rect 349738 232070 350120 232098
rect 340156 230314 340184 232070
rect 340144 230308 340196 230314
rect 340144 230250 340196 230256
rect 350092 230246 350120 232070
rect 359568 230246 359596 253914
rect 376680 251940 376708 253982
rect 386328 253972 386380 253978
rect 386328 253914 386380 253920
rect 386340 251940 386368 253914
rect 361580 251320 361632 251326
rect 361580 251262 361632 251268
rect 361592 242185 361620 251262
rect 365628 251252 365680 251258
rect 365628 251194 365680 251200
rect 365824 251246 367034 251274
rect 365640 242321 365668 251194
rect 365626 242312 365682 242321
rect 365626 242247 365682 242256
rect 361578 242176 361634 242185
rect 361578 242111 361634 242120
rect 365824 230246 365852 251246
rect 386524 232778 386552 253982
rect 387064 253972 387116 253978
rect 387064 253914 387116 253920
rect 386354 232750 386552 232778
rect 366744 232070 367034 232098
rect 376588 232070 376694 232098
rect 366744 230314 366772 232070
rect 366732 230308 366784 230314
rect 366732 230250 366784 230256
rect 376588 230246 376616 232070
rect 387076 230246 387104 253914
rect 403636 251940 403664 253982
rect 413284 253972 413336 253978
rect 413284 253914 413336 253920
rect 413296 251940 413324 253914
rect 393424 251246 393990 251274
rect 391846 241904 391902 241913
rect 391846 241839 391902 241848
rect 389178 241632 389234 241641
rect 389178 241567 389234 241576
rect 389192 233238 389220 241567
rect 391860 233238 391888 241839
rect 389180 233232 389232 233238
rect 389180 233174 389232 233180
rect 391848 233232 391900 233238
rect 391848 233174 391900 233180
rect 393424 230246 393452 251246
rect 413480 232778 413508 254050
rect 421012 254040 421064 254046
rect 421012 253982 421064 253988
rect 414664 253972 414716 253978
rect 414664 253914 414716 253920
rect 413402 232750 413508 232778
rect 393608 232070 393990 232098
rect 403742 232070 404032 232098
rect 393608 230314 393636 232070
rect 393596 230308 393648 230314
rect 393596 230250 393648 230256
rect 404004 230246 404032 232070
rect 414676 230246 414704 253914
rect 421024 251940 421052 253982
rect 430684 251940 430712 254050
rect 440332 253972 440384 253978
rect 440332 253914 440384 253920
rect 440344 251940 440372 253914
rect 415400 251252 415452 251258
rect 415400 251194 415452 251200
rect 419448 251252 419500 251258
rect 419448 251194 419500 251200
rect 415412 241641 415440 251194
rect 419460 242321 419488 251194
rect 419446 242312 419502 242321
rect 419446 242247 419502 242256
rect 415398 241632 415454 241641
rect 415398 241567 415454 241576
rect 440528 232778 440556 254050
rect 443644 254040 443696 254046
rect 443644 253982 443696 253988
rect 442264 253972 442316 253978
rect 442264 253914 442316 253920
rect 440358 232750 440556 232778
rect 420932 232070 421038 232098
rect 430698 232070 431080 232098
rect 420932 230314 420960 232070
rect 431052 230314 431080 232070
rect 442276 230314 442304 253914
rect 442998 241632 443054 241641
rect 442998 241567 443054 241576
rect 443012 233238 443040 241567
rect 443000 233232 443052 233238
rect 443000 233174 443052 233180
rect 443656 230450 443684 253982
rect 457640 251940 457668 254050
rect 467288 253972 467340 253978
rect 467288 253914 467340 253920
rect 468484 253972 468536 253978
rect 468484 253914 468536 253920
rect 467300 251940 467328 253914
rect 447244 251246 447994 251274
rect 445666 242176 445722 242185
rect 445666 242111 445722 242120
rect 445680 233238 445708 242111
rect 445668 233232 445720 233238
rect 445668 233174 445720 233180
rect 443644 230444 443696 230450
rect 443644 230386 443696 230392
rect 447244 230314 447272 251246
rect 467656 233164 467708 233170
rect 467656 233106 467708 233112
rect 467668 232778 467696 233106
rect 467406 232750 467696 232778
rect 447704 232070 447994 232098
rect 457746 232070 458128 232098
rect 447704 230450 447732 232070
rect 447692 230444 447744 230450
rect 447692 230386 447744 230392
rect 420920 230308 420972 230314
rect 420920 230250 420972 230256
rect 431040 230308 431092 230314
rect 431040 230250 431092 230256
rect 442264 230308 442316 230314
rect 442264 230250 442316 230256
rect 447232 230308 447284 230314
rect 447232 230250 447284 230256
rect 458100 230246 458128 232070
rect 468496 230246 468524 253914
rect 468588 233170 468616 254050
rect 475028 251940 475056 254118
rect 484676 254108 484728 254114
rect 484676 254050 484728 254056
rect 484688 251940 484716 254050
rect 494520 254040 494572 254046
rect 494520 253982 494572 253988
rect 494336 253972 494388 253978
rect 494336 253914 494388 253920
rect 494348 251940 494376 253914
rect 469220 251252 469272 251258
rect 469220 251194 469272 251200
rect 473268 251252 473320 251258
rect 473268 251194 473320 251200
rect 469232 242185 469260 251194
rect 473280 242865 473308 251194
rect 473266 242856 473322 242865
rect 473266 242791 473322 242800
rect 469218 242176 469274 242185
rect 469218 242111 469274 242120
rect 468576 233164 468628 233170
rect 468576 233106 468628 233112
rect 494532 232778 494560 253982
rect 494362 232750 494560 232778
rect 474752 232070 475042 232098
rect 484702 232070 484992 232098
rect 474752 230314 474780 232070
rect 484964 230314 484992 232070
rect 494716 231878 494744 254118
rect 511632 254040 511684 254046
rect 511632 253982 511684 253988
rect 522396 254040 522448 254046
rect 522396 253982 522448 253988
rect 496084 253972 496136 253978
rect 496084 253914 496136 253920
rect 494704 231872 494756 231878
rect 494704 231814 494756 231820
rect 496096 230314 496124 253914
rect 511644 251940 511672 253982
rect 521292 253972 521344 253978
rect 521292 253914 521344 253920
rect 522304 253972 522356 253978
rect 522304 253914 522356 253920
rect 521304 251940 521332 253914
rect 500868 251320 500920 251326
rect 500868 251262 500920 251268
rect 500880 242321 500908 251262
rect 501064 251246 501998 251274
rect 500866 242312 500922 242321
rect 500866 242247 500922 242256
rect 496818 241632 496874 241641
rect 496818 241567 496874 241576
rect 496832 233238 496860 241567
rect 496820 233232 496872 233238
rect 496820 233174 496872 233180
rect 501064 230314 501092 251246
rect 521752 235408 521804 235414
rect 521752 235350 521804 235356
rect 521764 232778 521792 235350
rect 521410 232750 521792 232778
rect 501616 232070 501998 232098
rect 511750 232070 511948 232098
rect 501616 231878 501644 232070
rect 501604 231872 501656 231878
rect 501604 231814 501656 231820
rect 474740 230308 474792 230314
rect 474740 230250 474792 230256
rect 484952 230308 485004 230314
rect 484952 230250 485004 230256
rect 496084 230308 496136 230314
rect 496084 230250 496136 230256
rect 501052 230308 501104 230314
rect 501052 230250 501104 230256
rect 511920 230246 511948 232070
rect 522316 230246 522344 253914
rect 522408 235414 522436 253982
rect 529032 251940 529060 254526
rect 538680 254040 538732 254046
rect 538680 253982 538732 253988
rect 538692 251940 538720 253982
rect 548340 253972 548392 253978
rect 548340 253914 548392 253920
rect 548352 251940 548380 253914
rect 526444 251864 526496 251870
rect 526444 251806 526496 251812
rect 523040 251252 523092 251258
rect 523040 251194 523092 251200
rect 523052 241641 523080 251194
rect 526456 242321 526484 251806
rect 550640 251320 550692 251326
rect 550640 251262 550692 251268
rect 526442 242312 526498 242321
rect 526442 242247 526498 242256
rect 550652 241641 550680 251262
rect 523038 241632 523094 241641
rect 523038 241567 523094 241576
rect 550638 241632 550694 241641
rect 550638 241567 550694 241576
rect 522396 235408 522448 235414
rect 522396 235350 522448 235356
rect 528664 232070 529046 232098
rect 538416 232070 538706 232098
rect 547984 232070 548366 232098
rect 528664 230314 528692 232070
rect 528652 230308 528704 230314
rect 528652 230250 528704 230256
rect 160560 230240 160612 230246
rect 160560 230182 160612 230188
rect 171784 230240 171836 230246
rect 171784 230182 171836 230188
rect 215024 230240 215076 230246
rect 215024 230182 215076 230188
rect 225604 230240 225656 230246
rect 225604 230182 225656 230188
rect 268936 230240 268988 230246
rect 268936 230182 268988 230188
rect 279516 230240 279568 230246
rect 279516 230182 279568 230188
rect 285772 230240 285824 230246
rect 285772 230182 285824 230188
rect 295984 230240 296036 230246
rect 295984 230182 296036 230188
rect 307024 230240 307076 230246
rect 307024 230182 307076 230188
rect 311992 230240 312044 230246
rect 311992 230182 312044 230188
rect 322848 230240 322900 230246
rect 322848 230182 322900 230188
rect 333244 230240 333296 230246
rect 333244 230182 333296 230188
rect 339592 230240 339644 230246
rect 339592 230182 339644 230188
rect 350080 230240 350132 230246
rect 350080 230182 350132 230188
rect 359556 230240 359608 230246
rect 359556 230182 359608 230188
rect 365812 230240 365864 230246
rect 365812 230182 365864 230188
rect 376576 230240 376628 230246
rect 376576 230182 376628 230188
rect 387064 230240 387116 230246
rect 387064 230182 387116 230188
rect 393412 230240 393464 230246
rect 393412 230182 393464 230188
rect 403992 230240 404044 230246
rect 403992 230182 404044 230188
rect 414664 230240 414716 230246
rect 414664 230182 414716 230188
rect 458088 230240 458140 230246
rect 458088 230182 458140 230188
rect 468484 230240 468536 230246
rect 468484 230182 468536 230188
rect 511908 230240 511960 230246
rect 511908 230182 511960 230188
rect 522304 230240 522356 230246
rect 522304 230182 522356 230188
rect 538416 230178 538444 232070
rect 547984 230382 548012 232070
rect 547972 230376 548024 230382
rect 547972 230318 548024 230324
rect 538404 230172 538456 230178
rect 538404 230114 538456 230120
rect 528744 227044 528796 227050
rect 528744 226986 528796 226992
rect 259368 226568 259420 226574
rect 259368 226510 259420 226516
rect 279608 226568 279660 226574
rect 279608 226510 279660 226516
rect 448336 226568 448388 226574
rect 448336 226510 448388 226516
rect 468668 226568 468720 226574
rect 468668 226510 468720 226516
rect 170496 226500 170548 226506
rect 170496 226442 170548 226448
rect 187792 226500 187844 226506
rect 187792 226442 187844 226448
rect 197544 226500 197596 226506
rect 197544 226442 197596 226448
rect 214380 226500 214432 226506
rect 214380 226442 214432 226448
rect 224500 226500 224552 226506
rect 224500 226442 224552 226448
rect 241520 226500 241572 226506
rect 241520 226442 241572 226448
rect 251456 226500 251508 226506
rect 251456 226442 251508 226448
rect 170036 226432 170088 226438
rect 170036 226374 170088 226380
rect 160284 226364 160336 226370
rect 160284 226306 160336 226312
rect 160296 224890 160324 226306
rect 170048 224890 170076 226374
rect 160296 224862 160678 224890
rect 170048 224862 170338 224890
rect 150544 224318 151018 224346
rect 148966 215248 149022 215257
rect 148966 215183 149022 215192
rect 148980 205630 149008 215183
rect 148968 205624 149020 205630
rect 148968 205566 149020 205572
rect 148324 202768 148376 202774
rect 148324 202710 148376 202716
rect 150544 202706 150572 224318
rect 150532 202700 150584 202706
rect 150532 202642 150584 202648
rect 151004 202638 151032 205020
rect 160664 202638 160692 205020
rect 170324 204898 170352 205020
rect 170508 204898 170536 226442
rect 178408 226432 178460 226438
rect 178408 226374 178460 226380
rect 171784 226364 171836 226370
rect 171784 226306 171836 226312
rect 170324 204870 170536 204898
rect 171796 202638 171824 226306
rect 178420 224890 178448 226374
rect 187804 224890 187832 226442
rect 197452 226364 197504 226370
rect 197452 226306 197504 226312
rect 197464 224890 197492 226306
rect 178066 224862 178448 224890
rect 187726 224862 187832 224890
rect 197386 224862 197492 224890
rect 197556 219434 197584 226442
rect 200764 226432 200816 226438
rect 200764 226374 200816 226380
rect 199384 226364 199436 226370
rect 199384 226306 199436 226312
rect 197464 219406 197584 219434
rect 176566 214704 176622 214713
rect 176566 214639 176622 214648
rect 172518 214568 172574 214577
rect 172518 214503 172574 214512
rect 172532 205562 172560 214503
rect 176580 205562 176608 214639
rect 197464 205714 197492 219406
rect 197386 205686 197492 205714
rect 172520 205556 172572 205562
rect 172520 205498 172572 205504
rect 176568 205556 176620 205562
rect 176568 205498 176620 205504
rect 178052 202706 178080 205020
rect 187712 202706 187740 205020
rect 199396 202706 199424 226306
rect 200118 214568 200174 214577
rect 200118 214503 200174 214512
rect 200132 205630 200160 214503
rect 200120 205624 200172 205630
rect 200120 205566 200172 205572
rect 200776 205494 200804 226374
rect 214392 224890 214420 226442
rect 223948 226364 224000 226370
rect 223948 226306 224000 226312
rect 223960 224890 223988 226306
rect 214392 224862 214682 224890
rect 223960 224862 224342 224890
rect 204364 224318 205022 224346
rect 202786 215248 202842 215257
rect 202786 215183 202842 215192
rect 202800 205630 202828 215183
rect 202788 205624 202840 205630
rect 202788 205566 202840 205572
rect 200764 205488 200816 205494
rect 200764 205430 200816 205436
rect 204364 202706 204392 224318
rect 224512 205714 224540 226442
rect 232320 226432 232372 226438
rect 232320 226374 232372 226380
rect 225604 226364 225656 226370
rect 225604 226306 225656 226312
rect 224342 205686 224540 205714
rect 204628 205488 204680 205494
rect 204680 205436 205022 205442
rect 204628 205430 205022 205436
rect 204640 205414 205022 205430
rect 178040 202700 178092 202706
rect 178040 202642 178092 202648
rect 187700 202700 187752 202706
rect 187700 202642 187752 202648
rect 199384 202700 199436 202706
rect 199384 202642 199436 202648
rect 204352 202700 204404 202706
rect 204352 202642 204404 202648
rect 214668 202638 214696 205020
rect 225616 202638 225644 226306
rect 232332 224890 232360 226374
rect 232070 224862 232360 224890
rect 241532 224890 241560 226442
rect 251180 226364 251232 226370
rect 251180 226306 251232 226312
rect 251192 224890 251220 226306
rect 241532 224862 241730 224890
rect 251192 224862 251390 224890
rect 230386 215248 230442 215257
rect 230386 215183 230442 215192
rect 226338 214568 226394 214577
rect 226338 214503 226394 214512
rect 226352 205562 226380 214503
rect 230400 205562 230428 215183
rect 251468 205714 251496 226442
rect 251824 226432 251876 226438
rect 251824 226374 251876 226380
rect 251390 205686 251496 205714
rect 226340 205556 226392 205562
rect 226340 205498 226392 205504
rect 230388 205556 230440 205562
rect 230388 205498 230440 205504
rect 232056 202706 232084 205020
rect 241716 202706 241744 205020
rect 251836 202842 251864 226374
rect 253204 226364 253256 226370
rect 253204 226306 253256 226312
rect 251824 202836 251876 202842
rect 251824 202778 251876 202784
rect 253216 202706 253244 226306
rect 259380 224890 259408 226510
rect 268292 226500 268344 226506
rect 268292 226442 268344 226448
rect 259026 224862 259408 224890
rect 268304 224890 268332 226442
rect 279424 226432 279476 226438
rect 279424 226374 279476 226380
rect 278044 226364 278096 226370
rect 278044 226306 278096 226312
rect 278056 224890 278084 226306
rect 268304 224862 268686 224890
rect 278056 224862 278346 224890
rect 256606 215248 256662 215257
rect 256606 215183 256662 215192
rect 253938 214024 253994 214033
rect 253938 213959 253994 213968
rect 253952 205630 253980 213959
rect 256620 205630 256648 215183
rect 279436 209774 279464 226374
rect 279516 226364 279568 226370
rect 279516 226306 279568 226312
rect 278792 209746 279464 209774
rect 253940 205624 253992 205630
rect 253940 205566 253992 205572
rect 256608 205624 256660 205630
rect 278792 205578 278820 209746
rect 256608 205566 256660 205572
rect 278346 205550 278820 205578
rect 259012 202842 259040 205020
rect 259000 202836 259052 202842
rect 259000 202778 259052 202784
rect 268672 202706 268700 205020
rect 279528 202706 279556 226306
rect 279620 205698 279648 226510
rect 413468 226500 413520 226506
rect 413468 226442 413520 226448
rect 430580 226500 430632 226506
rect 430580 226442 430632 226448
rect 440516 226500 440568 226506
rect 440516 226442 440568 226448
rect 295800 226432 295852 226438
rect 295800 226374 295852 226380
rect 305644 226432 305696 226438
rect 305644 226374 305696 226380
rect 322388 226432 322440 226438
rect 322388 226374 322440 226380
rect 336004 226432 336056 226438
rect 336004 226374 336056 226380
rect 349804 226432 349856 226438
rect 349804 226374 349856 226380
rect 359556 226432 359608 226438
rect 359556 226374 359608 226380
rect 376300 226432 376352 226438
rect 376300 226374 376352 226380
rect 386512 226432 386564 226438
rect 386512 226374 386564 226380
rect 403348 226432 403400 226438
rect 403348 226374 403400 226380
rect 295812 224890 295840 226374
rect 305552 226364 305604 226370
rect 305552 226306 305604 226312
rect 305564 224890 305592 226306
rect 295734 224862 295840 224890
rect 305394 224862 305592 224890
rect 286074 224330 286180 224346
rect 285772 224324 285824 224330
rect 286074 224324 286192 224330
rect 286074 224318 286140 224324
rect 285772 224266 285824 224272
rect 286140 224266 286192 224272
rect 284206 214704 284262 214713
rect 284206 214639 284262 214648
rect 280158 214568 280214 214577
rect 280158 214503 280214 214512
rect 279608 205692 279660 205698
rect 279608 205634 279660 205640
rect 280172 205562 280200 214503
rect 284220 205562 284248 214639
rect 280160 205556 280212 205562
rect 280160 205498 280212 205504
rect 284208 205556 284260 205562
rect 284208 205498 284260 205504
rect 285784 202706 285812 224266
rect 305656 219434 305684 226374
rect 307024 226364 307076 226370
rect 307024 226306 307076 226312
rect 305472 219406 305684 219434
rect 305472 205714 305500 219406
rect 286140 205692 286192 205698
rect 305394 205686 305500 205714
rect 286140 205634 286192 205640
rect 286152 205578 286180 205634
rect 286074 205550 286180 205578
rect 232044 202700 232096 202706
rect 232044 202642 232096 202648
rect 241704 202700 241756 202706
rect 241704 202642 241756 202648
rect 253204 202700 253256 202706
rect 253204 202642 253256 202648
rect 268660 202700 268712 202706
rect 268660 202642 268712 202648
rect 279516 202700 279568 202706
rect 279516 202642 279568 202648
rect 285772 202700 285824 202706
rect 285772 202642 285824 202648
rect 295720 202638 295748 205020
rect 307036 202638 307064 226306
rect 322400 224890 322428 226374
rect 331956 226364 332008 226370
rect 331956 226306 332008 226312
rect 333244 226364 333296 226370
rect 333244 226306 333296 226312
rect 331968 224890 331996 226306
rect 322400 224862 322690 224890
rect 331968 224862 332350 224890
rect 312004 224318 313030 224346
rect 311806 215248 311862 215257
rect 311806 215183 311862 215192
rect 307758 214568 307814 214577
rect 307758 214503 307814 214512
rect 307772 205630 307800 214503
rect 307760 205624 307812 205630
rect 307760 205566 307812 205572
rect 311820 205494 311848 215183
rect 311808 205488 311860 205494
rect 311808 205430 311860 205436
rect 312004 202638 312032 224318
rect 313016 202706 313044 205020
rect 313004 202700 313056 202706
rect 313004 202642 313056 202648
rect 322676 202638 322704 205020
rect 332336 202842 332364 205020
rect 332324 202836 332376 202842
rect 332324 202778 332376 202784
rect 333256 202638 333284 226306
rect 335358 214568 335414 214577
rect 335358 214503 335414 214512
rect 335372 205562 335400 214503
rect 335360 205556 335412 205562
rect 335360 205498 335412 205504
rect 336016 202842 336044 226374
rect 349816 224890 349844 226374
rect 359464 226364 359516 226370
rect 359464 226306 359516 226312
rect 359476 224890 359504 226306
rect 349738 224862 349844 224890
rect 359398 224862 359504 224890
rect 340078 224330 340184 224346
rect 339592 224324 339644 224330
rect 340078 224324 340196 224330
rect 340078 224318 340144 224324
rect 339592 224266 339644 224272
rect 340144 224266 340196 224272
rect 338026 215248 338082 215257
rect 338026 215183 338082 215192
rect 338040 205630 338068 215183
rect 338028 205624 338080 205630
rect 338028 205566 338080 205572
rect 336004 202836 336056 202842
rect 336004 202778 336056 202784
rect 339604 202638 339632 224266
rect 359568 223122 359596 226374
rect 359740 226364 359792 226370
rect 359740 226306 359792 226312
rect 359476 223094 359596 223122
rect 359476 205714 359504 223094
rect 359752 222850 359780 226306
rect 376312 224890 376340 226374
rect 386052 226364 386104 226370
rect 386052 226306 386104 226312
rect 386064 224890 386092 226306
rect 376312 224862 376694 224890
rect 386064 224862 386354 224890
rect 359398 205686 359504 205714
rect 359568 222822 359780 222850
rect 365824 224318 367034 224346
rect 340064 202706 340092 205020
rect 340052 202700 340104 202706
rect 340052 202642 340104 202648
rect 349724 202638 349752 205020
rect 359568 202638 359596 222822
rect 365626 215248 365682 215257
rect 365626 215183 365682 215192
rect 361578 214024 361634 214033
rect 361578 213959 361634 213968
rect 361592 205494 361620 213959
rect 365640 205562 365668 215183
rect 365628 205556 365680 205562
rect 365628 205498 365680 205504
rect 361580 205488 361632 205494
rect 361580 205430 361632 205436
rect 365824 202638 365852 224318
rect 386524 205714 386552 226374
rect 387064 226364 387116 226370
rect 387064 226306 387116 226312
rect 386354 205686 386552 205714
rect 367020 202706 367048 205020
rect 367008 202700 367060 202706
rect 367008 202642 367060 202648
rect 376680 202638 376708 205020
rect 387076 202638 387104 226306
rect 403360 224890 403388 226374
rect 412916 226364 412968 226370
rect 412916 226306 412968 226312
rect 412928 224890 412956 226306
rect 403360 224862 403650 224890
rect 412928 224862 413310 224890
rect 393424 224318 393990 224346
rect 391846 215248 391902 215257
rect 391846 215183 391902 215192
rect 389178 214568 389234 214577
rect 389178 214503 389234 214512
rect 389192 205630 389220 214503
rect 391860 205630 391888 215183
rect 389180 205624 389232 205630
rect 389180 205566 389232 205572
rect 391848 205624 391900 205630
rect 391848 205566 391900 205572
rect 393424 202638 393452 224318
rect 413480 205714 413508 226442
rect 421288 226432 421340 226438
rect 421288 226374 421340 226380
rect 414664 226364 414716 226370
rect 414664 226306 414716 226312
rect 413402 205686 413508 205714
rect 393608 205006 393990 205034
rect 393608 202706 393636 205006
rect 393596 202700 393648 202706
rect 393596 202642 393648 202648
rect 403728 202638 403756 205020
rect 414676 202638 414704 226306
rect 421300 224890 421328 226374
rect 421038 224862 421328 224890
rect 430592 224890 430620 226442
rect 440240 226364 440292 226370
rect 440240 226306 440292 226312
rect 440252 224890 440280 226306
rect 430592 224862 430698 224890
rect 440252 224862 440358 224890
rect 419446 215248 419502 215257
rect 419446 215183 419502 215192
rect 415398 214568 415454 214577
rect 415398 214503 415454 214512
rect 415412 205562 415440 214503
rect 419460 205562 419488 215183
rect 440528 205714 440556 226442
rect 445024 226432 445076 226438
rect 445024 226374 445076 226380
rect 442264 226364 442316 226370
rect 442264 226306 442316 226312
rect 440358 205686 440556 205714
rect 415400 205556 415452 205562
rect 415400 205498 415452 205504
rect 419448 205556 419500 205562
rect 419448 205498 419500 205504
rect 421024 202706 421052 205020
rect 430684 202706 430712 205020
rect 442276 202706 442304 226306
rect 442998 214568 443054 214577
rect 442998 214503 443054 214512
rect 443012 205630 443040 214503
rect 445036 205698 445064 226374
rect 448348 224890 448376 226510
rect 457260 226500 457312 226506
rect 457260 226442 457312 226448
rect 448086 224862 448376 224890
rect 457272 224890 457300 226442
rect 468576 226432 468628 226438
rect 468576 226374 468628 226380
rect 467012 226364 467064 226370
rect 467012 226306 467064 226312
rect 468484 226364 468536 226370
rect 468484 226306 468536 226312
rect 467024 224890 467052 226306
rect 457272 224862 457654 224890
rect 467024 224862 467314 224890
rect 445666 215248 445722 215257
rect 445666 215183 445722 215192
rect 445024 205692 445076 205698
rect 445024 205634 445076 205640
rect 445680 205630 445708 215183
rect 447692 205692 447744 205698
rect 447692 205634 447744 205640
rect 443000 205624 443052 205630
rect 443000 205566 443052 205572
rect 445668 205624 445720 205630
rect 445668 205566 445720 205572
rect 447704 205578 447732 205634
rect 447704 205550 447994 205578
rect 467656 205488 467708 205494
rect 467406 205436 467656 205442
rect 467406 205430 467708 205436
rect 467406 205414 467696 205430
rect 457732 202706 457760 205020
rect 468496 202706 468524 226306
rect 468588 205494 468616 226374
rect 468680 206310 468708 226510
rect 484400 226432 484452 226438
rect 484400 226374 484452 226380
rect 494520 226432 494572 226438
rect 494520 226374 494572 226380
rect 511356 226432 511408 226438
rect 511356 226374 511408 226380
rect 522396 226432 522448 226438
rect 522396 226374 522448 226380
rect 484412 224890 484440 226374
rect 494060 226364 494112 226370
rect 494060 226306 494112 226312
rect 494072 224890 494100 226306
rect 484412 224862 484702 224890
rect 494072 224862 494362 224890
rect 474844 224318 475042 224346
rect 473266 214704 473322 214713
rect 473266 214639 473322 214648
rect 469218 214024 469274 214033
rect 469218 213959 469274 213968
rect 468668 206304 468720 206310
rect 468668 206246 468720 206252
rect 469232 205562 469260 213959
rect 473280 205562 473308 214639
rect 474740 206304 474792 206310
rect 474740 206246 474792 206252
rect 469220 205556 469272 205562
rect 469220 205498 469272 205504
rect 473268 205556 473320 205562
rect 473268 205498 473320 205504
rect 468576 205488 468628 205494
rect 468576 205430 468628 205436
rect 474752 205442 474780 206246
rect 474844 205766 474872 224318
rect 474832 205760 474884 205766
rect 494532 205714 494560 226374
rect 496084 226364 496136 226370
rect 496084 226306 496136 226312
rect 474832 205702 474884 205708
rect 475200 205692 475252 205698
rect 494362 205686 494560 205714
rect 475200 205634 475252 205640
rect 474752 205414 475042 205442
rect 475212 202706 475240 205634
rect 421012 202700 421064 202706
rect 421012 202642 421064 202648
rect 430672 202700 430724 202706
rect 430672 202642 430724 202648
rect 442264 202700 442316 202706
rect 442264 202642 442316 202648
rect 457720 202700 457772 202706
rect 457720 202642 457772 202648
rect 468484 202700 468536 202706
rect 468484 202642 468536 202648
rect 475200 202700 475252 202706
rect 475200 202642 475252 202648
rect 484688 202638 484716 205020
rect 496096 202638 496124 226306
rect 511368 224890 511396 226374
rect 520924 226364 520976 226370
rect 520924 226306 520976 226312
rect 522304 226364 522356 226370
rect 522304 226306 522356 226312
rect 520936 224890 520964 226306
rect 511368 224862 511658 224890
rect 520936 224862 521318 224890
rect 501064 224318 501998 224346
rect 500866 215248 500922 215257
rect 500866 215183 500922 215192
rect 496818 214568 496874 214577
rect 496818 214503 496874 214512
rect 496832 205630 496860 214503
rect 500880 205630 500908 215183
rect 496820 205624 496872 205630
rect 496820 205566 496872 205572
rect 500868 205624 500920 205630
rect 500868 205566 500920 205572
rect 501064 202638 501092 224318
rect 521752 205692 521804 205698
rect 521752 205634 521804 205640
rect 521764 205578 521792 205634
rect 521410 205550 521792 205578
rect 501984 202706 502012 205020
rect 501972 202700 502024 202706
rect 501972 202642 502024 202648
rect 511736 202638 511764 205020
rect 522316 202638 522344 226306
rect 522408 205698 522436 226374
rect 526444 225616 526496 225622
rect 526444 225558 526496 225564
rect 526456 215257 526484 225558
rect 528756 224890 528784 226986
rect 538404 226432 538456 226438
rect 538404 226374 538456 226380
rect 538416 224890 538444 226374
rect 548064 226364 548116 226370
rect 548064 226306 548116 226312
rect 548076 224890 548104 226306
rect 528756 224862 529046 224890
rect 538416 224862 538706 224890
rect 548076 224862 548366 224890
rect 526442 215248 526498 215257
rect 526442 215183 526498 215192
rect 523038 214568 523094 214577
rect 523038 214503 523094 214512
rect 550638 214568 550694 214577
rect 550638 214503 550694 214512
rect 522396 205692 522448 205698
rect 522396 205634 522448 205640
rect 523052 205562 523080 214503
rect 550652 205630 550680 214503
rect 550640 205624 550692 205630
rect 550640 205566 550692 205572
rect 523040 205556 523092 205562
rect 523040 205498 523092 205504
rect 529032 202706 529060 205020
rect 529020 202700 529072 202706
rect 529020 202642 529072 202648
rect 150992 202632 151044 202638
rect 150992 202574 151044 202580
rect 160652 202632 160704 202638
rect 160652 202574 160704 202580
rect 171784 202632 171836 202638
rect 171784 202574 171836 202580
rect 214656 202632 214708 202638
rect 214656 202574 214708 202580
rect 225604 202632 225656 202638
rect 225604 202574 225656 202580
rect 295708 202632 295760 202638
rect 295708 202574 295760 202580
rect 307024 202632 307076 202638
rect 307024 202574 307076 202580
rect 311992 202632 312044 202638
rect 311992 202574 312044 202580
rect 322664 202632 322716 202638
rect 322664 202574 322716 202580
rect 333244 202632 333296 202638
rect 333244 202574 333296 202580
rect 339592 202632 339644 202638
rect 339592 202574 339644 202580
rect 349712 202632 349764 202638
rect 349712 202574 349764 202580
rect 359556 202632 359608 202638
rect 359556 202574 359608 202580
rect 365812 202632 365864 202638
rect 365812 202574 365864 202580
rect 376668 202632 376720 202638
rect 376668 202574 376720 202580
rect 387064 202632 387116 202638
rect 387064 202574 387116 202580
rect 393412 202632 393464 202638
rect 393412 202574 393464 202580
rect 403716 202632 403768 202638
rect 403716 202574 403768 202580
rect 414664 202632 414716 202638
rect 414664 202574 414716 202580
rect 484676 202632 484728 202638
rect 484676 202574 484728 202580
rect 496084 202632 496136 202638
rect 496084 202574 496136 202580
rect 501052 202632 501104 202638
rect 501052 202574 501104 202580
rect 511724 202632 511776 202638
rect 511724 202574 511776 202580
rect 522304 202632 522356 202638
rect 522304 202574 522356 202580
rect 538692 202570 538720 205020
rect 548352 202774 548380 205020
rect 548340 202768 548392 202774
rect 548340 202710 548392 202716
rect 538680 202564 538732 202570
rect 538680 202506 538732 202512
rect 529020 200796 529072 200802
rect 529020 200738 529072 200744
rect 149704 200456 149756 200462
rect 149704 200398 149756 200404
rect 148966 188184 149022 188193
rect 148966 188119 149022 188128
rect 148980 179382 149008 188119
rect 148968 179376 149020 179382
rect 148968 179318 149020 179324
rect 146944 176656 146996 176662
rect 146944 176598 146996 176604
rect 123668 176588 123720 176594
rect 123668 176530 123720 176536
rect 133788 176588 133840 176594
rect 133788 176530 133840 176536
rect 144276 176588 144328 176594
rect 144276 176530 144328 176536
rect 79968 176520 80020 176526
rect 79968 176462 80020 176468
rect 90456 176520 90508 176526
rect 90456 176462 90508 176468
rect 106556 176520 106608 176526
rect 106556 176462 106608 176468
rect 116584 176520 116636 176526
rect 116584 176462 116636 176468
rect 122932 176520 122984 176526
rect 122932 176462 122984 176468
rect 146944 172848 146996 172854
rect 146944 172790 146996 172796
rect 52460 172780 52512 172786
rect 52460 172722 52512 172728
rect 43352 172576 43404 172582
rect 43352 172518 43404 172524
rect 43364 170898 43392 172518
rect 43102 170870 43392 170898
rect 52472 170898 52500 172722
rect 62488 172712 62540 172718
rect 62488 172654 62540 172660
rect 79324 172712 79376 172718
rect 79324 172654 79376 172660
rect 90456 172712 90508 172718
rect 90456 172654 90508 172660
rect 106464 172712 106516 172718
rect 106464 172654 106516 172660
rect 116492 172712 116544 172718
rect 116492 172654 116544 172660
rect 133420 172712 133472 172718
rect 133420 172654 133472 172660
rect 62120 172644 62172 172650
rect 62120 172586 62172 172592
rect 62132 170898 62160 172586
rect 52472 170870 52670 170898
rect 62132 170870 62330 170898
rect 37924 170400 37976 170406
rect 37924 170342 37976 170348
rect 41326 161256 41382 161265
rect 41326 161191 41382 161200
rect 37922 160168 37978 160177
rect 37922 160103 37978 160112
rect 36820 148912 36872 148918
rect 36820 148854 36872 148860
rect 36728 146532 36780 146538
rect 36728 146474 36780 146480
rect 36740 124846 36768 146474
rect 36820 146396 36872 146402
rect 36820 146338 36872 146344
rect 36728 124840 36780 124846
rect 36728 124782 36780 124788
rect 36832 122670 36860 146338
rect 37936 144226 37964 160103
rect 41340 151706 41368 161191
rect 62500 151722 62528 172654
rect 64144 172644 64196 172650
rect 64144 172586 64196 172592
rect 62764 172576 62816 172582
rect 62764 172518 62816 172524
rect 41328 151700 41380 151706
rect 62422 151694 62528 151722
rect 41328 151642 41380 151648
rect 42996 148986 43024 151028
rect 52748 149054 52776 151028
rect 52736 149048 52788 149054
rect 52736 148990 52788 148996
rect 62776 148986 62804 172518
rect 64156 149054 64184 172586
rect 79336 170898 79364 172654
rect 89076 172644 89128 172650
rect 89076 172586 89128 172592
rect 90364 172644 90416 172650
rect 90364 172586 90416 172592
rect 89088 170898 89116 172586
rect 79336 170870 79718 170898
rect 89088 170870 89378 170898
rect 69124 170326 70058 170354
rect 68926 160712 68982 160721
rect 68926 160647 68982 160656
rect 64878 160576 64934 160585
rect 64878 160511 64934 160520
rect 64892 151774 64920 160511
rect 64880 151768 64932 151774
rect 64880 151710 64932 151716
rect 68940 151638 68968 160647
rect 68928 151632 68980 151638
rect 68928 151574 68980 151580
rect 69124 149054 69152 170326
rect 89720 156664 89772 156670
rect 89720 156606 89772 156612
rect 89732 151722 89760 156606
rect 89378 151694 89760 151722
rect 64144 149048 64196 149054
rect 64144 148990 64196 148996
rect 69112 149048 69164 149054
rect 69112 148990 69164 148996
rect 70044 148986 70072 151028
rect 42984 148980 43036 148986
rect 42984 148922 43036 148928
rect 62764 148980 62816 148986
rect 62764 148922 62816 148928
rect 70032 148980 70084 148986
rect 70032 148922 70084 148928
rect 79704 148918 79732 151028
rect 90376 148918 90404 172586
rect 90468 156670 90496 172654
rect 106476 170898 106504 172654
rect 116124 172644 116176 172650
rect 116124 172586 116176 172592
rect 116136 170898 116164 172586
rect 106476 170870 106674 170898
rect 116136 170870 116334 170898
rect 96724 170326 97014 170354
rect 95146 161256 95202 161265
rect 95146 161191 95202 161200
rect 91098 160576 91154 160585
rect 91098 160511 91154 160520
rect 90456 156664 90508 156670
rect 90456 156606 90508 156612
rect 91112 151706 91140 160511
rect 95160 151774 95188 161191
rect 95148 151768 95200 151774
rect 95148 151710 95200 151716
rect 91100 151700 91152 151706
rect 91100 151642 91152 151648
rect 96724 149054 96752 170326
rect 96712 149048 96764 149054
rect 96712 148990 96764 148996
rect 97000 148986 97028 151028
rect 96988 148980 97040 148986
rect 96988 148922 97040 148928
rect 106660 148918 106688 151028
rect 116320 150906 116348 151028
rect 116504 150906 116532 172654
rect 116584 172644 116636 172650
rect 116584 172586 116636 172592
rect 116320 150878 116532 150906
rect 116596 148918 116624 172586
rect 133432 170898 133460 172654
rect 142988 172644 143040 172650
rect 142988 172586 143040 172592
rect 144184 172644 144236 172650
rect 144184 172586 144236 172592
rect 143000 170898 143028 172586
rect 133432 170870 133722 170898
rect 143000 170870 143382 170898
rect 122944 170326 124062 170354
rect 122746 161256 122802 161265
rect 122746 161191 122802 161200
rect 118698 160576 118754 160585
rect 118698 160511 118754 160520
rect 118712 151638 118740 160511
rect 122760 151706 122788 161191
rect 122748 151700 122800 151706
rect 122748 151642 122800 151648
rect 118700 151632 118752 151638
rect 118700 151574 118752 151580
rect 79692 148912 79744 148918
rect 79692 148854 79744 148860
rect 90364 148912 90416 148918
rect 90364 148854 90416 148860
rect 106648 148912 106700 148918
rect 106648 148854 106700 148860
rect 116584 148912 116636 148918
rect 116584 148854 116636 148860
rect 122944 148850 122972 170326
rect 143632 154352 143684 154358
rect 143632 154294 143684 154300
rect 143644 151722 143672 154294
rect 143382 151694 143672 151722
rect 124048 148986 124076 151028
rect 124036 148980 124088 148986
rect 124036 148922 124088 148928
rect 133708 148918 133736 151028
rect 144196 148918 144224 172586
rect 144276 172576 144328 172582
rect 144276 172518 144328 172524
rect 144288 154358 144316 172518
rect 146298 160168 146354 160177
rect 146298 160103 146354 160112
rect 144276 154352 144328 154358
rect 144276 154294 144328 154300
rect 146312 151774 146340 160103
rect 146300 151768 146352 151774
rect 146300 151710 146352 151716
rect 133696 148912 133748 148918
rect 133696 148854 133748 148860
rect 144184 148912 144236 148918
rect 144184 148854 144236 148860
rect 122932 148844 122984 148850
rect 122932 148786 122984 148792
rect 52644 146532 52696 146538
rect 52644 146474 52696 146480
rect 43076 146328 43128 146334
rect 43076 146270 43128 146276
rect 37924 144220 37976 144226
rect 37924 144162 37976 144168
rect 43088 143956 43116 146270
rect 52656 143956 52684 146474
rect 62488 146464 62540 146470
rect 62488 146406 62540 146412
rect 79692 146464 79744 146470
rect 79692 146406 79744 146412
rect 90456 146464 90508 146470
rect 90456 146406 90508 146412
rect 106648 146464 106700 146470
rect 106648 146406 106700 146412
rect 116492 146464 116544 146470
rect 116492 146406 116544 146412
rect 133696 146464 133748 146470
rect 133696 146406 133748 146412
rect 144184 146464 144236 146470
rect 144184 146406 144236 146412
rect 62304 146396 62356 146402
rect 62304 146338 62356 146344
rect 62316 143956 62344 146338
rect 41326 134192 41382 134201
rect 41326 134127 41382 134136
rect 37922 132968 37978 132977
rect 37922 132903 37978 132912
rect 36820 122664 36872 122670
rect 36820 122606 36872 122612
rect 36636 122528 36688 122534
rect 36636 122470 36688 122476
rect 36820 118924 36872 118930
rect 36820 118866 36872 118872
rect 36636 118788 36688 118794
rect 36636 118730 36688 118736
rect 36648 95062 36676 118730
rect 36728 116136 36780 116142
rect 36728 116078 36780 116084
rect 36636 95056 36688 95062
rect 36636 94998 36688 95004
rect 36544 94920 36596 94926
rect 36544 94862 36596 94868
rect 15292 91792 15344 91798
rect 15292 91734 15344 91740
rect 25688 91384 25740 91390
rect 25688 91326 25740 91332
rect 25700 89964 25728 91326
rect 36544 91316 36596 91322
rect 36544 91258 36596 91264
rect 15212 89270 16054 89298
rect 35374 89270 35664 89298
rect 13728 88392 13780 88398
rect 13728 88334 13780 88340
rect 13740 80345 13768 88334
rect 13726 80336 13782 80345
rect 13726 80271 13782 80280
rect 15212 68950 15240 89270
rect 35636 88466 35664 89270
rect 35624 88460 35676 88466
rect 35624 88402 35676 88408
rect 36556 74534 36584 91258
rect 36636 88460 36688 88466
rect 36636 88402 36688 88408
rect 35912 74506 36584 74534
rect 35912 71482 35940 74506
rect 35728 71454 35940 71482
rect 35728 70666 35756 71454
rect 35374 70638 35756 70666
rect 16054 70094 16344 70122
rect 25714 70094 26004 70122
rect 15200 68944 15252 68950
rect 15200 68886 15252 68892
rect 16316 65550 16344 70094
rect 25976 68882 26004 70094
rect 25964 68876 26016 68882
rect 25964 68818 26016 68824
rect 16304 65544 16356 65550
rect 16304 65486 16356 65492
rect 26056 65204 26108 65210
rect 26056 65146 26108 65152
rect 26068 62914 26096 65146
rect 25714 62886 26096 62914
rect 15212 62206 16054 62234
rect 35374 62206 36032 62234
rect 13726 53272 13782 53281
rect 13726 53207 13782 53216
rect 13740 44130 13768 53207
rect 13728 44124 13780 44130
rect 13728 44066 13780 44072
rect 15212 41342 15240 62206
rect 36004 55214 36032 62206
rect 36004 55186 36584 55214
rect 35624 44056 35676 44062
rect 35624 43998 35676 44004
rect 35636 43738 35664 43998
rect 35374 43710 35664 43738
rect 15200 41336 15252 41342
rect 15200 41278 15252 41284
rect 16040 38078 16068 43044
rect 25700 41274 25728 43044
rect 25688 41268 25740 41274
rect 25688 41210 25740 41216
rect 16028 38072 16080 38078
rect 16028 38014 16080 38020
rect 35348 38004 35400 38010
rect 35348 37946 35400 37952
rect 25688 37936 25740 37942
rect 25688 37878 25740 37884
rect 25700 35972 25728 37878
rect 35360 35972 35388 37946
rect 15212 35278 16054 35306
rect 13728 34536 13780 34542
rect 13728 34478 13780 34484
rect 13740 26353 13768 34478
rect 13726 26344 13782 26353
rect 13726 26279 13782 26288
rect 15212 13666 15240 35278
rect 35624 16584 35676 16590
rect 35374 16532 35624 16538
rect 35374 16526 35676 16532
rect 35374 16510 35664 16526
rect 16054 16102 16344 16130
rect 25714 16102 26004 16130
rect 15200 13660 15252 13666
rect 15200 13602 15252 13608
rect 16316 13462 16344 16102
rect 25976 13598 26004 16102
rect 36556 13734 36584 55186
rect 36648 41138 36676 88402
rect 36740 68746 36768 116078
rect 36832 97714 36860 118866
rect 37936 116618 37964 132903
rect 41340 125526 41368 134127
rect 41328 125520 41380 125526
rect 41328 125462 41380 125468
rect 62500 124794 62528 146406
rect 64144 146396 64196 146402
rect 64144 146338 64196 146344
rect 62764 146328 62816 146334
rect 62764 146270 62816 146276
rect 62422 124766 62528 124794
rect 42812 124086 43010 124114
rect 52762 124086 53144 124114
rect 42812 122738 42840 124086
rect 53116 122738 53144 124086
rect 62776 122806 62804 146270
rect 62764 122800 62816 122806
rect 62764 122742 62816 122748
rect 64156 122738 64184 146338
rect 79704 143956 79732 146406
rect 89352 146396 89404 146402
rect 89352 146338 89404 146344
rect 90364 146396 90416 146402
rect 90364 146338 90416 146344
rect 89364 143956 89392 146338
rect 69124 143262 70058 143290
rect 68926 133920 68982 133929
rect 68926 133855 68982 133864
rect 64878 133512 64934 133521
rect 64878 133447 64934 133456
rect 64892 125594 64920 133447
rect 64880 125588 64932 125594
rect 64880 125530 64932 125536
rect 68940 125458 68968 133855
rect 68928 125452 68980 125458
rect 68928 125394 68980 125400
rect 69124 122738 69152 143262
rect 89720 128308 89772 128314
rect 89720 128250 89772 128256
rect 89732 124794 89760 128250
rect 89378 124766 89760 124794
rect 69768 124086 70058 124114
rect 79718 124086 80008 124114
rect 69768 122806 69796 124086
rect 69756 122800 69808 122806
rect 69756 122742 69808 122748
rect 42800 122732 42852 122738
rect 42800 122674 42852 122680
rect 53104 122732 53156 122738
rect 53104 122674 53156 122680
rect 64144 122732 64196 122738
rect 64144 122674 64196 122680
rect 69112 122732 69164 122738
rect 69112 122674 69164 122680
rect 79980 122670 80008 124086
rect 90376 122670 90404 146338
rect 90468 128314 90496 146406
rect 106660 143956 106688 146406
rect 116308 146396 116360 146402
rect 116308 146338 116360 146344
rect 116320 143956 116348 146338
rect 96724 143262 97014 143290
rect 95146 134192 95202 134201
rect 95146 134127 95202 134136
rect 91098 133512 91154 133521
rect 91098 133447 91154 133456
rect 90456 128308 90508 128314
rect 90456 128250 90508 128256
rect 91112 125526 91140 133447
rect 95160 125594 95188 134127
rect 96724 132494 96752 143262
rect 96632 132466 96752 132494
rect 95148 125588 95200 125594
rect 95148 125530 95200 125536
rect 91100 125520 91152 125526
rect 91100 125462 91152 125468
rect 96632 122806 96660 132466
rect 116228 124642 116334 124658
rect 116504 124642 116532 146406
rect 116584 146396 116636 146402
rect 116584 146338 116636 146344
rect 116216 124636 116334 124642
rect 116268 124630 116334 124636
rect 116492 124636 116544 124642
rect 116216 124578 116268 124584
rect 116492 124578 116544 124584
rect 96724 124086 97014 124114
rect 106568 124086 106674 124114
rect 96620 122800 96672 122806
rect 96620 122742 96672 122748
rect 96724 122738 96752 124086
rect 96712 122732 96764 122738
rect 96712 122674 96764 122680
rect 106568 122670 106596 124086
rect 116596 122670 116624 146338
rect 133708 143956 133736 146406
rect 143356 146396 143408 146402
rect 143356 146338 143408 146344
rect 143368 143956 143396 146338
rect 122944 143262 124062 143290
rect 122746 134192 122802 134201
rect 122746 134127 122802 134136
rect 118698 133512 118754 133521
rect 118698 133447 118754 133456
rect 118712 125458 118740 133447
rect 122760 125526 122788 134127
rect 122748 125520 122800 125526
rect 122748 125462 122800 125468
rect 118700 125452 118752 125458
rect 118700 125394 118752 125400
rect 122944 122670 122972 143262
rect 144196 132494 144224 146406
rect 144276 146396 144328 146402
rect 144276 146338 144328 146344
rect 143736 132466 144224 132494
rect 143736 124794 143764 132466
rect 143382 124766 143764 124794
rect 123680 124086 124062 124114
rect 133722 124086 133828 124114
rect 123680 122738 123708 124086
rect 133800 122738 133828 124086
rect 144288 122738 144316 146338
rect 146298 132968 146354 132977
rect 146298 132903 146354 132912
rect 146312 125594 146340 132903
rect 146300 125588 146352 125594
rect 146300 125530 146352 125536
rect 146956 122738 146984 172790
rect 148966 161256 149022 161265
rect 148966 161191 149022 161200
rect 148980 151774 149008 161191
rect 148968 151768 149020 151774
rect 148968 151710 149020 151716
rect 149716 148986 149744 200398
rect 232044 200388 232096 200394
rect 232044 200330 232096 200336
rect 251824 200388 251876 200394
rect 251824 200330 251876 200336
rect 160652 200320 160704 200326
rect 160652 200262 160704 200268
rect 170496 200320 170548 200326
rect 170496 200262 170548 200268
rect 187700 200320 187752 200326
rect 187700 200262 187752 200268
rect 197452 200320 197504 200326
rect 197452 200262 197504 200268
rect 214656 200320 214708 200326
rect 214656 200262 214708 200268
rect 224500 200320 224552 200326
rect 224500 200262 224552 200268
rect 160664 197948 160692 200262
rect 170312 200252 170364 200258
rect 170312 200194 170364 200200
rect 170324 197948 170352 200194
rect 150544 197254 151018 197282
rect 150544 176594 150572 197254
rect 150728 178078 151018 178106
rect 160572 178078 160678 178106
rect 170232 178078 170338 178106
rect 150532 176588 150584 176594
rect 150532 176530 150584 176536
rect 150728 176526 150756 178078
rect 150716 176520 150768 176526
rect 150716 176462 150768 176468
rect 160572 176458 160600 178078
rect 170232 177970 170260 178078
rect 170508 177970 170536 200262
rect 178040 200252 178092 200258
rect 178040 200194 178092 200200
rect 171784 200184 171836 200190
rect 171784 200126 171836 200132
rect 170232 177942 170536 177970
rect 171796 176458 171824 200126
rect 178052 197948 178080 200194
rect 187712 197948 187740 200262
rect 197360 200184 197412 200190
rect 197360 200126 197412 200132
rect 197372 197948 197400 200126
rect 176566 187776 176622 187785
rect 176566 187711 176622 187720
rect 172518 187504 172574 187513
rect 172518 187439 172574 187448
rect 172532 179314 172560 187439
rect 176580 179314 176608 187711
rect 172520 179308 172572 179314
rect 172520 179250 172572 179256
rect 176568 179308 176620 179314
rect 176568 179250 176620 179256
rect 197464 178786 197492 200262
rect 200764 200252 200816 200258
rect 200764 200194 200816 200200
rect 199384 200184 199436 200190
rect 199384 200126 199436 200132
rect 197386 178758 197492 178786
rect 178066 178078 178172 178106
rect 187726 178078 188016 178106
rect 178144 176526 178172 178078
rect 187988 176526 188016 178078
rect 199396 176526 199424 200126
rect 200118 187504 200174 187513
rect 200118 187439 200174 187448
rect 200132 179382 200160 187439
rect 200120 179376 200172 179382
rect 200120 179318 200172 179324
rect 200776 176662 200804 200194
rect 214668 197948 214696 200262
rect 224316 200184 224368 200190
rect 224316 200126 224368 200132
rect 224328 197948 224356 200126
rect 204364 197254 205022 197282
rect 202786 188184 202842 188193
rect 202786 188119 202842 188128
rect 202800 179382 202828 188119
rect 202788 179376 202840 179382
rect 202788 179318 202840 179324
rect 200764 176656 200816 176662
rect 200764 176598 200816 176604
rect 204364 176526 204392 197254
rect 224512 178786 224540 200262
rect 225604 200184 225656 200190
rect 225604 200126 225656 200132
rect 224342 178758 224540 178786
rect 204640 178078 205022 178106
rect 214682 178078 215064 178106
rect 204640 176662 204668 178078
rect 204628 176656 204680 176662
rect 204628 176598 204680 176604
rect 178132 176520 178184 176526
rect 178132 176462 178184 176468
rect 187976 176520 188028 176526
rect 187976 176462 188028 176468
rect 199384 176520 199436 176526
rect 199384 176462 199436 176468
rect 204352 176520 204404 176526
rect 204352 176462 204404 176468
rect 215036 176458 215064 178078
rect 225616 176458 225644 200126
rect 232056 197948 232084 200330
rect 241704 200320 241756 200326
rect 241704 200262 241756 200268
rect 241716 197948 241744 200262
rect 251456 200252 251508 200258
rect 251456 200194 251508 200200
rect 251364 200184 251416 200190
rect 251364 200126 251416 200132
rect 251376 197948 251404 200126
rect 230386 188184 230442 188193
rect 230386 188119 230442 188128
rect 226338 187504 226394 187513
rect 226338 187439 226394 187448
rect 226352 179314 226380 187439
rect 230400 179314 230428 188119
rect 226340 179308 226392 179314
rect 226340 179250 226392 179256
rect 230388 179308 230440 179314
rect 230388 179250 230440 179256
rect 251468 178786 251496 200194
rect 251390 178758 251496 178786
rect 231872 178078 232070 178106
rect 241730 178078 242112 178106
rect 231872 176526 231900 178078
rect 242084 176526 242112 178078
rect 251836 176662 251864 200330
rect 413468 200320 413520 200326
rect 413468 200262 413520 200268
rect 430672 200320 430724 200326
rect 430672 200262 430724 200268
rect 440516 200320 440568 200326
rect 440516 200262 440568 200268
rect 457628 200320 457680 200326
rect 457628 200262 457680 200268
rect 468576 200320 468628 200326
rect 468576 200262 468628 200268
rect 484676 200320 484728 200326
rect 484676 200262 484728 200268
rect 494520 200320 494572 200326
rect 494520 200262 494572 200268
rect 511632 200320 511684 200326
rect 511632 200262 511684 200268
rect 268660 200252 268712 200258
rect 268660 200194 268712 200200
rect 279424 200252 279476 200258
rect 279424 200194 279476 200200
rect 295708 200252 295760 200258
rect 295708 200194 295760 200200
rect 305460 200252 305512 200258
rect 305460 200194 305512 200200
rect 322664 200252 322716 200258
rect 322664 200194 322716 200200
rect 336004 200252 336056 200258
rect 336004 200194 336056 200200
rect 349712 200252 349764 200258
rect 349712 200194 349764 200200
rect 359464 200252 359516 200258
rect 359464 200194 359516 200200
rect 376668 200252 376720 200258
rect 376668 200194 376720 200200
rect 386512 200252 386564 200258
rect 386512 200194 386564 200200
rect 403624 200252 403676 200258
rect 403624 200194 403676 200200
rect 253204 200184 253256 200190
rect 253204 200126 253256 200132
rect 251824 176656 251876 176662
rect 251824 176598 251876 176604
rect 253216 176526 253244 200126
rect 268672 197948 268700 200194
rect 278320 200184 278372 200190
rect 278320 200126 278372 200132
rect 278332 197948 278360 200126
rect 258184 197254 259026 197282
rect 256606 188184 256662 188193
rect 256606 188119 256662 188128
rect 253938 186960 253994 186969
rect 253938 186895 253994 186904
rect 253952 179382 253980 186895
rect 256620 179382 256648 188119
rect 253940 179376 253992 179382
rect 253940 179318 253992 179324
rect 256608 179376 256660 179382
rect 256608 179318 256660 179324
rect 258184 176526 258212 197254
rect 279436 180794 279464 200194
rect 279516 200184 279568 200190
rect 279516 200126 279568 200132
rect 278792 180766 279464 180794
rect 278792 178786 278820 180766
rect 278346 178758 278820 178786
rect 258736 178078 259026 178106
rect 268686 178078 268976 178106
rect 258736 176662 258764 178078
rect 258724 176656 258776 176662
rect 258724 176598 258776 176604
rect 231860 176520 231912 176526
rect 231860 176462 231912 176468
rect 242072 176520 242124 176526
rect 242072 176462 242124 176468
rect 253204 176520 253256 176526
rect 253204 176462 253256 176468
rect 258172 176520 258224 176526
rect 258172 176462 258224 176468
rect 268948 176458 268976 178078
rect 279528 176458 279556 200126
rect 285784 198070 286088 198098
rect 284206 187776 284262 187785
rect 284206 187711 284262 187720
rect 280158 187504 280214 187513
rect 280158 187439 280214 187448
rect 280172 179314 280200 187439
rect 284220 179314 284248 187711
rect 280160 179308 280212 179314
rect 280160 179250 280212 179256
rect 284208 179308 284260 179314
rect 284208 179250 284260 179256
rect 285784 176458 285812 198070
rect 286060 197948 286088 198070
rect 295720 197948 295748 200194
rect 305368 200184 305420 200190
rect 305368 200126 305420 200132
rect 305380 197948 305408 200126
rect 305472 178786 305500 200194
rect 307024 200184 307076 200190
rect 307024 200126 307076 200132
rect 305394 178758 305500 178786
rect 286074 178078 286180 178106
rect 295734 178078 296024 178106
rect 286152 176526 286180 178078
rect 286140 176520 286192 176526
rect 286140 176462 286192 176468
rect 295996 176458 296024 178078
rect 307036 176458 307064 200126
rect 322676 197948 322704 200194
rect 332324 200184 332376 200190
rect 332324 200126 332376 200132
rect 333244 200184 333296 200190
rect 333244 200126 333296 200132
rect 332336 197948 332364 200126
rect 312004 197254 313030 197282
rect 311806 188184 311862 188193
rect 311806 188119 311862 188128
rect 307758 187504 307814 187513
rect 307758 187439 307814 187448
rect 307772 179382 307800 187439
rect 307760 179376 307812 179382
rect 307760 179318 307812 179324
rect 311820 179246 311848 188119
rect 311808 179240 311860 179246
rect 311808 179182 311860 179188
rect 312004 176458 312032 197254
rect 312648 178078 313030 178106
rect 322690 178078 322888 178106
rect 332350 178078 332548 178106
rect 312648 176526 312676 178078
rect 312636 176520 312688 176526
rect 312636 176462 312688 176468
rect 322860 176458 322888 178078
rect 332520 176662 332548 178078
rect 332508 176656 332560 176662
rect 332508 176598 332560 176604
rect 333256 176458 333284 200126
rect 335358 187504 335414 187513
rect 335358 187439 335414 187448
rect 335372 179314 335400 187439
rect 335360 179308 335412 179314
rect 335360 179250 335412 179256
rect 336016 176662 336044 200194
rect 339604 198070 340092 198098
rect 338026 188184 338082 188193
rect 338026 188119 338082 188128
rect 338040 179382 338068 188119
rect 338028 179376 338080 179382
rect 338028 179318 338080 179324
rect 336004 176656 336056 176662
rect 336004 176598 336056 176604
rect 339604 176458 339632 198070
rect 340064 197948 340092 198070
rect 349724 197948 349752 200194
rect 359372 200184 359424 200190
rect 359372 200126 359424 200132
rect 359384 197948 359412 200126
rect 359476 178786 359504 200194
rect 359556 200184 359608 200190
rect 359556 200126 359608 200132
rect 359398 178758 359504 178786
rect 340078 178078 340184 178106
rect 349738 178078 350120 178106
rect 340156 176526 340184 178078
rect 340144 176520 340196 176526
rect 340144 176462 340196 176468
rect 350092 176458 350120 178078
rect 359568 176458 359596 200126
rect 376680 197948 376708 200194
rect 386328 200184 386380 200190
rect 386328 200126 386380 200132
rect 386340 197948 386368 200126
rect 365824 197254 367034 197282
rect 365626 188184 365682 188193
rect 365626 188119 365682 188128
rect 361578 186960 361634 186969
rect 361578 186895 361634 186904
rect 361592 179246 361620 186895
rect 365640 179314 365668 188119
rect 365628 179308 365680 179314
rect 365628 179250 365680 179256
rect 361580 179240 361632 179246
rect 361580 179182 361632 179188
rect 365824 176458 365852 197254
rect 386524 178786 386552 200194
rect 387064 200184 387116 200190
rect 387064 200126 387116 200132
rect 386354 178758 386552 178786
rect 366744 178078 367034 178106
rect 376588 178078 376694 178106
rect 366744 176526 366772 178078
rect 366732 176520 366784 176526
rect 366732 176462 366784 176468
rect 376588 176458 376616 178078
rect 387076 176458 387104 200126
rect 403636 197948 403664 200194
rect 413284 200184 413336 200190
rect 413284 200126 413336 200132
rect 413296 197948 413324 200126
rect 393424 197254 393990 197282
rect 391846 187776 391902 187785
rect 391846 187711 391902 187720
rect 389178 187504 389234 187513
rect 389178 187439 389234 187448
rect 389192 179382 389220 187439
rect 391860 179382 391888 187711
rect 389180 179376 389232 179382
rect 389180 179318 389232 179324
rect 391848 179376 391900 179382
rect 391848 179318 391900 179324
rect 393424 176458 393452 197254
rect 413480 178786 413508 200262
rect 421012 200252 421064 200258
rect 421012 200194 421064 200200
rect 414664 200184 414716 200190
rect 414664 200126 414716 200132
rect 413402 178758 413508 178786
rect 393608 178078 393990 178106
rect 403742 178078 404032 178106
rect 393608 176526 393636 178078
rect 393596 176520 393648 176526
rect 393596 176462 393648 176468
rect 404004 176458 404032 178078
rect 414676 176458 414704 200126
rect 421024 197948 421052 200194
rect 430684 197948 430712 200262
rect 440332 200184 440384 200190
rect 440332 200126 440384 200132
rect 440344 197948 440372 200126
rect 419446 188184 419502 188193
rect 419446 188119 419502 188128
rect 415398 187504 415454 187513
rect 415398 187439 415454 187448
rect 415412 179314 415440 187439
rect 419460 179314 419488 188119
rect 415400 179308 415452 179314
rect 415400 179250 415452 179256
rect 419448 179308 419500 179314
rect 419448 179250 419500 179256
rect 440528 178786 440556 200262
rect 446404 200252 446456 200258
rect 446404 200194 446456 200200
rect 442264 200184 442316 200190
rect 442264 200126 442316 200132
rect 440358 178758 440556 178786
rect 420932 178078 421038 178106
rect 430698 178078 431080 178106
rect 420932 176526 420960 178078
rect 431052 176526 431080 178078
rect 442276 176526 442304 200126
rect 445666 188184 445722 188193
rect 445666 188119 445722 188128
rect 442998 186960 443054 186969
rect 442998 186895 443054 186904
rect 443012 179382 443040 186895
rect 445680 179450 445708 188119
rect 445668 179444 445720 179450
rect 445668 179386 445720 179392
rect 446416 179382 446444 200194
rect 457640 197948 457668 200262
rect 467288 200184 467340 200190
rect 467288 200126 467340 200132
rect 468484 200184 468536 200190
rect 468484 200126 468536 200132
rect 467300 197948 467328 200126
rect 447244 197254 447994 197282
rect 443000 179376 443052 179382
rect 443000 179318 443052 179324
rect 446404 179376 446456 179382
rect 446404 179318 446456 179324
rect 447244 176526 447272 197254
rect 447692 179376 447744 179382
rect 447692 179318 447744 179324
rect 447704 178786 447732 179318
rect 467656 179240 467708 179246
rect 467656 179182 467708 179188
rect 467668 178786 467696 179182
rect 447704 178758 447994 178786
rect 467406 178758 467696 178786
rect 457746 178078 458128 178106
rect 420920 176520 420972 176526
rect 420920 176462 420972 176468
rect 431040 176520 431092 176526
rect 431040 176462 431092 176468
rect 442264 176520 442316 176526
rect 442264 176462 442316 176468
rect 447232 176520 447284 176526
rect 447232 176462 447284 176468
rect 458100 176458 458128 178078
rect 468496 176458 468524 200126
rect 468588 179246 468616 200262
rect 475016 200252 475068 200258
rect 475016 200194 475068 200200
rect 475028 197948 475056 200194
rect 484688 197948 484716 200262
rect 494336 200184 494388 200190
rect 494336 200126 494388 200132
rect 494348 197948 494376 200126
rect 473266 187776 473322 187785
rect 473266 187711 473322 187720
rect 469218 186960 469274 186969
rect 469218 186895 469274 186904
rect 469232 179314 469260 186895
rect 473280 179314 473308 187711
rect 469220 179308 469272 179314
rect 469220 179250 469272 179256
rect 473268 179308 473320 179314
rect 473268 179250 473320 179256
rect 468576 179240 468628 179246
rect 468576 179182 468628 179188
rect 494532 178786 494560 200262
rect 494704 200252 494756 200258
rect 494704 200194 494756 200200
rect 494362 178758 494560 178786
rect 474752 178078 475042 178106
rect 484702 178078 484992 178106
rect 474752 176526 474780 178078
rect 484964 176526 484992 178078
rect 494716 176662 494744 200194
rect 496084 200184 496136 200190
rect 496084 200126 496136 200132
rect 494704 176656 494756 176662
rect 494704 176598 494756 176604
rect 496096 176526 496124 200126
rect 511644 197948 511672 200262
rect 522396 200252 522448 200258
rect 522396 200194 522448 200200
rect 521292 200184 521344 200190
rect 521292 200126 521344 200132
rect 522304 200184 522356 200190
rect 522304 200126 522356 200132
rect 521304 197948 521332 200126
rect 501064 197254 501998 197282
rect 500866 187776 500922 187785
rect 500866 187711 500922 187720
rect 496818 187504 496874 187513
rect 496818 187439 496874 187448
rect 496832 179382 496860 187439
rect 500880 179382 500908 187711
rect 496820 179376 496872 179382
rect 496820 179318 496872 179324
rect 500868 179376 500920 179382
rect 500868 179318 500920 179324
rect 501064 176526 501092 197254
rect 521752 179444 521804 179450
rect 521752 179386 521804 179392
rect 521764 178786 521792 179386
rect 521410 178758 521792 178786
rect 501616 178078 501998 178106
rect 511750 178078 511948 178106
rect 501616 176662 501644 178078
rect 501604 176656 501656 176662
rect 501604 176598 501656 176604
rect 474740 176520 474792 176526
rect 474740 176462 474792 176468
rect 484952 176520 485004 176526
rect 484952 176462 485004 176468
rect 496084 176520 496136 176526
rect 496084 176462 496136 176468
rect 501052 176520 501104 176526
rect 501052 176462 501104 176468
rect 511920 176458 511948 178078
rect 522316 176458 522344 200126
rect 522408 179450 522436 200194
rect 526444 198008 526496 198014
rect 526444 197950 526496 197956
rect 526456 188329 526484 197950
rect 529032 197948 529060 200738
rect 538680 200252 538732 200258
rect 538680 200194 538732 200200
rect 538692 197948 538720 200194
rect 548340 200184 548392 200190
rect 548340 200126 548392 200132
rect 548352 197948 548380 200126
rect 526442 188320 526498 188329
rect 526442 188255 526498 188264
rect 523038 187504 523094 187513
rect 523038 187439 523094 187448
rect 522396 179444 522448 179450
rect 522396 179386 522448 179392
rect 523052 179314 523080 187439
rect 550638 186960 550694 186969
rect 550638 186895 550694 186904
rect 550652 179382 550680 186895
rect 550640 179376 550692 179382
rect 550640 179318 550692 179324
rect 523040 179308 523092 179314
rect 523040 179250 523092 179256
rect 528664 178078 529046 178106
rect 538416 178078 538706 178106
rect 547984 178078 548366 178106
rect 528664 176526 528692 178078
rect 528652 176520 528704 176526
rect 528652 176462 528704 176468
rect 160560 176452 160612 176458
rect 160560 176394 160612 176400
rect 171784 176452 171836 176458
rect 171784 176394 171836 176400
rect 215024 176452 215076 176458
rect 215024 176394 215076 176400
rect 225604 176452 225656 176458
rect 225604 176394 225656 176400
rect 268936 176452 268988 176458
rect 268936 176394 268988 176400
rect 279516 176452 279568 176458
rect 279516 176394 279568 176400
rect 285772 176452 285824 176458
rect 285772 176394 285824 176400
rect 295984 176452 296036 176458
rect 295984 176394 296036 176400
rect 307024 176452 307076 176458
rect 307024 176394 307076 176400
rect 311992 176452 312044 176458
rect 311992 176394 312044 176400
rect 322848 176452 322900 176458
rect 322848 176394 322900 176400
rect 333244 176452 333296 176458
rect 333244 176394 333296 176400
rect 339592 176452 339644 176458
rect 339592 176394 339644 176400
rect 350080 176452 350132 176458
rect 350080 176394 350132 176400
rect 359556 176452 359608 176458
rect 359556 176394 359608 176400
rect 365812 176452 365864 176458
rect 365812 176394 365864 176400
rect 376576 176452 376628 176458
rect 376576 176394 376628 176400
rect 387064 176452 387116 176458
rect 387064 176394 387116 176400
rect 393412 176452 393464 176458
rect 393412 176394 393464 176400
rect 403992 176452 404044 176458
rect 403992 176394 404044 176400
rect 414664 176452 414716 176458
rect 414664 176394 414716 176400
rect 458088 176452 458140 176458
rect 458088 176394 458140 176400
rect 468484 176452 468536 176458
rect 468484 176394 468536 176400
rect 511908 176452 511960 176458
rect 511908 176394 511960 176400
rect 522304 176452 522356 176458
rect 522304 176394 522356 176400
rect 538416 176390 538444 178078
rect 547984 176594 548012 178078
rect 547972 176588 548024 176594
rect 547972 176530 548024 176536
rect 538404 176384 538456 176390
rect 538404 176326 538456 176332
rect 528652 173188 528704 173194
rect 528652 173130 528704 173136
rect 232320 172780 232372 172786
rect 232320 172722 232372 172728
rect 251824 172780 251876 172786
rect 251824 172722 251876 172728
rect 475384 172780 475436 172786
rect 475384 172722 475436 172728
rect 494704 172780 494756 172786
rect 494704 172722 494756 172728
rect 170496 172712 170548 172718
rect 170496 172654 170548 172660
rect 187792 172712 187844 172718
rect 187792 172654 187844 172660
rect 197544 172712 197596 172718
rect 197544 172654 197596 172660
rect 214380 172712 214432 172718
rect 214380 172654 214432 172660
rect 224500 172712 224552 172718
rect 224500 172654 224552 172660
rect 170036 172644 170088 172650
rect 170036 172586 170088 172592
rect 160284 172576 160336 172582
rect 160284 172518 160336 172524
rect 160296 170898 160324 172518
rect 170048 170898 170076 172586
rect 160296 170870 160678 170898
rect 170048 170870 170338 170898
rect 150544 170326 151018 170354
rect 149704 148980 149756 148986
rect 149704 148922 149756 148928
rect 150544 148918 150572 170326
rect 150532 148912 150584 148918
rect 150532 148854 150584 148860
rect 151004 148850 151032 151028
rect 160664 148850 160692 151028
rect 170324 150906 170352 151028
rect 170508 150906 170536 172654
rect 178408 172644 178460 172650
rect 178408 172586 178460 172592
rect 171784 172576 171836 172582
rect 171784 172518 171836 172524
rect 170324 150878 170536 150906
rect 171796 148850 171824 172518
rect 178420 170898 178448 172586
rect 187804 170898 187832 172654
rect 197452 172576 197504 172582
rect 197452 172518 197504 172524
rect 197464 170898 197492 172518
rect 178066 170870 178448 170898
rect 187726 170870 187832 170898
rect 197386 170870 197492 170898
rect 197556 161474 197584 172654
rect 200764 172644 200816 172650
rect 200764 172586 200816 172592
rect 199384 172576 199436 172582
rect 199384 172518 199436 172524
rect 197464 161446 197584 161474
rect 176566 160712 176622 160721
rect 176566 160647 176622 160656
rect 172518 160576 172574 160585
rect 172518 160511 172574 160520
rect 172532 151706 172560 160511
rect 176580 151706 176608 160647
rect 197464 151722 197492 161446
rect 172520 151700 172572 151706
rect 172520 151642 172572 151648
rect 176568 151700 176620 151706
rect 197386 151694 197492 151722
rect 176568 151642 176620 151648
rect 178052 148918 178080 151028
rect 187712 148918 187740 151028
rect 199396 148918 199424 172518
rect 200118 160576 200174 160585
rect 200118 160511 200174 160520
rect 200132 151774 200160 160511
rect 200120 151768 200172 151774
rect 200120 151710 200172 151716
rect 200776 151638 200804 172586
rect 214392 170898 214420 172654
rect 223948 172576 224000 172582
rect 223948 172518 224000 172524
rect 223960 170898 223988 172518
rect 214392 170870 214682 170898
rect 223960 170870 224342 170898
rect 204364 170326 205022 170354
rect 202786 161256 202842 161265
rect 202786 161191 202842 161200
rect 202800 151774 202828 161191
rect 202788 151768 202840 151774
rect 202788 151710 202840 151716
rect 200764 151632 200816 151638
rect 200764 151574 200816 151580
rect 204364 148918 204392 170326
rect 224512 151722 224540 172654
rect 225604 172576 225656 172582
rect 225604 172518 225656 172524
rect 224342 151694 224540 151722
rect 204628 151632 204680 151638
rect 204680 151580 205022 151586
rect 204628 151574 205022 151580
rect 204640 151558 205022 151574
rect 178040 148912 178092 148918
rect 178040 148854 178092 148860
rect 187700 148912 187752 148918
rect 187700 148854 187752 148860
rect 199384 148912 199436 148918
rect 199384 148854 199436 148860
rect 204352 148912 204404 148918
rect 204352 148854 204404 148860
rect 214668 148850 214696 151028
rect 225616 148850 225644 172518
rect 232332 170898 232360 172722
rect 241612 172712 241664 172718
rect 241612 172654 241664 172660
rect 232070 170870 232360 170898
rect 241624 170898 241652 172654
rect 251456 172644 251508 172650
rect 251456 172586 251508 172592
rect 251272 172576 251324 172582
rect 251272 172518 251324 172524
rect 251284 170898 251312 172518
rect 241624 170870 241730 170898
rect 251284 170870 251390 170898
rect 230386 161256 230442 161265
rect 230386 161191 230442 161200
rect 226338 160576 226394 160585
rect 226338 160511 226394 160520
rect 226352 151706 226380 160511
rect 230400 151706 230428 161191
rect 251468 151722 251496 172586
rect 226340 151700 226392 151706
rect 226340 151642 226392 151648
rect 230388 151700 230440 151706
rect 251390 151694 251496 151722
rect 230388 151642 230440 151648
rect 232056 148918 232084 151028
rect 241716 148918 241744 151028
rect 251836 149054 251864 172722
rect 413468 172712 413520 172718
rect 413468 172654 413520 172660
rect 430580 172712 430632 172718
rect 430580 172654 430632 172660
rect 440516 172712 440568 172718
rect 440516 172654 440568 172660
rect 457260 172712 457312 172718
rect 457260 172654 457312 172660
rect 468484 172712 468536 172718
rect 468484 172654 468536 172660
rect 268292 172644 268344 172650
rect 268292 172586 268344 172592
rect 279424 172644 279476 172650
rect 279424 172586 279476 172592
rect 295800 172644 295852 172650
rect 295800 172586 295852 172592
rect 305552 172644 305604 172650
rect 305552 172586 305604 172592
rect 322388 172644 322440 172650
rect 322388 172586 322440 172592
rect 334624 172644 334676 172650
rect 334624 172586 334676 172592
rect 349804 172644 349856 172650
rect 349804 172586 349856 172592
rect 359648 172644 359700 172650
rect 359648 172586 359700 172592
rect 376300 172644 376352 172650
rect 376300 172586 376352 172592
rect 386512 172644 386564 172650
rect 386512 172586 386564 172592
rect 403348 172644 403400 172650
rect 403348 172586 403400 172592
rect 253204 172576 253256 172582
rect 253204 172518 253256 172524
rect 251824 149048 251876 149054
rect 251824 148990 251876 148996
rect 253216 148918 253244 172518
rect 268304 170898 268332 172586
rect 278044 172576 278096 172582
rect 278044 172518 278096 172524
rect 278056 170898 278084 172518
rect 268304 170870 268686 170898
rect 278056 170870 278346 170898
rect 258184 170326 259026 170354
rect 256606 161256 256662 161265
rect 256606 161191 256662 161200
rect 253938 160168 253994 160177
rect 253938 160103 253994 160112
rect 253952 151774 253980 160103
rect 256620 151774 256648 161191
rect 253940 151768 253992 151774
rect 253940 151710 253992 151716
rect 256608 151768 256660 151774
rect 256608 151710 256660 151716
rect 258184 148918 258212 170326
rect 279436 151814 279464 172586
rect 279516 172576 279568 172582
rect 279516 172518 279568 172524
rect 278792 151786 279464 151814
rect 278792 151722 278820 151786
rect 278346 151694 278820 151722
rect 259012 149054 259040 151028
rect 259000 149048 259052 149054
rect 259000 148990 259052 148996
rect 232044 148912 232096 148918
rect 232044 148854 232096 148860
rect 241704 148912 241756 148918
rect 241704 148854 241756 148860
rect 253204 148912 253256 148918
rect 253204 148854 253256 148860
rect 258172 148912 258224 148918
rect 258172 148854 258224 148860
rect 268672 148850 268700 151028
rect 279528 148850 279556 172518
rect 295812 170898 295840 172586
rect 305460 172576 305512 172582
rect 305460 172518 305512 172524
rect 305472 170898 305500 172518
rect 295734 170870 295840 170898
rect 305394 170870 305500 170898
rect 286074 170338 286180 170354
rect 285772 170332 285824 170338
rect 286074 170332 286192 170338
rect 286074 170326 286140 170332
rect 285772 170274 285824 170280
rect 286140 170274 286192 170280
rect 284206 160712 284262 160721
rect 284206 160647 284262 160656
rect 280158 160576 280214 160585
rect 280158 160511 280214 160520
rect 280172 151706 280200 160511
rect 284220 151706 284248 160647
rect 280160 151700 280212 151706
rect 280160 151642 280212 151648
rect 284208 151700 284260 151706
rect 284208 151642 284260 151648
rect 285784 148850 285812 170274
rect 305564 161474 305592 172586
rect 307024 172576 307076 172582
rect 307024 172518 307076 172524
rect 305472 161446 305592 161474
rect 305472 151722 305500 161446
rect 305394 151694 305500 151722
rect 286060 148918 286088 151028
rect 286048 148912 286100 148918
rect 286048 148854 286100 148860
rect 295720 148850 295748 151028
rect 307036 148850 307064 172518
rect 322400 170898 322428 172586
rect 331956 172576 332008 172582
rect 331956 172518 332008 172524
rect 333244 172576 333296 172582
rect 333244 172518 333296 172524
rect 331968 170898 331996 172518
rect 322400 170870 322690 170898
rect 331968 170870 332350 170898
rect 312004 170326 313030 170354
rect 311806 161256 311862 161265
rect 311806 161191 311862 161200
rect 307758 160576 307814 160585
rect 307758 160511 307814 160520
rect 307772 151774 307800 160511
rect 307760 151768 307812 151774
rect 307760 151710 307812 151716
rect 311820 151638 311848 161191
rect 311808 151632 311860 151638
rect 311808 151574 311860 151580
rect 312004 148850 312032 170326
rect 332508 151768 332560 151774
rect 332350 151716 332508 151722
rect 332350 151710 332560 151716
rect 332350 151694 332548 151710
rect 313016 148918 313044 151028
rect 313004 148912 313056 148918
rect 313004 148854 313056 148860
rect 322676 148850 322704 151028
rect 333256 148850 333284 172518
rect 334636 151774 334664 172586
rect 349816 170898 349844 172586
rect 359464 172576 359516 172582
rect 359464 172518 359516 172524
rect 359556 172576 359608 172582
rect 359556 172518 359608 172524
rect 359476 170898 359504 172518
rect 349738 170870 349844 170898
rect 359398 170870 359504 170898
rect 340078 170338 340184 170354
rect 339592 170332 339644 170338
rect 340078 170332 340196 170338
rect 340078 170326 340144 170332
rect 339592 170274 339644 170280
rect 340144 170274 340196 170280
rect 338026 161256 338082 161265
rect 338026 161191 338082 161200
rect 335358 160576 335414 160585
rect 335358 160511 335414 160520
rect 334624 151768 334676 151774
rect 334624 151710 334676 151716
rect 335372 151706 335400 160511
rect 338040 151774 338068 161191
rect 338028 151768 338080 151774
rect 338028 151710 338080 151716
rect 335360 151700 335412 151706
rect 335360 151642 335412 151648
rect 339604 148850 339632 170274
rect 359568 166394 359596 172518
rect 359556 166388 359608 166394
rect 359556 166330 359608 166336
rect 359660 166274 359688 172586
rect 376312 170898 376340 172586
rect 386052 172576 386104 172582
rect 386052 172518 386104 172524
rect 386064 170898 386092 172518
rect 376312 170870 376694 170898
rect 386064 170870 386354 170898
rect 359476 166246 359688 166274
rect 365824 170326 367034 170354
rect 359476 151722 359504 166246
rect 359556 166184 359608 166190
rect 359556 166126 359608 166132
rect 359398 151694 359504 151722
rect 340064 148918 340092 151028
rect 340052 148912 340104 148918
rect 340052 148854 340104 148860
rect 349724 148850 349752 151028
rect 359568 148850 359596 166126
rect 365626 161256 365682 161265
rect 365626 161191 365682 161200
rect 361578 160168 361634 160177
rect 361578 160103 361634 160112
rect 361592 151638 361620 160103
rect 365640 151706 365668 161191
rect 365628 151700 365680 151706
rect 365628 151642 365680 151648
rect 361580 151632 361632 151638
rect 361580 151574 361632 151580
rect 365824 148850 365852 170326
rect 386524 151722 386552 172586
rect 387064 172576 387116 172582
rect 387064 172518 387116 172524
rect 386354 151694 386552 151722
rect 367020 148918 367048 151028
rect 367008 148912 367060 148918
rect 367008 148854 367060 148860
rect 376680 148850 376708 151028
rect 387076 148850 387104 172518
rect 403360 170898 403388 172586
rect 412916 172576 412968 172582
rect 412916 172518 412968 172524
rect 412928 170898 412956 172518
rect 403360 170870 403650 170898
rect 412928 170870 413310 170898
rect 393424 170326 393990 170354
rect 391846 161256 391902 161265
rect 391846 161191 391902 161200
rect 389178 160576 389234 160585
rect 389178 160511 389234 160520
rect 389192 151774 389220 160511
rect 391860 151774 391888 161191
rect 389180 151768 389232 151774
rect 389180 151710 389232 151716
rect 391848 151768 391900 151774
rect 391848 151710 391900 151716
rect 393424 148850 393452 170326
rect 413480 151722 413508 172654
rect 421288 172644 421340 172650
rect 421288 172586 421340 172592
rect 414664 172576 414716 172582
rect 414664 172518 414716 172524
rect 413402 151694 413508 151722
rect 393976 148918 394004 151028
rect 393964 148912 394016 148918
rect 393964 148854 394016 148860
rect 403728 148850 403756 151028
rect 414676 148850 414704 172518
rect 421300 170898 421328 172586
rect 421038 170870 421328 170898
rect 430592 170898 430620 172654
rect 440240 172576 440292 172582
rect 440240 172518 440292 172524
rect 440252 170898 440280 172518
rect 430592 170870 430698 170898
rect 440252 170870 440358 170898
rect 419446 161256 419502 161265
rect 419446 161191 419502 161200
rect 415398 160576 415454 160585
rect 415398 160511 415454 160520
rect 415412 151706 415440 160511
rect 419460 151706 419488 161191
rect 440528 151722 440556 172654
rect 443644 172644 443696 172650
rect 443644 172586 443696 172592
rect 442264 172576 442316 172582
rect 442264 172518 442316 172524
rect 415400 151700 415452 151706
rect 415400 151642 415452 151648
rect 419448 151700 419500 151706
rect 440358 151694 440556 151722
rect 419448 151642 419500 151648
rect 421024 148918 421052 151028
rect 430684 148918 430712 151028
rect 442276 148918 442304 172518
rect 442998 160576 443054 160585
rect 442998 160511 443054 160520
rect 443012 151774 443040 160511
rect 443000 151768 443052 151774
rect 443000 151710 443052 151716
rect 443656 151638 443684 172586
rect 457272 170898 457300 172654
rect 467012 172576 467064 172582
rect 467012 172518 467064 172524
rect 467024 170898 467052 172518
rect 457272 170870 457654 170898
rect 467024 170870 467314 170898
rect 447244 170326 447994 170354
rect 445666 161256 445722 161265
rect 445666 161191 445722 161200
rect 445680 151774 445708 161191
rect 445668 151768 445720 151774
rect 445668 151710 445720 151716
rect 443644 151632 443696 151638
rect 443644 151574 443696 151580
rect 447244 148918 447272 170326
rect 468496 151814 468524 172654
rect 468576 172576 468628 172582
rect 468576 172518 468628 172524
rect 467760 151786 468524 151814
rect 467760 151722 467788 151786
rect 467406 151694 467788 151722
rect 447692 151632 447744 151638
rect 447744 151580 447994 151586
rect 447692 151574 447994 151580
rect 447704 151558 447994 151574
rect 421012 148912 421064 148918
rect 421012 148854 421064 148860
rect 430672 148912 430724 148918
rect 430672 148854 430724 148860
rect 442264 148912 442316 148918
rect 442264 148854 442316 148860
rect 447232 148912 447284 148918
rect 447232 148854 447284 148860
rect 457732 148850 457760 151028
rect 468588 148850 468616 172518
rect 475396 170898 475424 172722
rect 484400 172712 484452 172718
rect 484400 172654 484452 172660
rect 475042 170870 475424 170898
rect 484412 170898 484440 172654
rect 494520 172644 494572 172650
rect 494520 172586 494572 172592
rect 494060 172576 494112 172582
rect 494060 172518 494112 172524
rect 494072 170898 494100 172518
rect 484412 170870 484702 170898
rect 494072 170870 494362 170898
rect 473266 160712 473322 160721
rect 473266 160647 473322 160656
rect 469218 160168 469274 160177
rect 469218 160103 469274 160112
rect 469232 151706 469260 160103
rect 473280 151706 473308 160647
rect 494532 151722 494560 172586
rect 469220 151700 469272 151706
rect 469220 151642 469272 151648
rect 473268 151700 473320 151706
rect 494362 151694 494560 151722
rect 473268 151642 473320 151648
rect 475028 148918 475056 151028
rect 484688 148918 484716 151028
rect 494716 149054 494744 172722
rect 511356 172644 511408 172650
rect 511356 172586 511408 172592
rect 522304 172644 522356 172650
rect 522304 172586 522356 172592
rect 496084 172576 496136 172582
rect 496084 172518 496136 172524
rect 494704 149048 494756 149054
rect 494704 148990 494756 148996
rect 496096 148918 496124 172518
rect 511368 170898 511396 172586
rect 520924 172576 520976 172582
rect 520924 172518 520976 172524
rect 520936 170898 520964 172518
rect 511368 170870 511658 170898
rect 520936 170870 521318 170898
rect 501064 170326 501998 170354
rect 500866 161256 500922 161265
rect 500866 161191 500922 161200
rect 496818 160576 496874 160585
rect 496818 160511 496874 160520
rect 496832 151774 496860 160511
rect 500880 151774 500908 161191
rect 496820 151768 496872 151774
rect 496820 151710 496872 151716
rect 500868 151768 500920 151774
rect 500868 151710 500920 151716
rect 501064 148918 501092 170326
rect 522316 151814 522344 172586
rect 522396 172576 522448 172582
rect 522396 172518 522448 172524
rect 521856 151786 522344 151814
rect 521856 151722 521884 151786
rect 521410 151694 521884 151722
rect 501984 149054 502012 151028
rect 501972 149048 502024 149054
rect 501972 148990 502024 148996
rect 475016 148912 475068 148918
rect 475016 148854 475068 148860
rect 484676 148912 484728 148918
rect 484676 148854 484728 148860
rect 496084 148912 496136 148918
rect 496084 148854 496136 148860
rect 501052 148912 501104 148918
rect 501052 148854 501104 148860
rect 511736 148850 511764 151028
rect 522408 148850 522436 172518
rect 528664 170898 528692 173130
rect 538404 172644 538456 172650
rect 538404 172586 538456 172592
rect 538416 170898 538444 172586
rect 547972 172576 548024 172582
rect 547972 172518 548024 172524
rect 547984 170898 548012 172518
rect 528664 170870 529046 170898
rect 538416 170870 538706 170898
rect 547984 170870 548366 170898
rect 526444 170400 526496 170406
rect 526444 170342 526496 170348
rect 526456 161401 526484 170342
rect 526442 161392 526498 161401
rect 526442 161327 526498 161336
rect 523038 160576 523094 160585
rect 523038 160511 523094 160520
rect 550638 160576 550694 160585
rect 550638 160511 550694 160520
rect 523052 151706 523080 160511
rect 550652 151774 550680 160511
rect 550640 151768 550692 151774
rect 550640 151710 550692 151716
rect 523040 151700 523092 151706
rect 523040 151642 523092 151648
rect 529032 148918 529060 151028
rect 529020 148912 529072 148918
rect 529020 148854 529072 148860
rect 150992 148844 151044 148850
rect 150992 148786 151044 148792
rect 160652 148844 160704 148850
rect 160652 148786 160704 148792
rect 171784 148844 171836 148850
rect 171784 148786 171836 148792
rect 214656 148844 214708 148850
rect 214656 148786 214708 148792
rect 225604 148844 225656 148850
rect 225604 148786 225656 148792
rect 268660 148844 268712 148850
rect 268660 148786 268712 148792
rect 279516 148844 279568 148850
rect 279516 148786 279568 148792
rect 285772 148844 285824 148850
rect 285772 148786 285824 148792
rect 295708 148844 295760 148850
rect 295708 148786 295760 148792
rect 307024 148844 307076 148850
rect 307024 148786 307076 148792
rect 311992 148844 312044 148850
rect 311992 148786 312044 148792
rect 322664 148844 322716 148850
rect 322664 148786 322716 148792
rect 333244 148844 333296 148850
rect 333244 148786 333296 148792
rect 339592 148844 339644 148850
rect 339592 148786 339644 148792
rect 349712 148844 349764 148850
rect 349712 148786 349764 148792
rect 359556 148844 359608 148850
rect 359556 148786 359608 148792
rect 365812 148844 365864 148850
rect 365812 148786 365864 148792
rect 376668 148844 376720 148850
rect 376668 148786 376720 148792
rect 387064 148844 387116 148850
rect 387064 148786 387116 148792
rect 393412 148844 393464 148850
rect 393412 148786 393464 148792
rect 403716 148844 403768 148850
rect 403716 148786 403768 148792
rect 414664 148844 414716 148850
rect 414664 148786 414716 148792
rect 457720 148844 457772 148850
rect 457720 148786 457772 148792
rect 468576 148844 468628 148850
rect 468576 148786 468628 148792
rect 511724 148844 511776 148850
rect 511724 148786 511776 148792
rect 522396 148844 522448 148850
rect 522396 148786 522448 148792
rect 538692 148782 538720 151028
rect 548352 148986 548380 151028
rect 548340 148980 548392 148986
rect 548340 148922 548392 148928
rect 538680 148776 538732 148782
rect 538680 148718 538732 148724
rect 529020 146940 529072 146946
rect 529020 146882 529072 146888
rect 149704 146600 149756 146606
rect 149704 146542 149756 146548
rect 148966 134192 149022 134201
rect 148966 134127 149022 134136
rect 148980 125594 149008 134127
rect 148968 125588 149020 125594
rect 148968 125530 149020 125536
rect 123668 122732 123720 122738
rect 123668 122674 123720 122680
rect 133788 122732 133840 122738
rect 133788 122674 133840 122680
rect 144276 122732 144328 122738
rect 144276 122674 144328 122680
rect 146944 122732 146996 122738
rect 146944 122674 146996 122680
rect 79968 122664 80020 122670
rect 79968 122606 80020 122612
rect 90364 122664 90416 122670
rect 90364 122606 90416 122612
rect 106556 122664 106608 122670
rect 106556 122606 106608 122612
rect 116584 122664 116636 122670
rect 116584 122606 116636 122612
rect 122932 122664 122984 122670
rect 122932 122606 122984 122612
rect 146944 118992 146996 118998
rect 146944 118934 146996 118940
rect 52460 118924 52512 118930
rect 52460 118866 52512 118872
rect 43352 118720 43404 118726
rect 43352 118662 43404 118668
rect 43364 116906 43392 118662
rect 43102 116878 43392 116906
rect 52472 116906 52500 118866
rect 62488 118856 62540 118862
rect 62488 118798 62540 118804
rect 79324 118856 79376 118862
rect 79324 118798 79376 118804
rect 90456 118856 90508 118862
rect 90456 118798 90508 118804
rect 106372 118856 106424 118862
rect 106372 118798 106424 118804
rect 116492 118856 116544 118862
rect 116492 118798 116544 118804
rect 133420 118856 133472 118862
rect 133420 118798 133472 118804
rect 62120 118788 62172 118794
rect 62120 118730 62172 118736
rect 62132 116906 62160 118730
rect 52472 116878 52670 116906
rect 62132 116878 62330 116906
rect 37924 116612 37976 116618
rect 37924 116554 37976 116560
rect 41326 107264 41382 107273
rect 41326 107199 41382 107208
rect 37922 106584 37978 106593
rect 37922 106519 37978 106528
rect 36820 97708 36872 97714
rect 36820 97650 36872 97656
rect 36820 91180 36872 91186
rect 36820 91122 36872 91128
rect 36832 68882 36860 91122
rect 37936 90370 37964 106519
rect 41340 97918 41368 107199
rect 41328 97912 41380 97918
rect 41328 97854 41380 97860
rect 62500 97730 62528 118798
rect 64144 118788 64196 118794
rect 64144 118730 64196 118736
rect 62764 118720 62816 118726
rect 62764 118662 62816 118668
rect 62422 97702 62528 97730
rect 42996 95130 43024 97036
rect 52748 95130 52776 97036
rect 62776 95198 62804 118662
rect 62764 95192 62816 95198
rect 62764 95134 62816 95140
rect 64156 95130 64184 118730
rect 79336 116906 79364 118798
rect 89076 118788 89128 118794
rect 89076 118730 89128 118736
rect 90364 118788 90416 118794
rect 90364 118730 90416 118736
rect 89088 116906 89116 118730
rect 79336 116878 79718 116906
rect 89088 116878 89378 116906
rect 69124 116334 70058 116362
rect 68926 106720 68982 106729
rect 68926 106655 68982 106664
rect 64878 106584 64934 106593
rect 64878 106519 64934 106528
rect 64892 97986 64920 106519
rect 64880 97980 64932 97986
rect 64880 97922 64932 97928
rect 68940 97850 68968 106655
rect 68928 97844 68980 97850
rect 68928 97786 68980 97792
rect 69124 95130 69152 116334
rect 89720 100292 89772 100298
rect 89720 100234 89772 100240
rect 89732 97730 89760 100234
rect 89378 97702 89760 97730
rect 70044 95198 70072 97036
rect 70032 95192 70084 95198
rect 70032 95134 70084 95140
rect 42984 95124 43036 95130
rect 42984 95066 43036 95072
rect 52736 95124 52788 95130
rect 52736 95066 52788 95072
rect 64144 95124 64196 95130
rect 64144 95066 64196 95072
rect 69112 95124 69164 95130
rect 69112 95066 69164 95072
rect 79704 95062 79732 97036
rect 90376 95062 90404 118730
rect 90468 100298 90496 118798
rect 106384 116906 106412 118798
rect 115940 118788 115992 118794
rect 115940 118730 115992 118736
rect 115952 116906 115980 118730
rect 106384 116878 106674 116906
rect 115952 116878 116334 116906
rect 96724 116334 97014 116362
rect 95146 107264 95202 107273
rect 95146 107199 95202 107208
rect 91098 106584 91154 106593
rect 91098 106519 91154 106528
rect 90456 100292 90508 100298
rect 90456 100234 90508 100240
rect 91112 97918 91140 106519
rect 95160 97986 95188 107199
rect 95148 97980 95200 97986
rect 95148 97922 95200 97928
rect 91100 97912 91152 97918
rect 91100 97854 91152 97860
rect 96724 95198 96752 116334
rect 96712 95192 96764 95198
rect 96712 95134 96764 95140
rect 97000 95130 97028 97036
rect 96988 95124 97040 95130
rect 96988 95066 97040 95072
rect 106660 95062 106688 97036
rect 116320 96914 116348 97036
rect 116504 96914 116532 118798
rect 116584 118788 116636 118794
rect 116584 118730 116636 118736
rect 116320 96886 116532 96914
rect 116596 95062 116624 118730
rect 133432 116906 133460 118798
rect 142988 118788 143040 118794
rect 142988 118730 143040 118736
rect 144184 118788 144236 118794
rect 144184 118730 144236 118736
rect 143000 116906 143028 118730
rect 133432 116878 133722 116906
rect 143000 116878 143382 116906
rect 122944 116334 124062 116362
rect 122746 107264 122802 107273
rect 122746 107199 122802 107208
rect 118698 106584 118754 106593
rect 118698 106519 118754 106528
rect 118712 97850 118740 106519
rect 122760 97918 122788 107199
rect 122748 97912 122800 97918
rect 122748 97854 122800 97860
rect 118700 97844 118752 97850
rect 118700 97786 118752 97792
rect 79692 95056 79744 95062
rect 79692 94998 79744 95004
rect 90364 95056 90416 95062
rect 90364 94998 90416 95004
rect 106648 95056 106700 95062
rect 106648 94998 106700 95004
rect 116584 95056 116636 95062
rect 116584 94998 116636 95004
rect 122944 94994 122972 116334
rect 143632 100292 143684 100298
rect 143632 100234 143684 100240
rect 143644 97730 143672 100234
rect 143382 97702 143672 97730
rect 124048 95130 124076 97036
rect 124036 95124 124088 95130
rect 124036 95066 124088 95072
rect 133708 95062 133736 97036
rect 144196 95062 144224 118730
rect 144276 118720 144328 118726
rect 144276 118662 144328 118668
rect 144288 100298 144316 118662
rect 146298 106312 146354 106321
rect 146298 106247 146354 106256
rect 144276 100292 144328 100298
rect 144276 100234 144328 100240
rect 146312 97986 146340 106247
rect 146300 97980 146352 97986
rect 146300 97922 146352 97928
rect 133696 95056 133748 95062
rect 133696 94998 133748 95004
rect 144184 95056 144236 95062
rect 144184 94998 144236 95004
rect 122932 94988 122984 94994
rect 122932 94930 122984 94936
rect 52644 91316 52696 91322
rect 52644 91258 52696 91264
rect 43076 91248 43128 91254
rect 43076 91190 43128 91196
rect 37924 90364 37976 90370
rect 37924 90306 37976 90312
rect 43088 89964 43116 91190
rect 52656 89964 52684 91258
rect 62764 91248 62816 91254
rect 62764 91190 62816 91196
rect 90456 91248 90508 91254
rect 90456 91190 90508 91196
rect 106648 91248 106700 91254
rect 106648 91190 106700 91196
rect 116492 91248 116544 91254
rect 116492 91190 116544 91196
rect 133696 91248 133748 91254
rect 133696 91190 133748 91196
rect 144276 91248 144328 91254
rect 144276 91190 144328 91196
rect 62304 91180 62356 91186
rect 62304 91122 62356 91128
rect 62316 89964 62344 91122
rect 62488 91112 62540 91118
rect 62488 91054 62540 91060
rect 41328 88460 41380 88466
rect 41328 88402 41380 88408
rect 41340 80345 41368 88402
rect 41326 80336 41382 80345
rect 41326 80271 41382 80280
rect 37922 78976 37978 78985
rect 37922 78911 37978 78920
rect 36820 68876 36872 68882
rect 36820 68818 36872 68824
rect 36728 68740 36780 68746
rect 36728 68682 36780 68688
rect 36728 65136 36780 65142
rect 36728 65078 36780 65084
rect 36740 44062 36768 65078
rect 36820 65000 36872 65006
rect 36820 64942 36872 64948
rect 36728 44056 36780 44062
rect 36728 43998 36780 44004
rect 36832 41274 36860 64942
rect 37936 62830 37964 78911
rect 62500 70666 62528 91054
rect 62422 70638 62528 70666
rect 42812 70094 43010 70122
rect 52762 70094 53144 70122
rect 42812 68950 42840 70094
rect 53116 69018 53144 70094
rect 53104 69012 53156 69018
rect 53104 68954 53156 68960
rect 62776 68950 62804 91190
rect 64144 91180 64196 91186
rect 64144 91122 64196 91128
rect 89352 91180 89404 91186
rect 89352 91122 89404 91128
rect 90364 91180 90416 91186
rect 90364 91122 90416 91128
rect 64156 69018 64184 91122
rect 79692 91112 79744 91118
rect 79692 91054 79744 91060
rect 79704 89964 79732 91054
rect 89364 89964 89392 91122
rect 69124 89270 70058 89298
rect 68928 88528 68980 88534
rect 68928 88470 68980 88476
rect 64880 88392 64932 88398
rect 64880 88334 64932 88340
rect 64892 79665 64920 88334
rect 68940 80889 68968 88470
rect 68926 80880 68982 80889
rect 68926 80815 68982 80824
rect 64878 79656 64934 79665
rect 64878 79591 64934 79600
rect 69124 69018 69152 89270
rect 89720 72344 89772 72350
rect 89720 72286 89772 72292
rect 89732 70666 89760 72286
rect 89378 70638 89760 70666
rect 69768 70094 70058 70122
rect 79718 70094 80008 70122
rect 64144 69012 64196 69018
rect 64144 68954 64196 68960
rect 69112 69012 69164 69018
rect 69112 68954 69164 68960
rect 69768 68950 69796 70094
rect 42800 68944 42852 68950
rect 42800 68886 42852 68892
rect 62764 68944 62816 68950
rect 62764 68886 62816 68892
rect 69756 68944 69808 68950
rect 69756 68886 69808 68892
rect 79980 68882 80008 70094
rect 90376 68882 90404 91122
rect 90468 72350 90496 91190
rect 106660 89964 106688 91190
rect 116308 91180 116360 91186
rect 116308 91122 116360 91128
rect 116320 89964 116348 91122
rect 96724 89270 97014 89298
rect 91100 88460 91152 88466
rect 91100 88402 91152 88408
rect 91112 79665 91140 88402
rect 95148 88392 95200 88398
rect 95148 88334 95200 88340
rect 95160 80345 95188 88334
rect 95146 80336 95202 80345
rect 95146 80271 95202 80280
rect 91098 79656 91154 79665
rect 91098 79591 91154 79600
rect 90456 72344 90508 72350
rect 90456 72286 90508 72292
rect 96724 69018 96752 89270
rect 116228 70650 116334 70666
rect 116504 70650 116532 91190
rect 116584 91180 116636 91186
rect 116584 91122 116636 91128
rect 116216 70644 116334 70650
rect 116268 70638 116334 70644
rect 116492 70644 116544 70650
rect 116216 70586 116268 70592
rect 116492 70586 116544 70592
rect 96816 70094 97014 70122
rect 106568 70094 106674 70122
rect 96712 69012 96764 69018
rect 96712 68954 96764 68960
rect 96816 68950 96844 70094
rect 96804 68944 96856 68950
rect 96804 68886 96856 68892
rect 106568 68882 106596 70094
rect 116596 68882 116624 91122
rect 133708 89964 133736 91190
rect 143356 91180 143408 91186
rect 143356 91122 143408 91128
rect 144184 91180 144236 91186
rect 144184 91122 144236 91128
rect 143368 89964 143396 91122
rect 122944 89270 124062 89298
rect 118700 88528 118752 88534
rect 118700 88470 118752 88476
rect 118712 79665 118740 88470
rect 122748 88460 122800 88466
rect 122748 88402 122800 88408
rect 122760 80345 122788 88402
rect 122746 80336 122802 80345
rect 122746 80271 122802 80280
rect 118698 79656 118754 79665
rect 118698 79591 118754 79600
rect 122944 68882 122972 89270
rect 143632 72344 143684 72350
rect 143632 72286 143684 72292
rect 143644 70666 143672 72286
rect 143382 70638 143672 70666
rect 123680 70094 124062 70122
rect 133722 70094 133828 70122
rect 123680 68950 123708 70094
rect 133800 68950 133828 70094
rect 144196 68950 144224 91122
rect 144288 72350 144316 91190
rect 146300 88392 146352 88398
rect 146300 88334 146352 88340
rect 146312 80073 146340 88334
rect 146298 80064 146354 80073
rect 146298 79999 146354 80008
rect 144276 72344 144328 72350
rect 144276 72286 144328 72292
rect 146956 69018 146984 118934
rect 148966 107264 149022 107273
rect 148966 107199 149022 107208
rect 148980 97986 149008 107199
rect 148968 97980 149020 97986
rect 148968 97922 149020 97928
rect 149716 95130 149744 146542
rect 232044 146532 232096 146538
rect 232044 146474 232096 146480
rect 251824 146532 251876 146538
rect 251824 146474 251876 146480
rect 475016 146532 475068 146538
rect 475016 146474 475068 146480
rect 494704 146532 494756 146538
rect 494704 146474 494756 146480
rect 160652 146464 160704 146470
rect 160652 146406 160704 146412
rect 170496 146464 170548 146470
rect 170496 146406 170548 146412
rect 187700 146464 187752 146470
rect 187700 146406 187752 146412
rect 197452 146464 197504 146470
rect 197452 146406 197504 146412
rect 214656 146464 214708 146470
rect 214656 146406 214708 146412
rect 224500 146464 224552 146470
rect 224500 146406 224552 146412
rect 160664 143956 160692 146406
rect 170312 146396 170364 146402
rect 170312 146338 170364 146344
rect 170324 143956 170352 146338
rect 150544 143262 151018 143290
rect 150544 122670 150572 143262
rect 170232 124642 170338 124658
rect 170508 124642 170536 146406
rect 178040 146396 178092 146402
rect 178040 146338 178092 146344
rect 171784 146328 171836 146334
rect 171784 146270 171836 146276
rect 170220 124636 170338 124642
rect 170272 124630 170338 124636
rect 170496 124636 170548 124642
rect 170220 124578 170272 124584
rect 170496 124578 170548 124584
rect 150728 124086 151018 124114
rect 160572 124086 160678 124114
rect 150532 122664 150584 122670
rect 150532 122606 150584 122612
rect 150728 122602 150756 124086
rect 160572 122602 160600 124086
rect 171796 122602 171824 146270
rect 178052 143956 178080 146338
rect 187712 143956 187740 146406
rect 197360 146328 197412 146334
rect 197360 146270 197412 146276
rect 197372 143956 197400 146270
rect 176566 133920 176622 133929
rect 176566 133855 176622 133864
rect 172518 133512 172574 133521
rect 172518 133447 172574 133456
rect 172532 125526 172560 133447
rect 176580 125526 176608 133855
rect 172520 125520 172572 125526
rect 172520 125462 172572 125468
rect 176568 125520 176620 125526
rect 176568 125462 176620 125468
rect 197464 124794 197492 146406
rect 200764 146396 200816 146402
rect 200764 146338 200816 146344
rect 199384 146328 199436 146334
rect 199384 146270 199436 146276
rect 197386 124766 197492 124794
rect 178066 124086 178172 124114
rect 187726 124086 188016 124114
rect 178144 122670 178172 124086
rect 187988 122670 188016 124086
rect 199396 122670 199424 146270
rect 200118 133512 200174 133521
rect 200118 133447 200174 133456
rect 200132 125594 200160 133447
rect 200120 125588 200172 125594
rect 200120 125530 200172 125536
rect 200776 122806 200804 146338
rect 214668 143956 214696 146406
rect 224316 146328 224368 146334
rect 224316 146270 224368 146276
rect 224328 143956 224356 146270
rect 204364 143262 205022 143290
rect 202786 134192 202842 134201
rect 202786 134127 202842 134136
rect 202800 125594 202828 134127
rect 202788 125588 202840 125594
rect 202788 125530 202840 125536
rect 200764 122800 200816 122806
rect 200764 122742 200816 122748
rect 204364 122670 204392 143262
rect 224512 124794 224540 146406
rect 225604 146328 225656 146334
rect 225604 146270 225656 146276
rect 224342 124766 224540 124794
rect 204640 124086 205022 124114
rect 214682 124086 215064 124114
rect 204640 122806 204668 124086
rect 204628 122800 204680 122806
rect 204628 122742 204680 122748
rect 178132 122664 178184 122670
rect 178132 122606 178184 122612
rect 187976 122664 188028 122670
rect 187976 122606 188028 122612
rect 199384 122664 199436 122670
rect 199384 122606 199436 122612
rect 204352 122664 204404 122670
rect 204352 122606 204404 122612
rect 215036 122602 215064 124086
rect 225616 122602 225644 146270
rect 232056 143956 232084 146474
rect 241704 146464 241756 146470
rect 241704 146406 241756 146412
rect 241716 143956 241744 146406
rect 251456 146396 251508 146402
rect 251456 146338 251508 146344
rect 251364 146328 251416 146334
rect 251364 146270 251416 146276
rect 251376 143956 251404 146270
rect 230386 134192 230442 134201
rect 230386 134127 230442 134136
rect 226338 133512 226394 133521
rect 226338 133447 226394 133456
rect 226352 125526 226380 133447
rect 230400 125526 230428 134127
rect 226340 125520 226392 125526
rect 226340 125462 226392 125468
rect 230388 125520 230440 125526
rect 230388 125462 230440 125468
rect 251468 124794 251496 146338
rect 251390 124766 251496 124794
rect 231964 124086 232070 124114
rect 241730 124086 242112 124114
rect 231964 122670 231992 124086
rect 242084 122670 242112 124086
rect 251836 122806 251864 146474
rect 413468 146464 413520 146470
rect 413468 146406 413520 146412
rect 430672 146464 430724 146470
rect 430672 146406 430724 146412
rect 440516 146464 440568 146470
rect 440516 146406 440568 146412
rect 457628 146464 457680 146470
rect 457628 146406 457680 146412
rect 468484 146464 468536 146470
rect 468484 146406 468536 146412
rect 268660 146396 268712 146402
rect 268660 146338 268712 146344
rect 279516 146396 279568 146402
rect 279516 146338 279568 146344
rect 295708 146396 295760 146402
rect 295708 146338 295760 146344
rect 305460 146396 305512 146402
rect 305460 146338 305512 146344
rect 322664 146396 322716 146402
rect 322664 146338 322716 146344
rect 336004 146396 336056 146402
rect 336004 146338 336056 146344
rect 349712 146396 349764 146402
rect 349712 146338 349764 146344
rect 359464 146396 359516 146402
rect 359464 146338 359516 146344
rect 376668 146396 376720 146402
rect 376668 146338 376720 146344
rect 386512 146396 386564 146402
rect 386512 146338 386564 146344
rect 403624 146396 403676 146402
rect 403624 146338 403676 146344
rect 253204 146328 253256 146334
rect 253204 146270 253256 146276
rect 251824 122800 251876 122806
rect 251824 122742 251876 122748
rect 253216 122670 253244 146270
rect 268672 143956 268700 146338
rect 278320 146328 278372 146334
rect 278320 146270 278372 146276
rect 279424 146328 279476 146334
rect 279424 146270 279476 146276
rect 278332 143956 278360 146270
rect 258184 143262 259026 143290
rect 256606 134192 256662 134201
rect 256606 134127 256662 134136
rect 253938 132968 253994 132977
rect 253938 132903 253994 132912
rect 253952 125594 253980 132903
rect 256620 125594 256648 134127
rect 253940 125588 253992 125594
rect 253940 125530 253992 125536
rect 256608 125588 256660 125594
rect 256608 125530 256660 125536
rect 258184 122670 258212 143262
rect 278688 125520 278740 125526
rect 278688 125462 278740 125468
rect 278700 124794 278728 125462
rect 278346 124766 278728 124794
rect 258736 124086 259026 124114
rect 268686 124086 268976 124114
rect 258736 122806 258764 124086
rect 258724 122800 258776 122806
rect 258724 122742 258776 122748
rect 231952 122664 232004 122670
rect 231952 122606 232004 122612
rect 242072 122664 242124 122670
rect 242072 122606 242124 122612
rect 253204 122664 253256 122670
rect 253204 122606 253256 122612
rect 258172 122664 258224 122670
rect 258172 122606 258224 122612
rect 268948 122602 268976 124086
rect 279436 122602 279464 146270
rect 279528 125526 279556 146338
rect 285784 144078 286088 144106
rect 284206 133920 284262 133929
rect 284206 133855 284262 133864
rect 280158 133512 280214 133521
rect 280158 133447 280214 133456
rect 279516 125520 279568 125526
rect 279516 125462 279568 125468
rect 280172 125458 280200 133447
rect 284220 125526 284248 133855
rect 284208 125520 284260 125526
rect 284208 125462 284260 125468
rect 280160 125452 280212 125458
rect 280160 125394 280212 125400
rect 285784 122670 285812 144078
rect 286060 143956 286088 144078
rect 295720 143956 295748 146338
rect 305368 146328 305420 146334
rect 305368 146270 305420 146276
rect 305380 143956 305408 146270
rect 305472 124794 305500 146338
rect 307024 146328 307076 146334
rect 307024 146270 307076 146276
rect 305394 124766 305500 124794
rect 286074 124086 286180 124114
rect 295734 124086 296024 124114
rect 285772 122664 285824 122670
rect 285772 122606 285824 122612
rect 286152 122602 286180 124086
rect 295996 122602 296024 124086
rect 307036 122602 307064 146270
rect 322676 143956 322704 146338
rect 332324 146328 332376 146334
rect 332324 146270 332376 146276
rect 333244 146328 333296 146334
rect 333244 146270 333296 146276
rect 332336 143956 332364 146270
rect 312004 143262 313030 143290
rect 311806 134192 311862 134201
rect 311806 134127 311862 134136
rect 307758 133512 307814 133521
rect 307758 133447 307814 133456
rect 307772 125594 307800 133447
rect 307760 125588 307812 125594
rect 307760 125530 307812 125536
rect 311820 125458 311848 134127
rect 311808 125452 311860 125458
rect 311808 125394 311860 125400
rect 312004 122602 312032 143262
rect 312648 124086 313030 124114
rect 322690 124086 322888 124114
rect 332350 124086 332548 124114
rect 312648 122670 312676 124086
rect 312636 122664 312688 122670
rect 312636 122606 312688 122612
rect 322860 122602 322888 124086
rect 332520 122806 332548 124086
rect 332508 122800 332560 122806
rect 332508 122742 332560 122748
rect 333256 122602 333284 146270
rect 335358 133512 335414 133521
rect 335358 133447 335414 133456
rect 335372 125526 335400 133447
rect 335360 125520 335412 125526
rect 335360 125462 335412 125468
rect 336016 122806 336044 146338
rect 339604 144078 340092 144106
rect 338026 134192 338082 134201
rect 338026 134127 338082 134136
rect 338040 125594 338068 134127
rect 338028 125588 338080 125594
rect 338028 125530 338080 125536
rect 336004 122800 336056 122806
rect 336004 122742 336056 122748
rect 339604 122670 339632 144078
rect 340064 143956 340092 144078
rect 349724 143956 349752 146338
rect 359372 146328 359424 146334
rect 359372 146270 359424 146276
rect 359384 143956 359412 146270
rect 359476 124794 359504 146338
rect 359556 146328 359608 146334
rect 359556 146270 359608 146276
rect 359398 124766 359504 124794
rect 340078 124086 340184 124114
rect 349738 124086 350120 124114
rect 339592 122664 339644 122670
rect 339592 122606 339644 122612
rect 340156 122602 340184 124086
rect 350092 122602 350120 124086
rect 359568 122602 359596 146270
rect 376680 143956 376708 146338
rect 386328 146328 386380 146334
rect 386328 146270 386380 146276
rect 386340 143956 386368 146270
rect 365824 143262 367034 143290
rect 365626 134192 365682 134201
rect 365626 134127 365682 134136
rect 361578 132968 361634 132977
rect 361578 132903 361634 132912
rect 361592 125458 361620 132903
rect 365640 125526 365668 134127
rect 365628 125520 365680 125526
rect 365628 125462 365680 125468
rect 361580 125452 361632 125458
rect 361580 125394 361632 125400
rect 365824 122602 365852 143262
rect 386524 124794 386552 146338
rect 387064 146328 387116 146334
rect 387064 146270 387116 146276
rect 386354 124766 386552 124794
rect 366744 124086 367034 124114
rect 376588 124086 376694 124114
rect 366744 122670 366772 124086
rect 366732 122664 366784 122670
rect 366732 122606 366784 122612
rect 376588 122602 376616 124086
rect 387076 122602 387104 146270
rect 403636 143956 403664 146338
rect 413284 146328 413336 146334
rect 413284 146270 413336 146276
rect 413296 143956 413324 146270
rect 393424 143262 393990 143290
rect 391846 133920 391902 133929
rect 391846 133855 391902 133864
rect 389178 133512 389234 133521
rect 389178 133447 389234 133456
rect 389192 125594 389220 133447
rect 391860 125594 391888 133855
rect 389180 125588 389232 125594
rect 389180 125530 389232 125536
rect 391848 125588 391900 125594
rect 391848 125530 391900 125536
rect 393424 122602 393452 143262
rect 413480 124794 413508 146406
rect 421012 146396 421064 146402
rect 421012 146338 421064 146344
rect 414664 146328 414716 146334
rect 414664 146270 414716 146276
rect 413402 124766 413508 124794
rect 393608 124086 393990 124114
rect 403742 124086 404032 124114
rect 393608 122670 393636 124086
rect 393596 122664 393648 122670
rect 393596 122606 393648 122612
rect 404004 122602 404032 124086
rect 414676 122602 414704 146270
rect 421024 143956 421052 146338
rect 430684 143956 430712 146406
rect 440332 146328 440384 146334
rect 440332 146270 440384 146276
rect 440344 143956 440372 146270
rect 419446 134192 419502 134201
rect 419446 134127 419502 134136
rect 415398 133512 415454 133521
rect 415398 133447 415454 133456
rect 415412 125526 415440 133447
rect 419460 125526 419488 134127
rect 415400 125520 415452 125526
rect 415400 125462 415452 125468
rect 419448 125520 419500 125526
rect 419448 125462 419500 125468
rect 440528 124794 440556 146406
rect 445024 146396 445076 146402
rect 445024 146338 445076 146344
rect 442264 146328 442316 146334
rect 442264 146270 442316 146276
rect 440358 124766 440556 124794
rect 420932 124086 421038 124114
rect 430698 124086 431080 124114
rect 420932 122670 420960 124086
rect 431052 122670 431080 124086
rect 442276 122670 442304 146270
rect 442998 133512 443054 133521
rect 442998 133447 443054 133456
rect 443012 125594 443040 133447
rect 443000 125588 443052 125594
rect 443000 125530 443052 125536
rect 445036 125458 445064 146338
rect 457640 143956 457668 146406
rect 467288 146328 467340 146334
rect 467288 146270 467340 146276
rect 467300 143956 467328 146270
rect 447244 143262 447994 143290
rect 445666 134192 445722 134201
rect 445666 134127 445722 134136
rect 445680 125594 445708 134127
rect 445668 125588 445720 125594
rect 445668 125530 445720 125536
rect 445024 125452 445076 125458
rect 445024 125394 445076 125400
rect 447244 122670 447272 143262
rect 468496 132494 468524 146406
rect 468576 146328 468628 146334
rect 468576 146270 468628 146276
rect 467852 132466 468524 132494
rect 447692 125452 447744 125458
rect 447692 125394 447744 125400
rect 447704 124794 447732 125394
rect 467852 124930 467880 132466
rect 467760 124902 467880 124930
rect 467760 124794 467788 124902
rect 447704 124766 447994 124794
rect 467406 124766 467788 124794
rect 457746 124086 458128 124114
rect 420920 122664 420972 122670
rect 420920 122606 420972 122612
rect 431040 122664 431092 122670
rect 431040 122606 431092 122612
rect 442264 122664 442316 122670
rect 442264 122606 442316 122612
rect 447232 122664 447284 122670
rect 447232 122606 447284 122612
rect 458100 122602 458128 124086
rect 468588 122602 468616 146270
rect 475028 143956 475056 146474
rect 484676 146464 484728 146470
rect 484676 146406 484728 146412
rect 484688 143956 484716 146406
rect 494520 146396 494572 146402
rect 494520 146338 494572 146344
rect 494336 146328 494388 146334
rect 494336 146270 494388 146276
rect 494348 143956 494376 146270
rect 473266 133920 473322 133929
rect 473266 133855 473322 133864
rect 469218 132968 469274 132977
rect 469218 132903 469274 132912
rect 469232 125526 469260 132903
rect 473280 125526 473308 133855
rect 469220 125520 469272 125526
rect 469220 125462 469272 125468
rect 473268 125520 473320 125526
rect 473268 125462 473320 125468
rect 494532 124794 494560 146338
rect 494362 124766 494560 124794
rect 474752 124086 475042 124114
rect 484702 124086 484992 124114
rect 474752 122670 474780 124086
rect 484964 122670 484992 124086
rect 494716 122806 494744 146474
rect 511632 146396 511684 146402
rect 511632 146338 511684 146344
rect 522396 146396 522448 146402
rect 522396 146338 522448 146344
rect 496084 146328 496136 146334
rect 496084 146270 496136 146276
rect 494704 122800 494756 122806
rect 494704 122742 494756 122748
rect 496096 122670 496124 146270
rect 511644 143956 511672 146338
rect 521292 146328 521344 146334
rect 521292 146270 521344 146276
rect 522304 146328 522356 146334
rect 522304 146270 522356 146276
rect 521304 143956 521332 146270
rect 501064 143262 501998 143290
rect 500866 134192 500922 134201
rect 500866 134127 500922 134136
rect 496818 133512 496874 133521
rect 496818 133447 496874 133456
rect 496832 125594 496860 133447
rect 500880 125594 500908 134127
rect 496820 125588 496872 125594
rect 496820 125530 496872 125536
rect 500868 125588 500920 125594
rect 500868 125530 500920 125536
rect 501064 122670 501092 143262
rect 501616 124086 501998 124114
rect 511750 124086 511856 124114
rect 521410 124086 521516 124114
rect 501616 122806 501644 124086
rect 501604 122800 501656 122806
rect 501604 122742 501656 122748
rect 474740 122664 474792 122670
rect 474740 122606 474792 122612
rect 484952 122664 485004 122670
rect 484952 122606 485004 122612
rect 496084 122664 496136 122670
rect 496084 122606 496136 122612
rect 501052 122664 501104 122670
rect 501052 122606 501104 122612
rect 511828 122602 511856 124086
rect 521488 122806 521516 124086
rect 521476 122800 521528 122806
rect 521476 122742 521528 122748
rect 522316 122602 522344 146270
rect 522408 122806 522436 146338
rect 526444 144220 526496 144226
rect 526444 144162 526496 144168
rect 526456 134337 526484 144162
rect 529032 143956 529060 146882
rect 538680 146396 538732 146402
rect 538680 146338 538732 146344
rect 538692 143956 538720 146338
rect 548340 146328 548392 146334
rect 548340 146270 548392 146276
rect 548352 143956 548380 146270
rect 526442 134328 526498 134337
rect 526442 134263 526498 134272
rect 523038 133512 523094 133521
rect 523038 133447 523094 133456
rect 523052 125526 523080 133447
rect 550638 132968 550694 132977
rect 550638 132903 550694 132912
rect 550652 125594 550680 132903
rect 550640 125588 550692 125594
rect 550640 125530 550692 125536
rect 523040 125520 523092 125526
rect 523040 125462 523092 125468
rect 528664 124086 529046 124114
rect 538416 124086 538706 124114
rect 547984 124086 548366 124114
rect 522396 122800 522448 122806
rect 522396 122742 522448 122748
rect 528664 122670 528692 124086
rect 528652 122664 528704 122670
rect 528652 122606 528704 122612
rect 150716 122596 150768 122602
rect 150716 122538 150768 122544
rect 160560 122596 160612 122602
rect 160560 122538 160612 122544
rect 171784 122596 171836 122602
rect 171784 122538 171836 122544
rect 215024 122596 215076 122602
rect 215024 122538 215076 122544
rect 225604 122596 225656 122602
rect 225604 122538 225656 122544
rect 268936 122596 268988 122602
rect 268936 122538 268988 122544
rect 279424 122596 279476 122602
rect 279424 122538 279476 122544
rect 286140 122596 286192 122602
rect 286140 122538 286192 122544
rect 295984 122596 296036 122602
rect 295984 122538 296036 122544
rect 307024 122596 307076 122602
rect 307024 122538 307076 122544
rect 311992 122596 312044 122602
rect 311992 122538 312044 122544
rect 322848 122596 322900 122602
rect 322848 122538 322900 122544
rect 333244 122596 333296 122602
rect 333244 122538 333296 122544
rect 340144 122596 340196 122602
rect 340144 122538 340196 122544
rect 350080 122596 350132 122602
rect 350080 122538 350132 122544
rect 359556 122596 359608 122602
rect 359556 122538 359608 122544
rect 365812 122596 365864 122602
rect 365812 122538 365864 122544
rect 376576 122596 376628 122602
rect 376576 122538 376628 122544
rect 387064 122596 387116 122602
rect 387064 122538 387116 122544
rect 393412 122596 393464 122602
rect 393412 122538 393464 122544
rect 403992 122596 404044 122602
rect 403992 122538 404044 122544
rect 414664 122596 414716 122602
rect 414664 122538 414716 122544
rect 458088 122596 458140 122602
rect 458088 122538 458140 122544
rect 468576 122596 468628 122602
rect 468576 122538 468628 122544
rect 511816 122596 511868 122602
rect 511816 122538 511868 122544
rect 522304 122596 522356 122602
rect 522304 122538 522356 122544
rect 538416 122534 538444 124086
rect 547984 122738 548012 124086
rect 547972 122732 548024 122738
rect 547972 122674 548024 122680
rect 538404 122528 538456 122534
rect 538404 122470 538456 122476
rect 528744 119400 528796 119406
rect 528744 119342 528796 119348
rect 232320 118924 232372 118930
rect 232320 118866 232372 118872
rect 251824 118924 251876 118930
rect 251824 118866 251876 118872
rect 170496 118856 170548 118862
rect 170496 118798 170548 118804
rect 187792 118856 187844 118862
rect 187792 118798 187844 118804
rect 197544 118856 197596 118862
rect 197544 118798 197596 118804
rect 214380 118856 214432 118862
rect 214380 118798 214432 118804
rect 224500 118856 224552 118862
rect 224500 118798 224552 118804
rect 170036 118788 170088 118794
rect 170036 118730 170088 118736
rect 160284 118720 160336 118726
rect 160284 118662 160336 118668
rect 160296 116906 160324 118662
rect 170048 116906 170076 118730
rect 160296 116878 160678 116906
rect 170048 116878 170338 116906
rect 150544 116334 151018 116362
rect 149704 95124 149756 95130
rect 149704 95066 149756 95072
rect 150544 95062 150572 116334
rect 150532 95056 150584 95062
rect 150532 94998 150584 95004
rect 151004 94994 151032 97036
rect 160664 94994 160692 97036
rect 170324 96914 170352 97036
rect 170508 96914 170536 118798
rect 178408 118788 178460 118794
rect 178408 118730 178460 118736
rect 171784 118720 171836 118726
rect 171784 118662 171836 118668
rect 170324 96886 170536 96914
rect 171796 94994 171824 118662
rect 178420 116906 178448 118730
rect 187804 116906 187832 118798
rect 197452 118720 197504 118726
rect 197452 118662 197504 118668
rect 197464 116906 197492 118662
rect 178066 116878 178448 116906
rect 187726 116878 187832 116906
rect 197386 116878 197492 116906
rect 176566 106720 176622 106729
rect 176566 106655 176622 106664
rect 172518 106584 172574 106593
rect 172518 106519 172574 106528
rect 172532 97918 172560 106519
rect 176580 97918 176608 106655
rect 197556 103514 197584 118798
rect 200764 118788 200816 118794
rect 200764 118730 200816 118736
rect 199384 118720 199436 118726
rect 199384 118662 199436 118668
rect 197464 103486 197584 103514
rect 172520 97912 172572 97918
rect 172520 97854 172572 97860
rect 176568 97912 176620 97918
rect 176568 97854 176620 97860
rect 197464 97730 197492 103486
rect 197386 97702 197492 97730
rect 178052 95062 178080 97036
rect 187712 95062 187740 97036
rect 199396 95062 199424 118662
rect 200118 106584 200174 106593
rect 200118 106519 200174 106528
rect 200132 97986 200160 106519
rect 200120 97980 200172 97986
rect 200120 97922 200172 97928
rect 200776 97850 200804 118730
rect 214392 116906 214420 118798
rect 223948 118720 224000 118726
rect 223948 118662 224000 118668
rect 223960 116906 223988 118662
rect 214392 116878 214682 116906
rect 223960 116878 224342 116906
rect 204364 116334 205022 116362
rect 202786 107264 202842 107273
rect 202786 107199 202842 107208
rect 202800 97986 202828 107199
rect 202788 97980 202840 97986
rect 202788 97922 202840 97928
rect 200764 97844 200816 97850
rect 200764 97786 200816 97792
rect 204364 95062 204392 116334
rect 204628 97844 204680 97850
rect 204628 97786 204680 97792
rect 204640 97730 204668 97786
rect 224512 97730 224540 118798
rect 225604 118720 225656 118726
rect 225604 118662 225656 118668
rect 204640 97702 205022 97730
rect 224342 97702 224540 97730
rect 178040 95056 178092 95062
rect 178040 94998 178092 95004
rect 187700 95056 187752 95062
rect 187700 94998 187752 95004
rect 199384 95056 199436 95062
rect 199384 94998 199436 95004
rect 204352 95056 204404 95062
rect 204352 94998 204404 95004
rect 214668 94994 214696 97036
rect 225616 94994 225644 118662
rect 232332 116906 232360 118866
rect 241520 118856 241572 118862
rect 241520 118798 241572 118804
rect 232070 116878 232360 116906
rect 241532 116906 241560 118798
rect 251456 118788 251508 118794
rect 251456 118730 251508 118736
rect 251180 118720 251232 118726
rect 251180 118662 251232 118668
rect 251192 116906 251220 118662
rect 241532 116878 241730 116906
rect 251192 116878 251390 116906
rect 230386 107264 230442 107273
rect 230386 107199 230442 107208
rect 226338 106584 226394 106593
rect 226338 106519 226394 106528
rect 226352 97918 226380 106519
rect 226340 97912 226392 97918
rect 226340 97854 226392 97860
rect 230400 97850 230428 107199
rect 230388 97844 230440 97850
rect 230388 97786 230440 97792
rect 251468 97730 251496 118730
rect 251390 97702 251496 97730
rect 232056 95062 232084 97036
rect 241716 95062 241744 97036
rect 251836 95198 251864 118866
rect 413468 118856 413520 118862
rect 413468 118798 413520 118804
rect 430580 118856 430632 118862
rect 430580 118798 430632 118804
rect 440516 118856 440568 118862
rect 440516 118798 440568 118804
rect 457260 118856 457312 118862
rect 457260 118798 457312 118804
rect 468576 118856 468628 118862
rect 468576 118798 468628 118804
rect 484400 118856 484452 118862
rect 484400 118798 484452 118804
rect 494520 118856 494572 118862
rect 494520 118798 494572 118804
rect 511356 118856 511408 118862
rect 511356 118798 511408 118804
rect 268292 118788 268344 118794
rect 268292 118730 268344 118736
rect 279424 118788 279476 118794
rect 279424 118730 279476 118736
rect 295800 118788 295852 118794
rect 295800 118730 295852 118736
rect 305644 118788 305696 118794
rect 305644 118730 305696 118736
rect 322388 118788 322440 118794
rect 322388 118730 322440 118736
rect 334624 118788 334676 118794
rect 334624 118730 334676 118736
rect 349804 118788 349856 118794
rect 349804 118730 349856 118736
rect 359556 118788 359608 118794
rect 359556 118730 359608 118736
rect 376300 118788 376352 118794
rect 376300 118730 376352 118736
rect 386512 118788 386564 118794
rect 386512 118730 386564 118736
rect 403348 118788 403400 118794
rect 403348 118730 403400 118736
rect 253204 118720 253256 118726
rect 253204 118662 253256 118668
rect 251824 95192 251876 95198
rect 251824 95134 251876 95140
rect 253216 95062 253244 118662
rect 268304 116906 268332 118730
rect 278044 118720 278096 118726
rect 278044 118662 278096 118668
rect 278056 116906 278084 118662
rect 268304 116878 268686 116906
rect 278056 116878 278346 116906
rect 258184 116334 259026 116362
rect 256606 107264 256662 107273
rect 256606 107199 256662 107208
rect 253938 106312 253994 106321
rect 253938 106247 253994 106256
rect 253952 97986 253980 106247
rect 253940 97980 253992 97986
rect 253940 97922 253992 97928
rect 256620 97918 256648 107199
rect 256608 97912 256660 97918
rect 256608 97854 256660 97860
rect 257988 96688 258040 96694
rect 257988 96630 258040 96636
rect 258000 95198 258028 96630
rect 257988 95192 258040 95198
rect 257988 95134 258040 95140
rect 258184 95062 258212 116334
rect 279436 103514 279464 118730
rect 279516 118720 279568 118726
rect 279516 118662 279568 118668
rect 278792 103486 279464 103514
rect 278792 97730 278820 103486
rect 278346 97702 278820 97730
rect 258736 97022 259026 97050
rect 258736 96694 258764 97022
rect 258724 96688 258776 96694
rect 258724 96630 258776 96636
rect 232044 95056 232096 95062
rect 232044 94998 232096 95004
rect 241704 95056 241756 95062
rect 241704 94998 241756 95004
rect 253204 95056 253256 95062
rect 253204 94998 253256 95004
rect 258172 95056 258224 95062
rect 258172 94998 258224 95004
rect 268672 94994 268700 97036
rect 279528 94994 279556 118662
rect 295812 116906 295840 118730
rect 305552 118720 305604 118726
rect 305552 118662 305604 118668
rect 305564 116906 305592 118662
rect 295734 116878 295840 116906
rect 305394 116878 305592 116906
rect 286074 116470 286180 116498
rect 286152 116414 286180 116470
rect 285772 116408 285824 116414
rect 285772 116350 285824 116356
rect 286140 116408 286192 116414
rect 286140 116350 286192 116356
rect 284206 106720 284262 106729
rect 284206 106655 284262 106664
rect 280158 106584 280214 106593
rect 280158 106519 280214 106528
rect 280172 97850 280200 106519
rect 284220 97986 284248 106655
rect 284208 97980 284260 97986
rect 284208 97922 284260 97928
rect 280160 97844 280212 97850
rect 280160 97786 280212 97792
rect 285784 94994 285812 116350
rect 305656 103514 305684 118730
rect 307024 118720 307076 118726
rect 307024 118662 307076 118668
rect 305472 103486 305684 103514
rect 305472 97730 305500 103486
rect 305394 97702 305500 97730
rect 286060 95062 286088 97036
rect 286048 95056 286100 95062
rect 286048 94998 286100 95004
rect 295720 94994 295748 97036
rect 307036 94994 307064 118662
rect 322400 116906 322428 118730
rect 331956 118720 332008 118726
rect 331956 118662 332008 118668
rect 333244 118720 333296 118726
rect 333244 118662 333296 118668
rect 331968 116906 331996 118662
rect 322400 116878 322690 116906
rect 331968 116878 332350 116906
rect 312004 116334 313030 116362
rect 311806 107264 311862 107273
rect 311806 107199 311862 107208
rect 307758 106584 307814 106593
rect 307758 106519 307814 106528
rect 307772 97918 307800 106519
rect 311820 97918 311848 107199
rect 307760 97912 307812 97918
rect 307760 97854 307812 97860
rect 311808 97912 311860 97918
rect 311808 97854 311860 97860
rect 312004 94994 312032 116334
rect 332508 97844 332560 97850
rect 332508 97786 332560 97792
rect 332520 97730 332548 97786
rect 332350 97702 332548 97730
rect 313016 95062 313044 97036
rect 313004 95056 313056 95062
rect 313004 94998 313056 95004
rect 322676 94994 322704 97036
rect 333256 94994 333284 118662
rect 334636 97850 334664 118730
rect 349816 116906 349844 118730
rect 359464 118720 359516 118726
rect 359464 118662 359516 118668
rect 359476 116906 359504 118662
rect 349738 116878 349844 116906
rect 359398 116878 359504 116906
rect 340078 116346 340184 116362
rect 339592 116340 339644 116346
rect 340078 116340 340196 116346
rect 340078 116334 340144 116340
rect 339592 116282 339644 116288
rect 340144 116282 340196 116288
rect 338026 107264 338082 107273
rect 338026 107199 338082 107208
rect 335358 106584 335414 106593
rect 335358 106519 335414 106528
rect 335372 97986 335400 106519
rect 338040 97986 338068 107199
rect 335360 97980 335412 97986
rect 335360 97922 335412 97928
rect 338028 97980 338080 97986
rect 338028 97922 338080 97928
rect 334624 97844 334676 97850
rect 334624 97786 334676 97792
rect 339604 94994 339632 116282
rect 359568 116090 359596 118730
rect 359740 118720 359792 118726
rect 359740 118662 359792 118668
rect 359476 116062 359596 116090
rect 359476 97730 359504 116062
rect 359752 115818 359780 118662
rect 376312 116906 376340 118730
rect 386052 118720 386104 118726
rect 386052 118662 386104 118668
rect 386064 116906 386092 118662
rect 376312 116878 376694 116906
rect 386064 116878 386354 116906
rect 359398 97702 359504 97730
rect 359568 115790 359780 115818
rect 365824 116334 367034 116362
rect 340064 95062 340092 97036
rect 340052 95056 340104 95062
rect 340052 94998 340104 95004
rect 349724 94994 349752 97036
rect 359568 94994 359596 115790
rect 365626 107264 365682 107273
rect 365626 107199 365682 107208
rect 361578 106312 361634 106321
rect 361578 106247 361634 106256
rect 361592 97918 361620 106247
rect 365640 97918 365668 107199
rect 361580 97912 361632 97918
rect 361580 97854 361632 97860
rect 365628 97912 365680 97918
rect 365628 97854 365680 97860
rect 365824 94994 365852 116334
rect 386524 97730 386552 118730
rect 387064 118720 387116 118726
rect 387064 118662 387116 118668
rect 386354 97702 386552 97730
rect 367020 95062 367048 97036
rect 367008 95056 367060 95062
rect 367008 94998 367060 95004
rect 376680 94994 376708 97036
rect 387076 94994 387104 118662
rect 403360 116906 403388 118730
rect 412916 118720 412968 118726
rect 412916 118662 412968 118668
rect 412928 116906 412956 118662
rect 403360 116878 403650 116906
rect 412928 116878 413310 116906
rect 393424 116334 393990 116362
rect 391846 107264 391902 107273
rect 391846 107199 391902 107208
rect 389178 106584 389234 106593
rect 389178 106519 389234 106528
rect 389192 97986 389220 106519
rect 391860 97986 391888 107199
rect 389180 97980 389232 97986
rect 389180 97922 389232 97928
rect 391848 97980 391900 97986
rect 391848 97922 391900 97928
rect 393424 94994 393452 116334
rect 413480 97730 413508 118798
rect 421288 118788 421340 118794
rect 421288 118730 421340 118736
rect 414664 118720 414716 118726
rect 414664 118662 414716 118668
rect 413402 97702 413508 97730
rect 393976 95062 394004 97036
rect 393964 95056 394016 95062
rect 393964 94998 394016 95004
rect 403728 94994 403756 97036
rect 414676 94994 414704 118662
rect 421300 116906 421328 118730
rect 421038 116878 421328 116906
rect 430592 116906 430620 118798
rect 440240 118720 440292 118726
rect 440240 118662 440292 118668
rect 440252 116906 440280 118662
rect 430592 116878 430698 116906
rect 440252 116878 440358 116906
rect 419446 107264 419502 107273
rect 419446 107199 419502 107208
rect 415398 106584 415454 106593
rect 415398 106519 415454 106528
rect 415412 97918 415440 106519
rect 419460 97918 419488 107199
rect 415400 97912 415452 97918
rect 415400 97854 415452 97860
rect 419448 97912 419500 97918
rect 419448 97854 419500 97860
rect 440528 97730 440556 118798
rect 443644 118788 443696 118794
rect 443644 118730 443696 118736
rect 442264 118720 442316 118726
rect 442264 118662 442316 118668
rect 440358 97702 440556 97730
rect 421024 95062 421052 97036
rect 430684 95062 430712 97036
rect 442276 95062 442304 118662
rect 442998 106584 443054 106593
rect 442998 106519 443054 106528
rect 443012 97986 443040 106519
rect 443000 97980 443052 97986
rect 443000 97922 443052 97928
rect 443656 97850 443684 118730
rect 457272 116906 457300 118798
rect 467012 118720 467064 118726
rect 467012 118662 467064 118668
rect 468484 118720 468536 118726
rect 468484 118662 468536 118668
rect 467024 116906 467052 118662
rect 457272 116878 457654 116906
rect 467024 116878 467314 116906
rect 447244 116334 447994 116362
rect 445666 107264 445722 107273
rect 445666 107199 445722 107208
rect 445680 97986 445708 107199
rect 445668 97980 445720 97986
rect 445668 97922 445720 97928
rect 443644 97844 443696 97850
rect 443644 97786 443696 97792
rect 447244 95062 447272 116334
rect 447692 97844 447744 97850
rect 447692 97786 447744 97792
rect 467656 97844 467708 97850
rect 467656 97786 467708 97792
rect 447704 97730 447732 97786
rect 467668 97730 467696 97786
rect 447704 97702 447994 97730
rect 467406 97702 467696 97730
rect 421012 95056 421064 95062
rect 421012 94998 421064 95004
rect 430672 95056 430724 95062
rect 430672 94998 430724 95004
rect 442264 95056 442316 95062
rect 442264 94998 442316 95004
rect 447232 95056 447284 95062
rect 447232 94998 447284 95004
rect 457732 94994 457760 97036
rect 468496 94994 468524 118662
rect 468588 97850 468616 118798
rect 475384 118788 475436 118794
rect 475384 118730 475436 118736
rect 475396 116906 475424 118730
rect 475042 116878 475424 116906
rect 484412 116906 484440 118798
rect 494060 118720 494112 118726
rect 494060 118662 494112 118668
rect 494072 116906 494100 118662
rect 484412 116878 484702 116906
rect 494072 116878 494362 116906
rect 473266 106720 473322 106729
rect 473266 106655 473322 106664
rect 469218 106312 469274 106321
rect 469218 106247 469274 106256
rect 469232 97918 469260 106247
rect 473280 97918 473308 106655
rect 469220 97912 469272 97918
rect 469220 97854 469272 97860
rect 473268 97912 473320 97918
rect 473268 97854 473320 97860
rect 468576 97844 468628 97850
rect 468576 97786 468628 97792
rect 494532 97730 494560 118798
rect 494704 118788 494756 118794
rect 494704 118730 494756 118736
rect 494362 97702 494560 97730
rect 475028 95062 475056 97036
rect 484688 95062 484716 97036
rect 494716 96694 494744 118730
rect 496084 118720 496136 118726
rect 496084 118662 496136 118668
rect 494704 96688 494756 96694
rect 494704 96630 494756 96636
rect 496096 95062 496124 118662
rect 511368 116906 511396 118798
rect 522396 118788 522448 118794
rect 522396 118730 522448 118736
rect 520924 118720 520976 118726
rect 520924 118662 520976 118668
rect 522304 118720 522356 118726
rect 522304 118662 522356 118668
rect 520936 116906 520964 118662
rect 511368 116878 511658 116906
rect 520936 116878 521318 116906
rect 501064 116334 501998 116362
rect 500866 107264 500922 107273
rect 500866 107199 500922 107208
rect 496818 106584 496874 106593
rect 496818 106519 496874 106528
rect 496832 97986 496860 106519
rect 500880 97986 500908 107199
rect 496820 97980 496872 97986
rect 496820 97922 496872 97928
rect 500868 97980 500920 97986
rect 500868 97922 500920 97928
rect 501064 95062 501092 116334
rect 521752 100292 521804 100298
rect 521752 100234 521804 100240
rect 521764 97730 521792 100234
rect 521410 97702 521792 97730
rect 501616 97022 501998 97050
rect 501616 96694 501644 97022
rect 501604 96688 501656 96694
rect 501604 96630 501656 96636
rect 475016 95056 475068 95062
rect 475016 94998 475068 95004
rect 484676 95056 484728 95062
rect 484676 94998 484728 95004
rect 496084 95056 496136 95062
rect 496084 94998 496136 95004
rect 501052 95056 501104 95062
rect 501052 94998 501104 95004
rect 511736 94994 511764 97036
rect 522316 94994 522344 118662
rect 522408 100298 522436 118730
rect 528756 116906 528784 119342
rect 538404 118788 538456 118794
rect 538404 118730 538456 118736
rect 538416 116906 538444 118730
rect 548064 118720 548116 118726
rect 548064 118662 548116 118668
rect 548076 116906 548104 118662
rect 528756 116878 529046 116906
rect 538416 116878 538706 116906
rect 548076 116878 548366 116906
rect 526444 116612 526496 116618
rect 526444 116554 526496 116560
rect 526456 107409 526484 116554
rect 526442 107400 526498 107409
rect 526442 107335 526498 107344
rect 523038 106584 523094 106593
rect 523038 106519 523094 106528
rect 550638 106584 550694 106593
rect 550638 106519 550694 106528
rect 522396 100292 522448 100298
rect 522396 100234 522448 100240
rect 523052 97918 523080 106519
rect 550652 97986 550680 106519
rect 550640 97980 550692 97986
rect 550640 97922 550692 97928
rect 523040 97912 523092 97918
rect 523040 97854 523092 97860
rect 529032 95062 529060 97036
rect 529020 95056 529072 95062
rect 529020 94998 529072 95004
rect 150992 94988 151044 94994
rect 150992 94930 151044 94936
rect 160652 94988 160704 94994
rect 160652 94930 160704 94936
rect 171784 94988 171836 94994
rect 171784 94930 171836 94936
rect 214656 94988 214708 94994
rect 214656 94930 214708 94936
rect 225604 94988 225656 94994
rect 225604 94930 225656 94936
rect 268660 94988 268712 94994
rect 268660 94930 268712 94936
rect 279516 94988 279568 94994
rect 279516 94930 279568 94936
rect 285772 94988 285824 94994
rect 285772 94930 285824 94936
rect 295708 94988 295760 94994
rect 295708 94930 295760 94936
rect 307024 94988 307076 94994
rect 307024 94930 307076 94936
rect 311992 94988 312044 94994
rect 311992 94930 312044 94936
rect 322664 94988 322716 94994
rect 322664 94930 322716 94936
rect 333244 94988 333296 94994
rect 333244 94930 333296 94936
rect 339592 94988 339644 94994
rect 339592 94930 339644 94936
rect 349712 94988 349764 94994
rect 349712 94930 349764 94936
rect 359556 94988 359608 94994
rect 359556 94930 359608 94936
rect 365812 94988 365864 94994
rect 365812 94930 365864 94936
rect 376668 94988 376720 94994
rect 376668 94930 376720 94936
rect 387064 94988 387116 94994
rect 387064 94930 387116 94936
rect 393412 94988 393464 94994
rect 393412 94930 393464 94936
rect 403716 94988 403768 94994
rect 403716 94930 403768 94936
rect 414664 94988 414716 94994
rect 414664 94930 414716 94936
rect 457720 94988 457772 94994
rect 457720 94930 457772 94936
rect 468484 94988 468536 94994
rect 468484 94930 468536 94936
rect 511724 94988 511776 94994
rect 511724 94930 511776 94936
rect 522304 94988 522356 94994
rect 522304 94930 522356 94936
rect 538692 94926 538720 97036
rect 548352 95130 548380 97036
rect 548340 95124 548392 95130
rect 548340 95066 548392 95072
rect 538680 94920 538732 94926
rect 538680 94862 538732 94868
rect 529020 91792 529072 91798
rect 529020 91734 529072 91740
rect 149704 91384 149756 91390
rect 149704 91326 149756 91332
rect 148968 88392 149020 88398
rect 148968 88334 149020 88340
rect 148980 80345 149008 88334
rect 148966 80336 149022 80345
rect 148966 80271 149022 80280
rect 146944 69012 146996 69018
rect 146944 68954 146996 68960
rect 123668 68944 123720 68950
rect 123668 68886 123720 68892
rect 133788 68944 133840 68950
rect 133788 68886 133840 68892
rect 144184 68944 144236 68950
rect 144184 68886 144236 68892
rect 79968 68876 80020 68882
rect 79968 68818 80020 68824
rect 90364 68876 90416 68882
rect 90364 68818 90416 68824
rect 106556 68876 106608 68882
rect 106556 68818 106608 68824
rect 116584 68876 116636 68882
rect 116584 68818 116636 68824
rect 122932 68876 122984 68882
rect 122932 68818 122984 68824
rect 146944 65204 146996 65210
rect 146944 65146 146996 65152
rect 52460 65136 52512 65142
rect 52460 65078 52512 65084
rect 43352 65068 43404 65074
rect 43352 65010 43404 65016
rect 43364 62914 43392 65010
rect 43102 62886 43392 62914
rect 52472 62914 52500 65078
rect 62764 65068 62816 65074
rect 62764 65010 62816 65016
rect 90456 65068 90508 65074
rect 90456 65010 90508 65016
rect 106464 65068 106516 65074
rect 106464 65010 106516 65016
rect 116492 65068 116544 65074
rect 116492 65010 116544 65016
rect 133420 65068 133472 65074
rect 133420 65010 133472 65016
rect 62120 65000 62172 65006
rect 62120 64942 62172 64948
rect 62132 62914 62160 64942
rect 62488 64932 62540 64938
rect 62488 64874 62540 64880
rect 52472 62886 52670 62914
rect 62132 62886 62330 62914
rect 37924 62824 37976 62830
rect 37924 62766 37976 62772
rect 41328 62144 41380 62150
rect 41328 62086 41380 62092
rect 41340 53417 41368 62086
rect 41326 53408 41382 53417
rect 41326 53343 41382 53352
rect 37922 52864 37978 52873
rect 37922 52799 37978 52808
rect 36820 41268 36872 41274
rect 36820 41210 36872 41216
rect 36636 41132 36688 41138
rect 36636 41074 36688 41080
rect 36636 37460 36688 37466
rect 36636 37402 36688 37408
rect 36648 16590 36676 37402
rect 36728 37324 36780 37330
rect 36728 37266 36780 37272
rect 36636 16584 36688 16590
rect 36636 16526 36688 16532
rect 36544 13728 36596 13734
rect 36544 13670 36596 13676
rect 36740 13598 36768 37266
rect 37936 36650 37964 52799
rect 62500 43738 62528 64874
rect 62422 43710 62528 43738
rect 42996 41342 43024 43044
rect 52748 41342 52776 43044
rect 62776 41410 62804 65010
rect 64144 65000 64196 65006
rect 64144 64942 64196 64948
rect 89076 65000 89128 65006
rect 89076 64942 89128 64948
rect 90364 65000 90416 65006
rect 90364 64942 90416 64948
rect 62764 41404 62816 41410
rect 62764 41346 62816 41352
rect 64156 41342 64184 64942
rect 79324 64932 79376 64938
rect 79324 64874 79376 64880
rect 79336 62914 79364 64874
rect 89088 62914 89116 64942
rect 79336 62886 79718 62914
rect 89088 62886 89378 62914
rect 68928 62212 68980 62218
rect 68928 62154 68980 62160
rect 69124 62206 70058 62234
rect 68940 53825 68968 62154
rect 68926 53816 68982 53825
rect 68926 53751 68982 53760
rect 64878 52592 64934 52601
rect 64878 52527 64934 52536
rect 64892 44130 64920 52527
rect 64880 44124 64932 44130
rect 64880 44066 64932 44072
rect 69124 41342 69152 62206
rect 89720 50380 89772 50386
rect 89720 50322 89772 50328
rect 89732 43738 89760 50322
rect 89378 43710 89760 43738
rect 70044 41410 70072 43044
rect 70032 41404 70084 41410
rect 70032 41346 70084 41352
rect 42984 41336 43036 41342
rect 42984 41278 43036 41284
rect 52736 41336 52788 41342
rect 52736 41278 52788 41284
rect 64144 41336 64196 41342
rect 64144 41278 64196 41284
rect 69112 41336 69164 41342
rect 69112 41278 69164 41284
rect 79704 41274 79732 43044
rect 90376 41274 90404 64942
rect 90468 50386 90496 65010
rect 106476 62914 106504 65010
rect 116124 65000 116176 65006
rect 116124 64942 116176 64948
rect 116136 62914 116164 64942
rect 106476 62886 106674 62914
rect 116136 62886 116334 62914
rect 96724 62206 97014 62234
rect 91100 62144 91152 62150
rect 91100 62086 91152 62092
rect 91112 52737 91140 62086
rect 95146 53272 95202 53281
rect 95146 53207 95202 53216
rect 91098 52728 91154 52737
rect 91098 52663 91154 52672
rect 90456 50380 90508 50386
rect 90456 50322 90508 50328
rect 95160 44130 95188 53207
rect 95148 44124 95200 44130
rect 95148 44066 95200 44072
rect 96724 41410 96752 62206
rect 96712 41404 96764 41410
rect 96712 41346 96764 41352
rect 97000 41342 97028 43044
rect 96988 41336 97040 41342
rect 96988 41278 97040 41284
rect 106660 41274 106688 43044
rect 116320 42922 116348 43044
rect 116504 42922 116532 65010
rect 116584 65000 116636 65006
rect 116584 64942 116636 64948
rect 116320 42894 116532 42922
rect 116596 41274 116624 64942
rect 133432 62914 133460 65010
rect 142988 65000 143040 65006
rect 142988 64942 143040 64948
rect 144276 65000 144328 65006
rect 144276 64942 144328 64948
rect 143000 62914 143028 64942
rect 144184 64932 144236 64938
rect 144184 64874 144236 64880
rect 133432 62886 133722 62914
rect 143000 62886 143382 62914
rect 118700 62212 118752 62218
rect 118700 62154 118752 62160
rect 122748 62212 122800 62218
rect 122748 62154 122800 62160
rect 122944 62206 124062 62234
rect 118712 52737 118740 62154
rect 122760 53417 122788 62154
rect 122746 53408 122802 53417
rect 122746 53343 122802 53352
rect 118698 52728 118754 52737
rect 118698 52663 118754 52672
rect 79692 41268 79744 41274
rect 79692 41210 79744 41216
rect 90364 41268 90416 41274
rect 90364 41210 90416 41216
rect 106648 41268 106700 41274
rect 106648 41210 106700 41216
rect 116584 41268 116636 41274
rect 116584 41210 116636 41216
rect 122944 41206 122972 62206
rect 144196 45554 144224 64874
rect 143736 45526 144224 45554
rect 143736 43738 143764 45526
rect 143382 43710 143764 43738
rect 124048 41342 124076 43044
rect 124036 41336 124088 41342
rect 124036 41278 124088 41284
rect 133708 41274 133736 43044
rect 144288 41274 144316 64942
rect 146298 52864 146354 52873
rect 146298 52799 146354 52808
rect 146312 44130 146340 52799
rect 146300 44124 146352 44130
rect 146300 44066 146352 44072
rect 133696 41268 133748 41274
rect 133696 41210 133748 41216
rect 144276 41268 144328 41274
rect 144276 41210 144328 41216
rect 122932 41200 122984 41206
rect 122932 41142 122984 41148
rect 43076 37528 43128 37534
rect 43076 37470 43128 37476
rect 62764 37528 62816 37534
rect 62764 37470 62816 37476
rect 37924 36644 37976 36650
rect 37924 36586 37976 36592
rect 38016 36576 38068 36582
rect 38016 36518 38068 36524
rect 38028 26217 38056 36518
rect 43088 35972 43116 37470
rect 52644 37460 52696 37466
rect 52644 37402 52696 37408
rect 52656 35972 52684 37402
rect 62488 37392 62540 37398
rect 62488 37334 62540 37340
rect 62304 37324 62356 37330
rect 62304 37266 62356 37272
rect 62316 35972 62344 37266
rect 41328 34604 41380 34610
rect 41328 34546 41380 34552
rect 41340 26353 41368 34546
rect 41326 26344 41382 26353
rect 41326 26279 41382 26288
rect 38014 26208 38070 26217
rect 38014 26143 38070 26152
rect 62500 16674 62528 37334
rect 62422 16646 62528 16674
rect 42812 16102 43010 16130
rect 52762 16102 53144 16130
rect 42812 13666 42840 16102
rect 53116 13666 53144 16102
rect 62776 13802 62804 37470
rect 79692 37392 79744 37398
rect 79692 37334 79744 37340
rect 90364 37392 90416 37398
rect 90364 37334 90416 37340
rect 106648 37392 106700 37398
rect 106648 37334 106700 37340
rect 116492 37392 116544 37398
rect 116492 37334 116544 37340
rect 133696 37392 133748 37398
rect 133696 37334 133748 37340
rect 144184 37392 144236 37398
rect 144184 37334 144236 37340
rect 64144 37324 64196 37330
rect 64144 37266 64196 37272
rect 62764 13796 62816 13802
rect 62764 13738 62816 13744
rect 64156 13666 64184 37266
rect 79704 35972 79732 37334
rect 89352 37324 89404 37330
rect 89352 37266 89404 37272
rect 89364 35972 89392 37266
rect 69124 35278 70058 35306
rect 68928 34672 68980 34678
rect 68928 34614 68980 34620
rect 64880 34536 64932 34542
rect 64880 34478 64932 34484
rect 64892 25673 64920 34478
rect 68940 26897 68968 34614
rect 68926 26888 68982 26897
rect 68926 26823 68982 26832
rect 64878 25664 64934 25673
rect 64878 25599 64934 25608
rect 69124 13666 69152 35278
rect 90376 16574 90404 37334
rect 90456 37324 90508 37330
rect 90456 37266 90508 37272
rect 89824 16546 90404 16574
rect 89824 16538 89852 16546
rect 89378 16510 89852 16538
rect 69768 16102 70058 16130
rect 79718 16102 80008 16130
rect 69768 13802 69796 16102
rect 69756 13796 69808 13802
rect 69756 13738 69808 13744
rect 42800 13660 42852 13666
rect 42800 13602 42852 13608
rect 53104 13660 53156 13666
rect 53104 13602 53156 13608
rect 64144 13660 64196 13666
rect 64144 13602 64196 13608
rect 69112 13660 69164 13666
rect 69112 13602 69164 13608
rect 79980 13598 80008 16102
rect 90468 13598 90496 37266
rect 106660 35972 106688 37334
rect 116308 37324 116360 37330
rect 116308 37266 116360 37272
rect 116320 35972 116348 37266
rect 96724 35278 97014 35306
rect 91100 34604 91152 34610
rect 91100 34546 91152 34552
rect 91112 25673 91140 34546
rect 95148 34536 95200 34542
rect 95148 34478 95200 34484
rect 95160 26353 95188 34478
rect 95146 26344 95202 26353
rect 95146 26279 95202 26288
rect 91098 25664 91154 25673
rect 91098 25599 91154 25608
rect 96724 13598 96752 35278
rect 96816 16102 97014 16130
rect 106568 16102 106674 16130
rect 116228 16102 116334 16130
rect 96816 13666 96844 16102
rect 96804 13660 96856 13666
rect 96804 13602 96856 13608
rect 106568 13598 106596 16102
rect 116228 15858 116256 16102
rect 116504 15858 116532 37334
rect 116584 37324 116636 37330
rect 116584 37266 116636 37272
rect 116228 15830 116532 15858
rect 116596 13598 116624 37266
rect 133708 35972 133736 37334
rect 143356 37324 143408 37330
rect 143356 37266 143408 37272
rect 143368 35972 143396 37266
rect 122944 35278 124062 35306
rect 118700 34672 118752 34678
rect 118700 34614 118752 34620
rect 118712 25673 118740 34614
rect 122748 34604 122800 34610
rect 122748 34546 122800 34552
rect 122760 26353 122788 34546
rect 122746 26344 122802 26353
rect 122746 26279 122802 26288
rect 118698 25664 118754 25673
rect 118698 25599 118754 25608
rect 122944 13598 122972 35278
rect 144196 16574 144224 37334
rect 144276 37324 144328 37330
rect 144276 37266 144328 37272
rect 143736 16546 144224 16574
rect 143736 16538 143764 16546
rect 143382 16510 143764 16538
rect 123680 16102 124062 16130
rect 133722 16102 133828 16130
rect 123680 13666 123708 16102
rect 133800 13666 133828 16102
rect 144288 13666 144316 37266
rect 146300 34536 146352 34542
rect 146300 34478 146352 34484
rect 146312 25945 146340 34478
rect 146298 25936 146354 25945
rect 146298 25871 146354 25880
rect 146956 13734 146984 65146
rect 148968 62144 149020 62150
rect 148968 62086 149020 62092
rect 148980 53417 149008 62086
rect 148966 53408 149022 53417
rect 148966 53343 149022 53352
rect 149716 41342 149744 91326
rect 475016 91316 475068 91322
rect 475016 91258 475068 91264
rect 494704 91316 494756 91322
rect 494704 91258 494756 91264
rect 160652 91248 160704 91254
rect 160652 91190 160704 91196
rect 170496 91248 170548 91254
rect 170496 91190 170548 91196
rect 187700 91248 187752 91254
rect 187700 91190 187752 91196
rect 197452 91248 197504 91254
rect 197452 91190 197504 91196
rect 214656 91248 214708 91254
rect 214656 91190 214708 91196
rect 224500 91248 224552 91254
rect 224500 91190 224552 91196
rect 241704 91248 241756 91254
rect 241704 91190 241756 91196
rect 251456 91248 251508 91254
rect 251456 91190 251508 91196
rect 268660 91248 268712 91254
rect 268660 91190 268712 91196
rect 413468 91248 413520 91254
rect 413468 91190 413520 91196
rect 430672 91248 430724 91254
rect 430672 91190 430724 91196
rect 440516 91248 440568 91254
rect 440516 91190 440568 91196
rect 457628 91248 457680 91254
rect 457628 91190 457680 91196
rect 468484 91248 468536 91254
rect 468484 91190 468536 91196
rect 160664 89964 160692 91190
rect 170312 91180 170364 91186
rect 170312 91122 170364 91128
rect 170324 89964 170352 91122
rect 150544 89270 151018 89298
rect 150544 68882 150572 89270
rect 170232 70650 170338 70666
rect 170508 70650 170536 91190
rect 178040 91180 178092 91186
rect 178040 91122 178092 91128
rect 171784 91112 171836 91118
rect 171784 91054 171836 91060
rect 170220 70644 170338 70650
rect 170272 70638 170338 70644
rect 170496 70644 170548 70650
rect 170220 70586 170272 70592
rect 170496 70586 170548 70592
rect 150728 70094 151018 70122
rect 160572 70094 160678 70122
rect 150728 68950 150756 70094
rect 150716 68944 150768 68950
rect 150716 68886 150768 68892
rect 150532 68876 150584 68882
rect 150532 68818 150584 68824
rect 160572 68814 160600 70094
rect 171796 68814 171824 91054
rect 178052 89964 178080 91122
rect 187712 89964 187740 91190
rect 197360 91112 197412 91118
rect 197360 91054 197412 91060
rect 197372 89964 197400 91054
rect 172520 88460 172572 88466
rect 172520 88402 172572 88408
rect 176568 88460 176620 88466
rect 176568 88402 176620 88408
rect 172532 79665 172560 88402
rect 176580 80889 176608 88402
rect 176566 80880 176622 80889
rect 176566 80815 176622 80824
rect 172518 79656 172574 79665
rect 172518 79591 172574 79600
rect 197464 70666 197492 91190
rect 200764 91180 200816 91186
rect 200764 91122 200816 91128
rect 199384 91112 199436 91118
rect 199384 91054 199436 91060
rect 197386 70638 197492 70666
rect 178066 70094 178172 70122
rect 187726 70094 188016 70122
rect 178144 68882 178172 70094
rect 187988 68882 188016 70094
rect 199396 68882 199424 91054
rect 200120 88392 200172 88398
rect 200120 88334 200172 88340
rect 200132 79665 200160 88334
rect 200118 79656 200174 79665
rect 200118 79591 200174 79600
rect 200776 69018 200804 91122
rect 214668 89964 214696 91190
rect 224316 91112 224368 91118
rect 224316 91054 224368 91060
rect 224328 89964 224356 91054
rect 204364 89270 205022 89298
rect 202788 88392 202840 88398
rect 202788 88334 202840 88340
rect 202800 80345 202828 88334
rect 202786 80336 202842 80345
rect 202786 80271 202842 80280
rect 200764 69012 200816 69018
rect 200764 68954 200816 68960
rect 204364 68882 204392 89270
rect 224512 70666 224540 91190
rect 232044 91180 232096 91186
rect 232044 91122 232096 91128
rect 225604 91112 225656 91118
rect 225604 91054 225656 91060
rect 224342 70638 224540 70666
rect 204640 70094 205022 70122
rect 214682 70094 215064 70122
rect 204640 69018 204668 70094
rect 204628 69012 204680 69018
rect 204628 68954 204680 68960
rect 178132 68876 178184 68882
rect 178132 68818 178184 68824
rect 187976 68876 188028 68882
rect 187976 68818 188028 68824
rect 199384 68876 199436 68882
rect 199384 68818 199436 68824
rect 204352 68876 204404 68882
rect 204352 68818 204404 68824
rect 215036 68814 215064 70094
rect 225616 68814 225644 91054
rect 232056 89964 232084 91122
rect 241716 89964 241744 91190
rect 251364 91112 251416 91118
rect 251364 91054 251416 91060
rect 251376 89964 251404 91054
rect 230388 88528 230440 88534
rect 230388 88470 230440 88476
rect 226340 88460 226392 88466
rect 226340 88402 226392 88408
rect 226352 79665 226380 88402
rect 230400 80345 230428 88470
rect 230386 80336 230442 80345
rect 230386 80271 230442 80280
rect 226338 79656 226394 79665
rect 226338 79591 226394 79600
rect 251468 70666 251496 91190
rect 251824 91180 251876 91186
rect 251824 91122 251876 91128
rect 251390 70638 251496 70666
rect 231872 70094 232070 70122
rect 241730 70094 242112 70122
rect 231872 68882 231900 70094
rect 242084 68882 242112 70094
rect 251836 69018 251864 91122
rect 253204 91112 253256 91118
rect 253204 91054 253256 91060
rect 251824 69012 251876 69018
rect 251824 68954 251876 68960
rect 253216 68882 253244 91054
rect 268672 89964 268700 91190
rect 279424 91180 279476 91186
rect 279424 91122 279476 91128
rect 295708 91180 295760 91186
rect 295708 91122 295760 91128
rect 305460 91180 305512 91186
rect 305460 91122 305512 91128
rect 322664 91180 322716 91186
rect 322664 91122 322716 91128
rect 334624 91180 334676 91186
rect 334624 91122 334676 91128
rect 349712 91180 349764 91186
rect 349712 91122 349764 91128
rect 359464 91180 359516 91186
rect 359464 91122 359516 91128
rect 376668 91180 376720 91186
rect 376668 91122 376720 91128
rect 386512 91180 386564 91186
rect 386512 91122 386564 91128
rect 403624 91180 403676 91186
rect 403624 91122 403676 91128
rect 278320 91112 278372 91118
rect 278320 91054 278372 91060
rect 278332 89964 278360 91054
rect 258184 89270 259026 89298
rect 256608 88460 256660 88466
rect 256608 88402 256660 88408
rect 253940 88392 253992 88398
rect 253940 88334 253992 88340
rect 253952 80073 253980 88334
rect 256620 80345 256648 88402
rect 256606 80336 256662 80345
rect 256606 80271 256662 80280
rect 253938 80064 253994 80073
rect 253938 79999 253994 80008
rect 258184 68882 258212 89270
rect 279436 74534 279464 91122
rect 279516 91112 279568 91118
rect 279516 91054 279568 91060
rect 278792 74506 279464 74534
rect 278792 70666 278820 74506
rect 278346 70638 278820 70666
rect 258736 70094 259026 70122
rect 268686 70094 268976 70122
rect 258736 69018 258764 70094
rect 258724 69012 258776 69018
rect 258724 68954 258776 68960
rect 231860 68876 231912 68882
rect 231860 68818 231912 68824
rect 242072 68876 242124 68882
rect 242072 68818 242124 68824
rect 253204 68876 253256 68882
rect 253204 68818 253256 68824
rect 258172 68876 258224 68882
rect 258172 68818 258224 68824
rect 268948 68814 268976 70094
rect 279528 68814 279556 91054
rect 285784 90086 286088 90114
rect 280160 88528 280212 88534
rect 280160 88470 280212 88476
rect 280172 79665 280200 88470
rect 284208 88392 284260 88398
rect 284208 88334 284260 88340
rect 284220 80889 284248 88334
rect 284206 80880 284262 80889
rect 284206 80815 284262 80824
rect 280158 79656 280214 79665
rect 280158 79591 280214 79600
rect 285784 68882 285812 90086
rect 286060 89964 286088 90086
rect 295720 89964 295748 91122
rect 305368 91112 305420 91118
rect 305368 91054 305420 91060
rect 305380 89964 305408 91054
rect 305472 70666 305500 91122
rect 307024 91112 307076 91118
rect 307024 91054 307076 91060
rect 305394 70638 305500 70666
rect 286074 70094 286180 70122
rect 295734 70094 296024 70122
rect 285772 68876 285824 68882
rect 285772 68818 285824 68824
rect 286152 68814 286180 70094
rect 295996 68814 296024 70094
rect 307036 68814 307064 91054
rect 322676 89964 322704 91122
rect 332324 91112 332376 91118
rect 332324 91054 332376 91060
rect 333244 91112 333296 91118
rect 333244 91054 333296 91060
rect 332336 89964 332364 91054
rect 312004 89270 313030 89298
rect 307760 88460 307812 88466
rect 307760 88402 307812 88408
rect 311808 88460 311860 88466
rect 311808 88402 311860 88408
rect 307772 79665 307800 88402
rect 311820 80345 311848 88402
rect 311806 80336 311862 80345
rect 311806 80271 311862 80280
rect 307758 79656 307814 79665
rect 307758 79591 307814 79600
rect 312004 68814 312032 89270
rect 332508 71732 332560 71738
rect 332508 71674 332560 71680
rect 332520 70666 332548 71674
rect 332350 70638 332548 70666
rect 312648 70094 313030 70122
rect 322690 70094 322888 70122
rect 312648 68882 312676 70094
rect 312636 68876 312688 68882
rect 312636 68818 312688 68824
rect 322860 68814 322888 70094
rect 333256 68814 333284 91054
rect 334636 71738 334664 91122
rect 339604 90086 340092 90114
rect 335360 88392 335412 88398
rect 335360 88334 335412 88340
rect 338028 88392 338080 88398
rect 338028 88334 338080 88340
rect 335372 79665 335400 88334
rect 338040 80345 338068 88334
rect 338026 80336 338082 80345
rect 338026 80271 338082 80280
rect 335358 79656 335414 79665
rect 335358 79591 335414 79600
rect 334624 71732 334676 71738
rect 334624 71674 334676 71680
rect 339604 68814 339632 90086
rect 340064 89964 340092 90086
rect 349724 89964 349752 91122
rect 359372 91112 359424 91118
rect 359372 91054 359424 91060
rect 359384 89964 359412 91054
rect 359476 70666 359504 91122
rect 359556 91112 359608 91118
rect 359556 91054 359608 91060
rect 359398 70638 359504 70666
rect 340078 70094 340184 70122
rect 349738 70094 350120 70122
rect 340156 68882 340184 70094
rect 340144 68876 340196 68882
rect 340144 68818 340196 68824
rect 350092 68814 350120 70094
rect 359568 68814 359596 91054
rect 376680 89964 376708 91122
rect 386328 91112 386380 91118
rect 386328 91054 386380 91060
rect 386340 89964 386368 91054
rect 365824 89270 367034 89298
rect 361580 88460 361632 88466
rect 361580 88402 361632 88408
rect 365628 88460 365680 88466
rect 365628 88402 365680 88408
rect 361592 80073 361620 88402
rect 365640 80345 365668 88402
rect 365626 80336 365682 80345
rect 365626 80271 365682 80280
rect 361578 80064 361634 80073
rect 361578 79999 361634 80008
rect 365824 68882 365852 89270
rect 386524 70666 386552 91122
rect 387064 91112 387116 91118
rect 387064 91054 387116 91060
rect 386354 70638 386552 70666
rect 366744 70094 367034 70122
rect 376588 70094 376694 70122
rect 365812 68876 365864 68882
rect 365812 68818 365864 68824
rect 366744 68814 366772 70094
rect 376588 68814 376616 70094
rect 387076 68814 387104 91054
rect 403636 89964 403664 91122
rect 413284 91112 413336 91118
rect 413284 91054 413336 91060
rect 413296 89964 413324 91054
rect 393424 89270 393990 89298
rect 389180 88392 389232 88398
rect 389180 88334 389232 88340
rect 391848 88392 391900 88398
rect 391848 88334 391900 88340
rect 389192 79665 389220 88334
rect 391860 80345 391888 88334
rect 391846 80336 391902 80345
rect 391846 80271 391902 80280
rect 389178 79656 389234 79665
rect 389178 79591 389234 79600
rect 393424 68814 393452 89270
rect 413480 70666 413508 91190
rect 421012 91180 421064 91186
rect 421012 91122 421064 91128
rect 414664 91112 414716 91118
rect 414664 91054 414716 91060
rect 413402 70638 413508 70666
rect 393608 70094 393990 70122
rect 403742 70094 404032 70122
rect 393608 68882 393636 70094
rect 393596 68876 393648 68882
rect 393596 68818 393648 68824
rect 404004 68814 404032 70094
rect 414676 68814 414704 91054
rect 421024 89964 421052 91122
rect 430684 89964 430712 91190
rect 440332 91112 440384 91118
rect 440332 91054 440384 91060
rect 440344 89964 440372 91054
rect 415400 88460 415452 88466
rect 415400 88402 415452 88408
rect 419448 88460 419500 88466
rect 419448 88402 419500 88408
rect 415412 79665 415440 88402
rect 419460 80345 419488 88402
rect 419446 80336 419502 80345
rect 419446 80271 419502 80280
rect 415398 79656 415454 79665
rect 415398 79591 415454 79600
rect 440528 70666 440556 91190
rect 443644 91180 443696 91186
rect 443644 91122 443696 91128
rect 442264 91112 442316 91118
rect 442264 91054 442316 91060
rect 440358 70638 440556 70666
rect 420932 70094 421038 70122
rect 430698 70094 431080 70122
rect 420932 68882 420960 70094
rect 431052 68882 431080 70094
rect 442276 68882 442304 91054
rect 443000 88392 443052 88398
rect 443000 88334 443052 88340
rect 443012 79665 443040 88334
rect 442998 79656 443054 79665
rect 442998 79591 443054 79600
rect 443656 69018 443684 91122
rect 457640 89964 457668 91190
rect 467288 91112 467340 91118
rect 467288 91054 467340 91060
rect 467300 89964 467328 91054
rect 447244 89270 447994 89298
rect 445668 88392 445720 88398
rect 445668 88334 445720 88340
rect 445680 80345 445708 88334
rect 445666 80336 445722 80345
rect 445666 80271 445722 80280
rect 443644 69012 443696 69018
rect 443644 68954 443696 68960
rect 447244 68882 447272 89270
rect 468496 74534 468524 91190
rect 468576 91112 468628 91118
rect 468576 91054 468628 91060
rect 467852 74506 468524 74534
rect 467852 70666 467880 74506
rect 467406 70638 467880 70666
rect 447704 70094 447994 70122
rect 457746 70094 458128 70122
rect 447704 69018 447732 70094
rect 447692 69012 447744 69018
rect 447692 68954 447744 68960
rect 420920 68876 420972 68882
rect 420920 68818 420972 68824
rect 431040 68876 431092 68882
rect 431040 68818 431092 68824
rect 442264 68876 442316 68882
rect 442264 68818 442316 68824
rect 447232 68876 447284 68882
rect 447232 68818 447284 68824
rect 458100 68814 458128 70094
rect 468588 68814 468616 91054
rect 475028 89964 475056 91258
rect 484676 91248 484728 91254
rect 484676 91190 484728 91196
rect 484688 89964 484716 91190
rect 494520 91180 494572 91186
rect 494520 91122 494572 91128
rect 494336 91112 494388 91118
rect 494336 91054 494388 91060
rect 494348 89964 494376 91054
rect 469220 88460 469272 88466
rect 469220 88402 469272 88408
rect 473268 88460 473320 88466
rect 473268 88402 473320 88408
rect 469232 80073 469260 88402
rect 473280 80889 473308 88402
rect 473266 80880 473322 80889
rect 473266 80815 473322 80824
rect 469218 80064 469274 80073
rect 469218 79999 469274 80008
rect 494532 70666 494560 91122
rect 494362 70638 494560 70666
rect 474752 70094 475042 70122
rect 484702 70094 484992 70122
rect 474752 68882 474780 70094
rect 484964 68882 484992 70094
rect 494716 69018 494744 91258
rect 511632 91180 511684 91186
rect 511632 91122 511684 91128
rect 522304 91180 522356 91186
rect 522304 91122 522356 91128
rect 496084 91112 496136 91118
rect 496084 91054 496136 91060
rect 494704 69012 494756 69018
rect 494704 68954 494756 68960
rect 496096 68882 496124 91054
rect 511644 89964 511672 91122
rect 521292 91112 521344 91118
rect 521292 91054 521344 91060
rect 521304 89964 521332 91054
rect 501064 89270 501998 89298
rect 496820 88392 496872 88398
rect 496820 88334 496872 88340
rect 500868 88392 500920 88398
rect 500868 88334 500920 88340
rect 496832 79665 496860 88334
rect 500880 80345 500908 88334
rect 500866 80336 500922 80345
rect 500866 80271 500922 80280
rect 496818 79656 496874 79665
rect 496818 79591 496874 79600
rect 501064 68882 501092 89270
rect 522316 74534 522344 91122
rect 522396 91112 522448 91118
rect 522396 91054 522448 91060
rect 521856 74506 522344 74534
rect 521856 70666 521884 74506
rect 521410 70638 521884 70666
rect 501616 70094 501998 70122
rect 511750 70094 511948 70122
rect 501616 69018 501644 70094
rect 501604 69012 501656 69018
rect 501604 68954 501656 68960
rect 474740 68876 474792 68882
rect 474740 68818 474792 68824
rect 484952 68876 485004 68882
rect 484952 68818 485004 68824
rect 496084 68876 496136 68882
rect 496084 68818 496136 68824
rect 501052 68876 501104 68882
rect 501052 68818 501104 68824
rect 511920 68814 511948 70094
rect 522408 68814 522436 91054
rect 526444 90364 526496 90370
rect 526444 90306 526496 90312
rect 523040 88460 523092 88466
rect 523040 88402 523092 88408
rect 523052 79665 523080 88402
rect 526456 80345 526484 90306
rect 529032 89964 529060 91734
rect 538680 91180 538732 91186
rect 538680 91122 538732 91128
rect 538692 89964 538720 91122
rect 548340 91112 548392 91118
rect 548340 91054 548392 91060
rect 548352 89964 548380 91054
rect 550640 88392 550692 88398
rect 550640 88334 550692 88340
rect 526442 80336 526498 80345
rect 526442 80271 526498 80280
rect 550652 79665 550680 88334
rect 523038 79656 523094 79665
rect 523038 79591 523094 79600
rect 550638 79656 550694 79665
rect 550638 79591 550694 79600
rect 528756 70094 529046 70122
rect 538416 70094 538706 70122
rect 548076 70094 548366 70122
rect 528756 68882 528784 70094
rect 528744 68876 528796 68882
rect 528744 68818 528796 68824
rect 160560 68808 160612 68814
rect 160560 68750 160612 68756
rect 171784 68808 171836 68814
rect 171784 68750 171836 68756
rect 215024 68808 215076 68814
rect 215024 68750 215076 68756
rect 225604 68808 225656 68814
rect 225604 68750 225656 68756
rect 268936 68808 268988 68814
rect 268936 68750 268988 68756
rect 279516 68808 279568 68814
rect 279516 68750 279568 68756
rect 286140 68808 286192 68814
rect 286140 68750 286192 68756
rect 295984 68808 296036 68814
rect 295984 68750 296036 68756
rect 307024 68808 307076 68814
rect 307024 68750 307076 68756
rect 311992 68808 312044 68814
rect 311992 68750 312044 68756
rect 322848 68808 322900 68814
rect 322848 68750 322900 68756
rect 333244 68808 333296 68814
rect 333244 68750 333296 68756
rect 339592 68808 339644 68814
rect 339592 68750 339644 68756
rect 350080 68808 350132 68814
rect 350080 68750 350132 68756
rect 359556 68808 359608 68814
rect 359556 68750 359608 68756
rect 366732 68808 366784 68814
rect 366732 68750 366784 68756
rect 376576 68808 376628 68814
rect 376576 68750 376628 68756
rect 387064 68808 387116 68814
rect 387064 68750 387116 68756
rect 393412 68808 393464 68814
rect 393412 68750 393464 68756
rect 403992 68808 404044 68814
rect 403992 68750 404044 68756
rect 414664 68808 414716 68814
rect 414664 68750 414716 68756
rect 458088 68808 458140 68814
rect 458088 68750 458140 68756
rect 468576 68808 468628 68814
rect 468576 68750 468628 68756
rect 511908 68808 511960 68814
rect 511908 68750 511960 68756
rect 522396 68808 522448 68814
rect 522396 68750 522448 68756
rect 538416 68746 538444 70094
rect 548076 68950 548104 70094
rect 548064 68944 548116 68950
rect 548064 68886 548116 68892
rect 538404 68740 538456 68746
rect 538404 68682 538456 68688
rect 528652 65544 528704 65550
rect 528652 65486 528704 65492
rect 232320 65136 232372 65142
rect 232320 65078 232372 65084
rect 251824 65136 251876 65142
rect 251824 65078 251876 65084
rect 475384 65136 475436 65142
rect 475384 65078 475436 65084
rect 494704 65136 494756 65142
rect 494704 65078 494756 65084
rect 170496 65068 170548 65074
rect 170496 65010 170548 65016
rect 187792 65068 187844 65074
rect 187792 65010 187844 65016
rect 197544 65068 197596 65074
rect 197544 65010 197596 65016
rect 214380 65068 214432 65074
rect 214380 65010 214432 65016
rect 224500 65068 224552 65074
rect 224500 65010 224552 65016
rect 170036 65000 170088 65006
rect 170036 64942 170088 64948
rect 160284 64932 160336 64938
rect 160284 64874 160336 64880
rect 160296 62914 160324 64874
rect 170048 62914 170076 64942
rect 160296 62886 160678 62914
rect 170048 62886 170338 62914
rect 150544 62206 151018 62234
rect 149704 41336 149756 41342
rect 149704 41278 149756 41284
rect 150544 41274 150572 62206
rect 150532 41268 150584 41274
rect 150532 41210 150584 41216
rect 151004 41206 151032 43044
rect 160664 41206 160692 43044
rect 170324 42922 170352 43044
rect 170508 42922 170536 65010
rect 178408 65000 178460 65006
rect 178408 64942 178460 64948
rect 171784 64932 171836 64938
rect 171784 64874 171836 64880
rect 170324 42894 170536 42922
rect 171796 41206 171824 64874
rect 178420 62914 178448 64942
rect 187804 62914 187832 65010
rect 197452 64932 197504 64938
rect 197452 64874 197504 64880
rect 197464 62914 197492 64874
rect 178066 62886 178448 62914
rect 187726 62886 187832 62914
rect 197386 62886 197492 62914
rect 172520 62212 172572 62218
rect 172520 62154 172572 62160
rect 172532 52737 172560 62154
rect 172518 52728 172574 52737
rect 172518 52663 172574 52672
rect 176566 52728 176622 52737
rect 176566 52663 176622 52672
rect 176580 44130 176608 52663
rect 197556 45554 197584 65010
rect 200764 65000 200816 65006
rect 200764 64942 200816 64948
rect 199384 64932 199436 64938
rect 199384 64874 199436 64880
rect 197464 45526 197584 45554
rect 176568 44124 176620 44130
rect 176568 44066 176620 44072
rect 197464 43738 197492 45526
rect 197386 43710 197492 43738
rect 178052 41274 178080 43044
rect 187712 41274 187740 43044
rect 199396 41274 199424 64874
rect 200120 62144 200172 62150
rect 200120 62086 200172 62092
rect 200132 52737 200160 62086
rect 200118 52728 200174 52737
rect 200118 52663 200174 52672
rect 200776 41410 200804 64942
rect 214392 62914 214420 65010
rect 223948 64932 224000 64938
rect 223948 64874 224000 64880
rect 223960 62914 223988 64874
rect 214392 62886 214682 62914
rect 223960 62886 224342 62914
rect 204364 62206 205022 62234
rect 202788 62144 202840 62150
rect 202788 62086 202840 62092
rect 202800 53417 202828 62086
rect 202786 53408 202842 53417
rect 202786 53343 202842 53352
rect 200764 41404 200816 41410
rect 200764 41346 200816 41352
rect 204364 41274 204392 62206
rect 224512 43738 224540 65010
rect 225604 64932 225656 64938
rect 225604 64874 225656 64880
rect 224342 43710 224540 43738
rect 205008 41410 205036 43044
rect 204996 41404 205048 41410
rect 204996 41346 205048 41352
rect 178040 41268 178092 41274
rect 178040 41210 178092 41216
rect 187700 41268 187752 41274
rect 187700 41210 187752 41216
rect 199384 41268 199436 41274
rect 199384 41210 199436 41216
rect 204352 41268 204404 41274
rect 204352 41210 204404 41216
rect 214668 41206 214696 43044
rect 225616 41206 225644 64874
rect 232332 62914 232360 65078
rect 241612 65068 241664 65074
rect 241612 65010 241664 65016
rect 232070 62886 232360 62914
rect 241624 62914 241652 65010
rect 251456 65000 251508 65006
rect 251456 64942 251508 64948
rect 251272 64932 251324 64938
rect 251272 64874 251324 64880
rect 251284 62914 251312 64874
rect 241624 62886 241730 62914
rect 251284 62886 251390 62914
rect 230388 62212 230440 62218
rect 230388 62154 230440 62160
rect 230400 53417 230428 62154
rect 230386 53408 230442 53417
rect 230386 53343 230442 53352
rect 226338 52592 226394 52601
rect 226338 52527 226394 52536
rect 226352 44130 226380 52527
rect 226340 44124 226392 44130
rect 226340 44066 226392 44072
rect 251468 43738 251496 64942
rect 251390 43710 251496 43738
rect 232056 41274 232084 43044
rect 241716 41274 241744 43044
rect 251836 41410 251864 65078
rect 413468 65068 413520 65074
rect 413468 65010 413520 65016
rect 430580 65068 430632 65074
rect 430580 65010 430632 65016
rect 440516 65068 440568 65074
rect 440516 65010 440568 65016
rect 457260 65068 457312 65074
rect 457260 65010 457312 65016
rect 468576 65068 468628 65074
rect 468576 65010 468628 65016
rect 268292 65000 268344 65006
rect 268292 64942 268344 64948
rect 279424 65000 279476 65006
rect 279424 64942 279476 64948
rect 295800 65000 295852 65006
rect 295800 64942 295852 64948
rect 305552 65000 305604 65006
rect 305552 64942 305604 64948
rect 322388 65000 322440 65006
rect 322388 64942 322440 64948
rect 334624 65000 334676 65006
rect 334624 64942 334676 64948
rect 349804 65000 349856 65006
rect 349804 64942 349856 64948
rect 359648 65000 359700 65006
rect 359648 64942 359700 64948
rect 376300 65000 376352 65006
rect 376300 64942 376352 64948
rect 386512 65000 386564 65006
rect 386512 64942 386564 64948
rect 403348 65000 403400 65006
rect 403348 64942 403400 64948
rect 253204 64932 253256 64938
rect 253204 64874 253256 64880
rect 251824 41404 251876 41410
rect 251824 41346 251876 41352
rect 253216 41274 253244 64874
rect 268304 62914 268332 64942
rect 278044 64932 278096 64938
rect 278044 64874 278096 64880
rect 278056 62914 278084 64874
rect 268304 62886 268686 62914
rect 278056 62886 278346 62914
rect 258184 62206 259026 62234
rect 253940 62144 253992 62150
rect 253940 62086 253992 62092
rect 253952 53281 253980 62086
rect 253938 53272 253994 53281
rect 253938 53207 253994 53216
rect 256606 53272 256662 53281
rect 256606 53207 256662 53216
rect 256620 44130 256648 53207
rect 256608 44124 256660 44130
rect 256608 44066 256660 44072
rect 258184 41274 258212 62206
rect 279436 45554 279464 64942
rect 279516 64932 279568 64938
rect 279516 64874 279568 64880
rect 278792 45526 279464 45554
rect 278792 43738 278820 45526
rect 278346 43710 278820 43738
rect 259012 41410 259040 43044
rect 259000 41404 259052 41410
rect 259000 41346 259052 41352
rect 232044 41268 232096 41274
rect 232044 41210 232096 41216
rect 241704 41268 241756 41274
rect 241704 41210 241756 41216
rect 253204 41268 253256 41274
rect 253204 41210 253256 41216
rect 258172 41268 258224 41274
rect 258172 41210 258224 41216
rect 268672 41206 268700 43044
rect 279528 41206 279556 64874
rect 295812 62914 295840 64942
rect 305460 64932 305512 64938
rect 305460 64874 305512 64880
rect 305472 62914 305500 64874
rect 295734 62886 295840 62914
rect 305394 62886 305500 62914
rect 286074 62478 286180 62506
rect 286152 62422 286180 62478
rect 285772 62416 285824 62422
rect 285772 62358 285824 62364
rect 286140 62416 286192 62422
rect 286140 62358 286192 62364
rect 280160 62212 280212 62218
rect 280160 62154 280212 62160
rect 280172 52737 280200 62154
rect 284208 62144 284260 62150
rect 284208 62086 284260 62092
rect 284220 53825 284248 62086
rect 284206 53816 284262 53825
rect 284206 53751 284262 53760
rect 280158 52728 280214 52737
rect 280158 52663 280214 52672
rect 285784 41206 285812 62358
rect 305564 45554 305592 64942
rect 307024 64932 307076 64938
rect 307024 64874 307076 64880
rect 305472 45526 305592 45554
rect 305472 43738 305500 45526
rect 305394 43710 305500 43738
rect 286060 41274 286088 43044
rect 286048 41268 286100 41274
rect 286048 41210 286100 41216
rect 295720 41206 295748 43044
rect 307036 41206 307064 64874
rect 322400 62914 322428 64942
rect 331956 64932 332008 64938
rect 331956 64874 332008 64880
rect 333244 64932 333296 64938
rect 333244 64874 333296 64880
rect 331968 62914 331996 64874
rect 322400 62886 322690 62914
rect 331968 62886 332350 62914
rect 311808 62212 311860 62218
rect 311808 62154 311860 62160
rect 312004 62206 313030 62234
rect 311820 53417 311848 62154
rect 311806 53408 311862 53417
rect 311806 53343 311862 53352
rect 307758 52592 307814 52601
rect 307758 52527 307814 52536
rect 307772 44130 307800 52527
rect 307760 44124 307812 44130
rect 307760 44066 307812 44072
rect 312004 41206 312032 62206
rect 332508 44124 332560 44130
rect 332508 44066 332560 44072
rect 332520 43738 332548 44066
rect 332350 43710 332548 43738
rect 313016 41274 313044 43044
rect 313004 41268 313056 41274
rect 313004 41210 313056 41216
rect 322676 41206 322704 43044
rect 333256 41206 333284 64874
rect 334636 44130 334664 64942
rect 349816 62914 349844 64942
rect 359464 64932 359516 64938
rect 359464 64874 359516 64880
rect 359556 64932 359608 64938
rect 359556 64874 359608 64880
rect 359476 62914 359504 64874
rect 349738 62886 349844 62914
rect 359398 62886 359504 62914
rect 340078 62354 340184 62370
rect 339592 62348 339644 62354
rect 340078 62348 340196 62354
rect 340078 62342 340144 62348
rect 339592 62290 339644 62296
rect 340144 62290 340196 62296
rect 335360 62144 335412 62150
rect 335360 62086 335412 62092
rect 335372 52737 335400 62086
rect 338026 53272 338082 53281
rect 338026 53207 338082 53216
rect 335358 52728 335414 52737
rect 335358 52663 335414 52672
rect 338040 44130 338068 53207
rect 334624 44124 334676 44130
rect 334624 44066 334676 44072
rect 338028 44124 338080 44130
rect 338028 44066 338080 44072
rect 339604 41206 339632 62290
rect 359568 60178 359596 64874
rect 359556 60172 359608 60178
rect 359556 60114 359608 60120
rect 359660 60058 359688 64942
rect 376312 62914 376340 64942
rect 386052 64932 386104 64938
rect 386052 64874 386104 64880
rect 386064 62914 386092 64874
rect 376312 62886 376694 62914
rect 386064 62886 386354 62914
rect 361580 62212 361632 62218
rect 361580 62154 361632 62160
rect 365824 62206 367034 62234
rect 359476 60030 359688 60058
rect 359476 43738 359504 60030
rect 359556 59968 359608 59974
rect 359556 59910 359608 59916
rect 359398 43710 359504 43738
rect 340064 41274 340092 43044
rect 340052 41268 340104 41274
rect 340052 41210 340104 41216
rect 349724 41206 349752 43044
rect 359568 41206 359596 59910
rect 361592 53281 361620 62154
rect 365628 62144 365680 62150
rect 365628 62086 365680 62092
rect 365640 53417 365668 62086
rect 365626 53408 365682 53417
rect 365626 53343 365682 53352
rect 361578 53272 361634 53281
rect 361578 53207 361634 53216
rect 365824 41206 365852 62206
rect 386524 43738 386552 64942
rect 387064 64932 387116 64938
rect 387064 64874 387116 64880
rect 386354 43710 386552 43738
rect 367020 41274 367048 43044
rect 367008 41268 367060 41274
rect 367008 41210 367060 41216
rect 376680 41206 376708 43044
rect 387076 41206 387104 64874
rect 403360 62914 403388 64942
rect 412916 64932 412968 64938
rect 412916 64874 412968 64880
rect 412928 62914 412956 64874
rect 403360 62886 403650 62914
rect 412928 62886 413310 62914
rect 393424 62206 393990 62234
rect 391846 53272 391902 53281
rect 391846 53207 391902 53216
rect 389178 52592 389234 52601
rect 389178 52527 389234 52536
rect 389192 44130 389220 52527
rect 391860 44130 391888 53207
rect 389180 44124 389232 44130
rect 389180 44066 389232 44072
rect 391848 44124 391900 44130
rect 391848 44066 391900 44072
rect 393424 41206 393452 62206
rect 413480 43738 413508 65010
rect 421288 65000 421340 65006
rect 421288 64942 421340 64948
rect 414664 64932 414716 64938
rect 414664 64874 414716 64880
rect 413402 43710 413508 43738
rect 393976 41274 394004 43044
rect 393964 41268 394016 41274
rect 393964 41210 394016 41216
rect 403728 41206 403756 43044
rect 414676 41206 414704 64874
rect 421300 62914 421328 64942
rect 421038 62886 421328 62914
rect 430592 62914 430620 65010
rect 440240 64932 440292 64938
rect 440240 64874 440292 64880
rect 440252 62914 440280 64874
rect 430592 62886 430698 62914
rect 440252 62886 440358 62914
rect 415400 62144 415452 62150
rect 415400 62086 415452 62092
rect 419448 62144 419500 62150
rect 419448 62086 419500 62092
rect 415412 52737 415440 62086
rect 419460 53417 419488 62086
rect 419446 53408 419502 53417
rect 419446 53343 419502 53352
rect 415398 52728 415454 52737
rect 415398 52663 415454 52672
rect 440528 43738 440556 65010
rect 443644 65000 443696 65006
rect 443644 64942 443696 64948
rect 442264 64932 442316 64938
rect 442264 64874 442316 64880
rect 440358 43710 440556 43738
rect 421024 41274 421052 43044
rect 430684 41274 430712 43044
rect 442276 41274 442304 64874
rect 442998 52592 443054 52601
rect 442998 52527 443054 52536
rect 443012 44130 443040 52527
rect 443000 44124 443052 44130
rect 443000 44066 443052 44072
rect 443656 41410 443684 64942
rect 457272 62914 457300 65010
rect 467012 64932 467064 64938
rect 467012 64874 467064 64880
rect 468484 64932 468536 64938
rect 468484 64874 468536 64880
rect 467024 62914 467052 64874
rect 457272 62886 457654 62914
rect 467024 62886 467314 62914
rect 447244 62206 447994 62234
rect 445666 53272 445722 53281
rect 445666 53207 445722 53216
rect 445680 44130 445708 53207
rect 445668 44124 445720 44130
rect 445668 44066 445720 44072
rect 443644 41404 443696 41410
rect 443644 41346 443696 41352
rect 447244 41274 447272 62206
rect 467656 44056 467708 44062
rect 467656 43998 467708 44004
rect 467668 43738 467696 43998
rect 467406 43710 467696 43738
rect 447980 41410 448008 43044
rect 447968 41404 448020 41410
rect 447968 41346 448020 41352
rect 421012 41268 421064 41274
rect 421012 41210 421064 41216
rect 430672 41268 430724 41274
rect 430672 41210 430724 41216
rect 442264 41268 442316 41274
rect 442264 41210 442316 41216
rect 447232 41268 447284 41274
rect 447232 41210 447284 41216
rect 457732 41206 457760 43044
rect 468496 41206 468524 64874
rect 468588 44062 468616 65010
rect 475396 62914 475424 65078
rect 484400 65068 484452 65074
rect 484400 65010 484452 65016
rect 475042 62886 475424 62914
rect 484412 62914 484440 65010
rect 494520 65000 494572 65006
rect 494520 64942 494572 64948
rect 494060 64932 494112 64938
rect 494060 64874 494112 64880
rect 494072 62914 494100 64874
rect 484412 62886 484702 62914
rect 494072 62886 494362 62914
rect 473268 62212 473320 62218
rect 473268 62154 473320 62160
rect 469220 62144 469272 62150
rect 469220 62086 469272 62092
rect 469232 53281 469260 62086
rect 473280 53825 473308 62154
rect 473266 53816 473322 53825
rect 473266 53751 473322 53760
rect 469218 53272 469274 53281
rect 469218 53207 469274 53216
rect 468576 44056 468628 44062
rect 468576 43998 468628 44004
rect 494532 43738 494560 64942
rect 494362 43710 494560 43738
rect 475028 41274 475056 43044
rect 484688 41274 484716 43044
rect 494716 41410 494744 65078
rect 511356 65000 511408 65006
rect 511356 64942 511408 64948
rect 522304 65000 522356 65006
rect 522304 64942 522356 64948
rect 496084 64932 496136 64938
rect 496084 64874 496136 64880
rect 494704 41404 494756 41410
rect 494704 41346 494756 41352
rect 496096 41274 496124 64874
rect 511368 62914 511396 64942
rect 520924 64932 520976 64938
rect 520924 64874 520976 64880
rect 520936 62914 520964 64874
rect 511368 62886 511658 62914
rect 520936 62886 521318 62914
rect 501064 62206 501998 62234
rect 500868 62144 500920 62150
rect 500868 62086 500920 62092
rect 500880 53825 500908 62086
rect 500866 53816 500922 53825
rect 500866 53751 500922 53760
rect 496818 52592 496874 52601
rect 496818 52527 496874 52536
rect 496832 44130 496860 52527
rect 496820 44124 496872 44130
rect 496820 44066 496872 44072
rect 501064 41274 501092 62206
rect 522316 45554 522344 64942
rect 522396 64932 522448 64938
rect 522396 64874 522448 64880
rect 521856 45526 522344 45554
rect 521856 43738 521884 45526
rect 521410 43710 521884 43738
rect 501984 41410 502012 43044
rect 501972 41404 502024 41410
rect 501972 41346 502024 41352
rect 475016 41268 475068 41274
rect 475016 41210 475068 41216
rect 484676 41268 484728 41274
rect 484676 41210 484728 41216
rect 496084 41268 496136 41274
rect 496084 41210 496136 41216
rect 501052 41268 501104 41274
rect 501052 41210 501104 41216
rect 511736 41206 511764 43044
rect 522408 41206 522436 64874
rect 528664 62914 528692 65486
rect 538404 65000 538456 65006
rect 538404 64942 538456 64948
rect 538416 62914 538444 64942
rect 547972 64932 548024 64938
rect 547972 64874 548024 64880
rect 547984 62914 548012 64874
rect 528664 62886 529046 62914
rect 538416 62886 538706 62914
rect 547984 62886 548366 62914
rect 526444 62824 526496 62830
rect 526444 62766 526496 62772
rect 523040 62212 523092 62218
rect 523040 62154 523092 62160
rect 523052 52737 523080 62154
rect 526456 53417 526484 62766
rect 550640 62144 550692 62150
rect 550640 62086 550692 62092
rect 526442 53408 526498 53417
rect 526442 53343 526498 53352
rect 550652 53281 550680 62086
rect 550638 53272 550694 53281
rect 550638 53207 550694 53216
rect 523038 52728 523094 52737
rect 523038 52663 523094 52672
rect 529032 41274 529060 43044
rect 529020 41268 529072 41274
rect 529020 41210 529072 41216
rect 150992 41200 151044 41206
rect 150992 41142 151044 41148
rect 160652 41200 160704 41206
rect 160652 41142 160704 41148
rect 171784 41200 171836 41206
rect 171784 41142 171836 41148
rect 214656 41200 214708 41206
rect 214656 41142 214708 41148
rect 225604 41200 225656 41206
rect 225604 41142 225656 41148
rect 268660 41200 268712 41206
rect 268660 41142 268712 41148
rect 279516 41200 279568 41206
rect 279516 41142 279568 41148
rect 285772 41200 285824 41206
rect 285772 41142 285824 41148
rect 295708 41200 295760 41206
rect 295708 41142 295760 41148
rect 307024 41200 307076 41206
rect 307024 41142 307076 41148
rect 311992 41200 312044 41206
rect 311992 41142 312044 41148
rect 322664 41200 322716 41206
rect 322664 41142 322716 41148
rect 333244 41200 333296 41206
rect 333244 41142 333296 41148
rect 339592 41200 339644 41206
rect 339592 41142 339644 41148
rect 349712 41200 349764 41206
rect 349712 41142 349764 41148
rect 359556 41200 359608 41206
rect 359556 41142 359608 41148
rect 365812 41200 365864 41206
rect 365812 41142 365864 41148
rect 376668 41200 376720 41206
rect 376668 41142 376720 41148
rect 387064 41200 387116 41206
rect 387064 41142 387116 41148
rect 393412 41200 393464 41206
rect 393412 41142 393464 41148
rect 403716 41200 403768 41206
rect 403716 41142 403768 41148
rect 414664 41200 414716 41206
rect 414664 41142 414716 41148
rect 457720 41200 457772 41206
rect 457720 41142 457772 41148
rect 468484 41200 468536 41206
rect 468484 41142 468536 41148
rect 511724 41200 511776 41206
rect 511724 41142 511776 41148
rect 522396 41200 522448 41206
rect 522396 41142 522448 41148
rect 538692 41138 538720 43044
rect 548352 41342 548380 43044
rect 548340 41336 548392 41342
rect 548340 41278 548392 41284
rect 538680 41132 538732 41138
rect 538680 41074 538732 41080
rect 529020 38072 529072 38078
rect 529020 38014 529072 38020
rect 232044 37528 232096 37534
rect 232044 37470 232096 37476
rect 251824 37528 251876 37534
rect 251824 37470 251876 37476
rect 170496 37460 170548 37466
rect 170496 37402 170548 37408
rect 187700 37460 187752 37466
rect 187700 37402 187752 37408
rect 197452 37460 197504 37466
rect 197452 37402 197504 37408
rect 214656 37460 214708 37466
rect 214656 37402 214708 37408
rect 224500 37460 224552 37466
rect 224500 37402 224552 37408
rect 160652 37392 160704 37398
rect 160652 37334 160704 37340
rect 160664 35972 160692 37334
rect 170312 37324 170364 37330
rect 170312 37266 170364 37272
rect 170324 35972 170352 37266
rect 150544 35278 151018 35306
rect 148968 34536 149020 34542
rect 148968 34478 149020 34484
rect 148980 26353 149008 34478
rect 148966 26344 149022 26353
rect 148966 26279 149022 26288
rect 146944 13728 146996 13734
rect 146944 13670 146996 13676
rect 123668 13660 123720 13666
rect 123668 13602 123720 13608
rect 133788 13660 133840 13666
rect 133788 13602 133840 13608
rect 144276 13660 144328 13666
rect 144276 13602 144328 13608
rect 150544 13598 150572 35278
rect 150728 16102 151018 16130
rect 160572 16102 160678 16130
rect 170232 16102 170338 16130
rect 150728 13666 150756 16102
rect 150716 13660 150768 13666
rect 150716 13602 150768 13608
rect 25964 13592 26016 13598
rect 25964 13534 26016 13540
rect 36728 13592 36780 13598
rect 36728 13534 36780 13540
rect 79968 13592 80020 13598
rect 79968 13534 80020 13540
rect 90456 13592 90508 13598
rect 90456 13534 90508 13540
rect 96712 13592 96764 13598
rect 96712 13534 96764 13540
rect 106556 13592 106608 13598
rect 106556 13534 106608 13540
rect 116584 13592 116636 13598
rect 116584 13534 116636 13540
rect 122932 13592 122984 13598
rect 122932 13534 122984 13540
rect 150532 13592 150584 13598
rect 150532 13534 150584 13540
rect 160572 13530 160600 16102
rect 170232 15858 170260 16102
rect 170508 15858 170536 37402
rect 178040 37392 178092 37398
rect 178040 37334 178092 37340
rect 171784 37324 171836 37330
rect 171784 37266 171836 37272
rect 170232 15830 170536 15858
rect 171796 13530 171824 37266
rect 178052 35972 178080 37334
rect 187712 35972 187740 37402
rect 197360 37324 197412 37330
rect 197360 37266 197412 37272
rect 197372 35972 197400 37266
rect 172520 34604 172572 34610
rect 172520 34546 172572 34552
rect 176568 34604 176620 34610
rect 176568 34546 176620 34552
rect 172532 25673 172560 34546
rect 176580 26897 176608 34546
rect 176566 26888 176622 26897
rect 176566 26823 176622 26832
rect 172518 25664 172574 25673
rect 172518 25599 172574 25608
rect 197464 16674 197492 37402
rect 200764 37392 200816 37398
rect 200764 37334 200816 37340
rect 199384 37324 199436 37330
rect 199384 37266 199436 37272
rect 197386 16646 197492 16674
rect 178066 16102 178172 16130
rect 187726 16102 188016 16130
rect 178144 13598 178172 16102
rect 187988 13598 188016 16102
rect 199396 13598 199424 37266
rect 200120 34536 200172 34542
rect 200120 34478 200172 34484
rect 200132 25673 200160 34478
rect 200118 25664 200174 25673
rect 200118 25599 200174 25608
rect 200776 16590 200804 37334
rect 214668 35972 214696 37402
rect 224316 37324 224368 37330
rect 224316 37266 224368 37272
rect 224328 35972 224356 37266
rect 204364 35278 205022 35306
rect 202788 34536 202840 34542
rect 202788 34478 202840 34484
rect 202800 26353 202828 34478
rect 202786 26344 202842 26353
rect 202786 26279 202842 26288
rect 200764 16584 200816 16590
rect 200764 16526 200816 16532
rect 204364 13598 204392 35278
rect 224512 16674 224540 37402
rect 225604 37324 225656 37330
rect 225604 37266 225656 37272
rect 224342 16646 224540 16674
rect 204628 16584 204680 16590
rect 204680 16532 205022 16538
rect 204628 16526 205022 16532
rect 204640 16510 205022 16526
rect 214682 16102 215064 16130
rect 178132 13592 178184 13598
rect 178132 13534 178184 13540
rect 187976 13592 188028 13598
rect 187976 13534 188028 13540
rect 199384 13592 199436 13598
rect 199384 13534 199436 13540
rect 204352 13592 204404 13598
rect 204352 13534 204404 13540
rect 215036 13530 215064 16102
rect 225616 13530 225644 37266
rect 232056 35972 232084 37470
rect 241704 37460 241756 37466
rect 241704 37402 241756 37408
rect 241716 35972 241744 37402
rect 251456 37392 251508 37398
rect 251456 37334 251508 37340
rect 251364 37324 251416 37330
rect 251364 37266 251416 37272
rect 251376 35972 251404 37266
rect 226340 34604 226392 34610
rect 226340 34546 226392 34552
rect 230388 34604 230440 34610
rect 230388 34546 230440 34552
rect 226352 25673 226380 34546
rect 230400 26353 230428 34546
rect 230386 26344 230442 26353
rect 230386 26279 230442 26288
rect 226338 25664 226394 25673
rect 226338 25599 226394 25608
rect 251468 16674 251496 37334
rect 251390 16646 251496 16674
rect 231872 16102 232070 16130
rect 241730 16102 242112 16130
rect 231872 13598 231900 16102
rect 242084 13598 242112 16102
rect 251836 13802 251864 37470
rect 413468 37460 413520 37466
rect 413468 37402 413520 37408
rect 430672 37460 430724 37466
rect 430672 37402 430724 37408
rect 440516 37460 440568 37466
rect 440516 37402 440568 37408
rect 457628 37460 457680 37466
rect 457628 37402 457680 37408
rect 468484 37460 468536 37466
rect 468484 37402 468536 37408
rect 484676 37460 484728 37466
rect 484676 37402 484728 37408
rect 494520 37460 494572 37466
rect 494520 37402 494572 37408
rect 511632 37460 511684 37466
rect 511632 37402 511684 37408
rect 268660 37392 268712 37398
rect 268660 37334 268712 37340
rect 279424 37392 279476 37398
rect 279424 37334 279476 37340
rect 295708 37392 295760 37398
rect 295708 37334 295760 37340
rect 305460 37392 305512 37398
rect 305460 37334 305512 37340
rect 322664 37392 322716 37398
rect 322664 37334 322716 37340
rect 336004 37392 336056 37398
rect 336004 37334 336056 37340
rect 349712 37392 349764 37398
rect 349712 37334 349764 37340
rect 359464 37392 359516 37398
rect 359464 37334 359516 37340
rect 376668 37392 376720 37398
rect 376668 37334 376720 37340
rect 386512 37392 386564 37398
rect 386512 37334 386564 37340
rect 403624 37392 403676 37398
rect 403624 37334 403676 37340
rect 253204 37324 253256 37330
rect 253204 37266 253256 37272
rect 251824 13796 251876 13802
rect 251824 13738 251876 13744
rect 253216 13598 253244 37266
rect 268672 35972 268700 37334
rect 278320 37324 278372 37330
rect 278320 37266 278372 37272
rect 278332 35972 278360 37266
rect 258184 35278 259026 35306
rect 253940 34536 253992 34542
rect 253940 34478 253992 34484
rect 256608 34536 256660 34542
rect 256608 34478 256660 34484
rect 253952 25945 253980 34478
rect 256620 26353 256648 34478
rect 256606 26344 256662 26353
rect 256606 26279 256662 26288
rect 253938 25936 253994 25945
rect 253938 25871 253994 25880
rect 258184 13598 258212 35278
rect 279436 16574 279464 37334
rect 279516 37324 279568 37330
rect 279516 37266 279568 37272
rect 278792 16546 279464 16574
rect 278792 16538 278820 16546
rect 278346 16510 278820 16538
rect 258736 16102 259026 16130
rect 268686 16102 268976 16130
rect 258736 13802 258764 16102
rect 258724 13796 258776 13802
rect 258724 13738 258776 13744
rect 231860 13592 231912 13598
rect 231860 13534 231912 13540
rect 242072 13592 242124 13598
rect 242072 13534 242124 13540
rect 253204 13592 253256 13598
rect 253204 13534 253256 13540
rect 258172 13592 258224 13598
rect 258172 13534 258224 13540
rect 268948 13530 268976 16102
rect 279528 13530 279556 37266
rect 285968 36094 286088 36122
rect 285968 35894 285996 36094
rect 286060 35972 286088 36094
rect 295720 35972 295748 37334
rect 305368 37324 305420 37330
rect 305368 37266 305420 37272
rect 305380 35972 305408 37266
rect 285784 35866 285996 35894
rect 280160 34604 280212 34610
rect 280160 34546 280212 34552
rect 284208 34604 284260 34610
rect 284208 34546 284260 34552
rect 280172 25673 280200 34546
rect 284220 26897 284248 34546
rect 284206 26888 284262 26897
rect 284206 26823 284262 26832
rect 280158 25664 280214 25673
rect 280158 25599 280214 25608
rect 285784 13598 285812 35866
rect 305472 16674 305500 37334
rect 307024 37324 307076 37330
rect 307024 37266 307076 37272
rect 305394 16646 305500 16674
rect 286074 16102 286180 16130
rect 295734 16102 296024 16130
rect 285772 13592 285824 13598
rect 285772 13534 285824 13540
rect 286152 13530 286180 16102
rect 295996 13530 296024 16102
rect 307036 13530 307064 37266
rect 322676 35972 322704 37334
rect 332324 37324 332376 37330
rect 332324 37266 332376 37272
rect 333244 37324 333296 37330
rect 333244 37266 333296 37272
rect 332336 35972 332364 37266
rect 312004 35278 313030 35306
rect 311808 34672 311860 34678
rect 311808 34614 311860 34620
rect 307760 34536 307812 34542
rect 307760 34478 307812 34484
rect 307772 25673 307800 34478
rect 311820 26353 311848 34614
rect 311806 26344 311862 26353
rect 311806 26279 311862 26288
rect 307758 25664 307814 25673
rect 307758 25599 307814 25608
rect 312004 13530 312032 35278
rect 332508 16584 332560 16590
rect 332350 16532 332508 16538
rect 332350 16526 332560 16532
rect 332350 16510 332548 16526
rect 312648 16102 313030 16130
rect 322690 16102 322888 16130
rect 312648 13598 312676 16102
rect 312636 13592 312688 13598
rect 312636 13534 312688 13540
rect 322860 13530 322888 16102
rect 333256 13530 333284 37266
rect 335360 34604 335412 34610
rect 335360 34546 335412 34552
rect 335372 25673 335400 34546
rect 335358 25664 335414 25673
rect 335358 25599 335414 25608
rect 336016 16590 336044 37334
rect 339972 36094 340092 36122
rect 339972 35894 340000 36094
rect 340064 35972 340092 36094
rect 349724 35972 349752 37334
rect 359372 37324 359424 37330
rect 359372 37266 359424 37272
rect 359384 35972 359412 37266
rect 339604 35866 340000 35894
rect 338028 34536 338080 34542
rect 338028 34478 338080 34484
rect 338040 26353 338068 34478
rect 338026 26344 338082 26353
rect 338026 26279 338082 26288
rect 336004 16584 336056 16590
rect 336004 16526 336056 16532
rect 339604 13530 339632 35866
rect 359476 16674 359504 37334
rect 359556 37324 359608 37330
rect 359556 37266 359608 37272
rect 359398 16646 359504 16674
rect 340078 16102 340184 16130
rect 349738 16102 350120 16130
rect 340156 13598 340184 16102
rect 350092 13802 350120 16102
rect 359568 13802 359596 37266
rect 376680 35972 376708 37334
rect 386328 37324 386380 37330
rect 386328 37266 386380 37272
rect 386340 35972 386368 37266
rect 365824 35278 367034 35306
rect 361580 34672 361632 34678
rect 361580 34614 361632 34620
rect 361592 25945 361620 34614
rect 365628 34604 365680 34610
rect 365628 34546 365680 34552
rect 365640 26353 365668 34546
rect 365626 26344 365682 26353
rect 365626 26279 365682 26288
rect 361578 25936 361634 25945
rect 361578 25871 361634 25880
rect 350080 13796 350132 13802
rect 350080 13738 350132 13744
rect 359556 13796 359608 13802
rect 359556 13738 359608 13744
rect 365824 13598 365852 35278
rect 386524 16538 386552 37334
rect 387064 37324 387116 37330
rect 387064 37266 387116 37272
rect 386354 16510 386552 16538
rect 366744 16102 367034 16130
rect 376588 16102 376694 16130
rect 340144 13592 340196 13598
rect 340144 13534 340196 13540
rect 365812 13592 365864 13598
rect 365812 13534 365864 13540
rect 366744 13530 366772 16102
rect 376588 13530 376616 16102
rect 387076 13530 387104 37266
rect 403636 35972 403664 37334
rect 413284 37324 413336 37330
rect 413284 37266 413336 37272
rect 413296 35972 413324 37266
rect 393424 35278 393990 35306
rect 389180 34536 389232 34542
rect 389180 34478 389232 34484
rect 391848 34536 391900 34542
rect 391848 34478 391900 34484
rect 389192 25673 389220 34478
rect 391860 26353 391888 34478
rect 391846 26344 391902 26353
rect 391846 26279 391902 26288
rect 389178 25664 389234 25673
rect 389178 25599 389234 25608
rect 393424 13530 393452 35278
rect 413480 16674 413508 37402
rect 421012 37392 421064 37398
rect 421012 37334 421064 37340
rect 414664 37324 414716 37330
rect 414664 37266 414716 37272
rect 413402 16646 413508 16674
rect 393608 16102 393990 16130
rect 403742 16102 404032 16130
rect 393608 13598 393636 16102
rect 393596 13592 393648 13598
rect 393596 13534 393648 13540
rect 404004 13530 404032 16102
rect 414676 13530 414704 37266
rect 421024 35972 421052 37334
rect 430684 35972 430712 37402
rect 440332 37324 440384 37330
rect 440332 37266 440384 37272
rect 440344 35972 440372 37266
rect 415400 34604 415452 34610
rect 415400 34546 415452 34552
rect 419448 34604 419500 34610
rect 419448 34546 419500 34552
rect 415412 25673 415440 34546
rect 419460 26353 419488 34546
rect 419446 26344 419502 26353
rect 419446 26279 419502 26288
rect 415398 25664 415454 25673
rect 415398 25599 415454 25608
rect 440528 16674 440556 37402
rect 446404 37392 446456 37398
rect 446404 37334 446456 37340
rect 442264 37324 442316 37330
rect 442264 37266 442316 37272
rect 440358 16646 440556 16674
rect 420932 16102 421038 16130
rect 430698 16102 431080 16130
rect 420932 13598 420960 16102
rect 431052 13598 431080 16102
rect 442276 13598 442304 37266
rect 443000 34536 443052 34542
rect 443000 34478 443052 34484
rect 445668 34536 445720 34542
rect 445668 34478 445720 34484
rect 443012 25673 443040 34478
rect 445680 26353 445708 34478
rect 445666 26344 445722 26353
rect 445666 26279 445722 26288
rect 442998 25664 443054 25673
rect 442998 25599 443054 25608
rect 446416 16590 446444 37334
rect 457640 35972 457668 37402
rect 467288 37324 467340 37330
rect 467288 37266 467340 37272
rect 467300 35972 467328 37266
rect 447244 35278 447994 35306
rect 446404 16584 446456 16590
rect 446404 16526 446456 16532
rect 447244 13598 447272 35278
rect 447692 16584 447744 16590
rect 468496 16574 468524 37402
rect 475016 37392 475068 37398
rect 475016 37334 475068 37340
rect 468576 37324 468628 37330
rect 468576 37266 468628 37272
rect 467760 16546 468524 16574
rect 467760 16538 467788 16546
rect 447744 16532 447994 16538
rect 447692 16526 447994 16532
rect 447704 16510 447994 16526
rect 467406 16510 467788 16538
rect 457746 16102 458128 16130
rect 420920 13592 420972 13598
rect 420920 13534 420972 13540
rect 431040 13592 431092 13598
rect 431040 13534 431092 13540
rect 442264 13592 442316 13598
rect 442264 13534 442316 13540
rect 447232 13592 447284 13598
rect 447232 13534 447284 13540
rect 458100 13530 458128 16102
rect 468588 13530 468616 37266
rect 475028 35972 475056 37334
rect 484688 35972 484716 37402
rect 494336 37324 494388 37330
rect 494336 37266 494388 37272
rect 494348 35972 494376 37266
rect 469220 34604 469272 34610
rect 469220 34546 469272 34552
rect 473268 34604 473320 34610
rect 473268 34546 473320 34552
rect 469232 25945 469260 34546
rect 473280 26897 473308 34546
rect 473266 26888 473322 26897
rect 473266 26823 473322 26832
rect 469218 25936 469274 25945
rect 469218 25871 469274 25880
rect 494532 16674 494560 37402
rect 494704 37392 494756 37398
rect 494704 37334 494756 37340
rect 494362 16646 494560 16674
rect 474752 16102 475042 16130
rect 484702 16102 484992 16130
rect 474752 13598 474780 16102
rect 484964 13598 484992 16102
rect 494716 13802 494744 37334
rect 496084 37324 496136 37330
rect 496084 37266 496136 37272
rect 494704 13796 494756 13802
rect 494704 13738 494756 13744
rect 496096 13598 496124 37266
rect 511644 35972 511672 37402
rect 522396 37392 522448 37398
rect 522396 37334 522448 37340
rect 521292 37324 521344 37330
rect 521292 37266 521344 37272
rect 522304 37324 522356 37330
rect 522304 37266 522356 37272
rect 521304 35972 521332 37266
rect 501064 35278 501998 35306
rect 496820 34536 496872 34542
rect 496820 34478 496872 34484
rect 500868 34536 500920 34542
rect 500868 34478 500920 34484
rect 496832 25673 496860 34478
rect 500880 26353 500908 34478
rect 500866 26344 500922 26353
rect 500866 26279 500922 26288
rect 496818 25664 496874 25673
rect 496818 25599 496874 25608
rect 501064 13598 501092 35278
rect 521752 16584 521804 16590
rect 521410 16532 521752 16538
rect 521410 16526 521804 16532
rect 521410 16510 521792 16526
rect 501616 16102 501998 16130
rect 511750 16102 511948 16130
rect 501616 13802 501644 16102
rect 501604 13796 501656 13802
rect 501604 13738 501656 13744
rect 474740 13592 474792 13598
rect 474740 13534 474792 13540
rect 484952 13592 485004 13598
rect 484952 13534 485004 13540
rect 496084 13592 496136 13598
rect 496084 13534 496136 13540
rect 501052 13592 501104 13598
rect 501052 13534 501104 13540
rect 511920 13530 511948 16102
rect 522316 13530 522344 37266
rect 522408 16590 522436 37334
rect 526444 36644 526496 36650
rect 526444 36586 526496 36592
rect 523040 34604 523092 34610
rect 523040 34546 523092 34552
rect 523052 25673 523080 34546
rect 526456 26353 526484 36586
rect 529032 35972 529060 38014
rect 538680 37392 538732 37398
rect 538680 37334 538732 37340
rect 538692 35972 538720 37334
rect 548340 37324 548392 37330
rect 548340 37266 548392 37272
rect 548352 35972 548380 37266
rect 550640 34536 550692 34542
rect 550640 34478 550692 34484
rect 526442 26344 526498 26353
rect 526442 26279 526498 26288
rect 550652 25673 550680 34478
rect 523038 25664 523094 25673
rect 523038 25599 523094 25608
rect 550638 25664 550694 25673
rect 550638 25599 550694 25608
rect 522396 16584 522448 16590
rect 522396 16526 522448 16532
rect 528756 16102 529046 16130
rect 538416 16102 538706 16130
rect 548076 16102 548366 16130
rect 528756 13598 528784 16102
rect 538416 13734 538444 16102
rect 538404 13728 538456 13734
rect 538404 13670 538456 13676
rect 548076 13666 548104 16102
rect 548064 13660 548116 13666
rect 548064 13602 548116 13608
rect 528744 13592 528796 13598
rect 528744 13534 528796 13540
rect 160560 13524 160612 13530
rect 160560 13466 160612 13472
rect 171784 13524 171836 13530
rect 171784 13466 171836 13472
rect 215024 13524 215076 13530
rect 215024 13466 215076 13472
rect 225604 13524 225656 13530
rect 225604 13466 225656 13472
rect 268936 13524 268988 13530
rect 268936 13466 268988 13472
rect 279516 13524 279568 13530
rect 279516 13466 279568 13472
rect 286140 13524 286192 13530
rect 286140 13466 286192 13472
rect 295984 13524 296036 13530
rect 295984 13466 296036 13472
rect 307024 13524 307076 13530
rect 307024 13466 307076 13472
rect 311992 13524 312044 13530
rect 311992 13466 312044 13472
rect 322848 13524 322900 13530
rect 322848 13466 322900 13472
rect 333244 13524 333296 13530
rect 333244 13466 333296 13472
rect 339592 13524 339644 13530
rect 339592 13466 339644 13472
rect 366732 13524 366784 13530
rect 366732 13466 366784 13472
rect 376576 13524 376628 13530
rect 376576 13466 376628 13472
rect 387064 13524 387116 13530
rect 387064 13466 387116 13472
rect 393412 13524 393464 13530
rect 393412 13466 393464 13472
rect 403992 13524 404044 13530
rect 403992 13466 404044 13472
rect 414664 13524 414716 13530
rect 414664 13466 414716 13472
rect 458088 13524 458140 13530
rect 458088 13466 458140 13472
rect 468576 13524 468628 13530
rect 468576 13466 468628 13472
rect 511908 13524 511960 13530
rect 511908 13466 511960 13472
rect 522304 13524 522356 13530
rect 522304 13466 522356 13472
rect 580276 13462 580304 511255
rect 580354 458144 580410 458153
rect 580354 458079 580410 458088
rect 580368 37942 580396 458079
rect 580446 404968 580502 404977
rect 580446 404903 580502 404912
rect 580356 37936 580408 37942
rect 580356 37878 580408 37884
rect 580460 36582 580488 404903
rect 580538 351928 580594 351937
rect 580538 351863 580594 351872
rect 580552 38010 580580 351863
rect 580540 38004 580592 38010
rect 580540 37946 580592 37952
rect 580448 36576 580500 36582
rect 580448 36518 580500 36524
rect 16304 13456 16356 13462
rect 16304 13398 16356 13404
rect 580264 13456 580316 13462
rect 580264 13398 580316 13404
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 13726 674192 13782 674248
rect 13726 647264 13782 647320
rect 41326 674328 41382 674384
rect 37922 673784 37978 673840
rect 13726 620200 13782 620256
rect 13726 593136 13782 593192
rect 68926 674736 68982 674792
rect 64878 673512 64934 673568
rect 95146 674192 95202 674248
rect 91098 673648 91154 673704
rect 122746 674328 122802 674384
rect 118698 673648 118754 673704
rect 148966 674328 149022 674384
rect 146298 673512 146354 673568
rect 41326 647264 41382 647320
rect 37922 645904 37978 645960
rect 68926 647808 68982 647864
rect 64878 646584 64934 646640
rect 95146 647264 95202 647320
rect 91098 646584 91154 646640
rect 122746 647264 122802 647320
rect 118698 646584 118754 646640
rect 146298 647128 146354 647184
rect 41326 620200 41382 620256
rect 37922 618976 37978 619032
rect 13726 566208 13782 566264
rect 13726 539144 13782 539200
rect 68926 619656 68982 619712
rect 64878 619520 64934 619576
rect 95146 620200 95202 620256
rect 91098 619520 91154 619576
rect 122746 620200 122802 620256
rect 118698 619520 118754 619576
rect 146298 618976 146354 619032
rect 148966 647264 149022 647320
rect 176566 673784 176622 673840
rect 172518 673648 172574 673704
rect 200118 673648 200174 673704
rect 202786 674328 202842 674384
rect 230386 674328 230442 674384
rect 226338 673512 226394 673568
rect 253938 674192 253994 674248
rect 256606 674192 256662 674248
rect 284206 674736 284262 674792
rect 280158 673648 280214 673704
rect 311806 674328 311862 674384
rect 307758 673512 307814 673568
rect 338026 674192 338082 674248
rect 335358 673648 335414 673704
rect 365626 674328 365682 674384
rect 361578 674192 361634 674248
rect 391846 674192 391902 674248
rect 389178 673512 389234 673568
rect 419446 674328 419502 674384
rect 415398 673648 415454 673704
rect 442998 673512 443054 673568
rect 445666 674192 445722 674248
rect 473266 674736 473322 674792
rect 469218 674192 469274 674248
rect 500866 674328 500922 674384
rect 496818 673512 496874 673568
rect 527086 674192 527142 674248
rect 523038 673648 523094 673704
rect 176566 647808 176622 647864
rect 172518 646584 172574 646640
rect 200118 646584 200174 646640
rect 202786 647264 202842 647320
rect 230386 647264 230442 647320
rect 226338 646584 226394 646640
rect 256606 647264 256662 647320
rect 253938 647128 253994 647184
rect 284206 647808 284262 647864
rect 280158 646584 280214 646640
rect 311806 647264 311862 647320
rect 307758 646584 307814 646640
rect 335358 646584 335414 646640
rect 338026 647264 338082 647320
rect 365626 647264 365682 647320
rect 361578 647128 361634 647184
rect 391846 647264 391902 647320
rect 389178 646584 389234 646640
rect 419446 647264 419502 647320
rect 415398 646584 415454 646640
rect 445666 647264 445722 647320
rect 442998 646584 443054 646640
rect 473266 647808 473322 647864
rect 469218 647128 469274 647184
rect 500866 647264 500922 647320
rect 496818 646584 496874 646640
rect 526442 647264 526498 647320
rect 523038 646584 523094 646640
rect 41326 593136 41382 593192
rect 37922 592048 37978 592104
rect 68926 592592 68982 592648
rect 64878 592456 64934 592512
rect 95146 593136 95202 593192
rect 91098 592456 91154 592512
rect 122746 593136 122802 593192
rect 118698 592456 118754 592512
rect 146298 592048 146354 592104
rect 41326 566208 41382 566264
rect 37922 564984 37978 565040
rect 13726 512352 13782 512408
rect 13726 485152 13782 485208
rect 13726 458360 13782 458416
rect 68926 565800 68982 565856
rect 64878 565528 64934 565584
rect 95146 566208 95202 566264
rect 91098 565528 91154 565584
rect 122746 566208 122802 566264
rect 118698 565528 118754 565584
rect 146298 564984 146354 565040
rect 148966 620200 149022 620256
rect 176566 619656 176622 619712
rect 172518 619520 172574 619576
rect 200118 619520 200174 619576
rect 202786 620200 202842 620256
rect 230386 620200 230442 620256
rect 226338 619520 226394 619576
rect 256606 620200 256662 620256
rect 253938 618976 253994 619032
rect 284206 619656 284262 619712
rect 280158 619520 280214 619576
rect 311806 620200 311862 620256
rect 307758 619520 307814 619576
rect 335358 619520 335414 619576
rect 338026 620200 338082 620256
rect 365626 620200 365682 620256
rect 361578 618976 361634 619032
rect 391846 620200 391902 620256
rect 389178 619520 389234 619576
rect 419446 620200 419502 620256
rect 415398 619520 415454 619576
rect 442998 619520 443054 619576
rect 445666 620200 445722 620256
rect 473266 619656 473322 619712
rect 469218 618976 469274 619032
rect 500866 620200 500922 620256
rect 496818 619520 496874 619576
rect 526442 620336 526498 620392
rect 523038 619520 523094 619576
rect 148966 593136 149022 593192
rect 176566 592592 176622 592648
rect 172518 592456 172574 592512
rect 200118 592456 200174 592512
rect 202786 593136 202842 593192
rect 230386 593136 230442 593192
rect 226338 592456 226394 592512
rect 256606 593136 256662 593192
rect 253938 592048 253994 592104
rect 284206 592592 284262 592648
rect 280158 592456 280214 592512
rect 311806 593136 311862 593192
rect 307758 592456 307814 592512
rect 335358 592456 335414 592512
rect 338026 593136 338082 593192
rect 365626 593136 365682 593192
rect 361578 592048 361634 592104
rect 391846 592592 391902 592648
rect 389178 592456 389234 592512
rect 419446 593136 419502 593192
rect 415398 592456 415454 592512
rect 442998 592456 443054 592512
rect 445666 593136 445722 593192
rect 473266 592592 473322 592648
rect 469218 592048 469274 592104
rect 500866 593136 500922 593192
rect 496818 592456 496874 592512
rect 526442 593272 526498 593328
rect 523038 592456 523094 592512
rect 148966 566208 149022 566264
rect 41326 539144 41382 539200
rect 37922 538192 37978 538248
rect 68926 538600 68982 538656
rect 64878 538464 64934 538520
rect 95146 539144 95202 539200
rect 91098 538464 91154 538520
rect 122746 539144 122802 539200
rect 118698 538464 118754 538520
rect 146298 538328 146354 538384
rect 41326 512352 41382 512408
rect 37922 510992 37978 511048
rect 68926 512896 68982 512952
rect 64878 511672 64934 511728
rect 91098 511672 91154 511728
rect 96894 512896 96950 512952
rect 122746 512352 122802 512408
rect 118698 511672 118754 511728
rect 146298 511944 146354 512000
rect 148966 539144 149022 539200
rect 176566 565800 176622 565856
rect 172518 565528 172574 565584
rect 200118 565528 200174 565584
rect 202786 566208 202842 566264
rect 230386 566208 230442 566264
rect 226338 565528 226394 565584
rect 256606 566208 256662 566264
rect 253938 564984 253994 565040
rect 284206 565800 284262 565856
rect 280158 565528 280214 565584
rect 311806 566208 311862 566264
rect 307758 565528 307814 565584
rect 335358 565528 335414 565584
rect 338026 566208 338082 566264
rect 365626 566208 365682 566264
rect 361578 564984 361634 565040
rect 391846 566208 391902 566264
rect 389178 565528 389234 565584
rect 419446 566208 419502 566264
rect 415398 565528 415454 565584
rect 445666 566208 445722 566264
rect 442998 565528 443054 565584
rect 473266 565800 473322 565856
rect 469218 564984 469274 565040
rect 500866 566208 500922 566264
rect 496818 565528 496874 565584
rect 526442 566344 526498 566400
rect 523038 565528 523094 565584
rect 176566 538600 176622 538656
rect 172518 538464 172574 538520
rect 200118 538464 200174 538520
rect 202786 539144 202842 539200
rect 230386 539144 230442 539200
rect 226338 538464 226394 538520
rect 256606 539144 256662 539200
rect 253938 538328 253994 538384
rect 284206 538600 284262 538656
rect 280158 538464 280214 538520
rect 311806 539144 311862 539200
rect 307758 538464 307814 538520
rect 338026 539144 338082 539200
rect 335358 538464 335414 538520
rect 365626 539144 365682 539200
rect 361578 538328 361634 538384
rect 391846 539144 391902 539200
rect 389178 538464 389234 538520
rect 419446 539144 419502 539200
rect 415398 538464 415454 538520
rect 442998 538464 443054 538520
rect 445666 539144 445722 539200
rect 473266 538600 473322 538656
rect 469218 538328 469274 538384
rect 500866 539144 500922 539200
rect 496818 538464 496874 538520
rect 526442 539280 526498 539336
rect 523038 538464 523094 538520
rect 550638 673648 550694 673704
rect 550638 646584 550694 646640
rect 550638 619520 550694 619576
rect 550638 592048 550694 592104
rect 550638 565528 550694 565584
rect 550638 538464 550694 538520
rect 579802 524456 579858 524512
rect 148966 512352 149022 512408
rect 41326 485288 41382 485344
rect 37922 484880 37978 484936
rect 13726 431296 13782 431352
rect 13726 404232 13782 404288
rect 68926 485696 68982 485752
rect 64878 484472 64934 484528
rect 95146 485152 95202 485208
rect 91098 484608 91154 484664
rect 122746 485288 122802 485344
rect 118698 484608 118754 484664
rect 146298 484472 146354 484528
rect 41326 458360 41382 458416
rect 37922 457000 37978 457056
rect 68926 458904 68982 458960
rect 64878 457680 64934 457736
rect 95146 458360 95202 458416
rect 91098 457680 91154 457736
rect 122746 458360 122802 458416
rect 118698 457680 118754 457736
rect 146298 458088 146354 458144
rect 148966 485288 149022 485344
rect 176566 512896 176622 512952
rect 172518 511672 172574 511728
rect 200118 511672 200174 511728
rect 204902 512896 204958 512952
rect 230386 512352 230442 512408
rect 226338 511672 226394 511728
rect 256606 512352 256662 512408
rect 253938 511944 253994 512000
rect 284206 512896 284262 512952
rect 280158 511672 280214 511728
rect 311806 512352 311862 512408
rect 307758 511672 307814 511728
rect 335358 511672 335414 511728
rect 339866 512896 339922 512952
rect 365626 512352 365682 512408
rect 361578 511944 361634 512000
rect 391846 512896 391902 512952
rect 389178 511672 389234 511728
rect 419446 512352 419502 512408
rect 415398 511672 415454 511728
rect 442998 511808 443054 511864
rect 445666 512352 445722 512408
rect 473266 512896 473322 512952
rect 469218 511944 469274 512000
rect 500866 512896 500922 512952
rect 496818 511672 496874 511728
rect 526442 512352 526498 512408
rect 550638 511944 550694 512000
rect 523038 511672 523094 511728
rect 580262 511264 580318 511320
rect 172518 484608 172574 484664
rect 176566 484608 176622 484664
rect 200118 484608 200174 484664
rect 202786 485288 202842 485344
rect 230386 485288 230442 485344
rect 226338 484472 226394 484528
rect 253938 485152 253994 485208
rect 256606 485152 256662 485208
rect 284206 485696 284262 485752
rect 280158 484608 280214 484664
rect 311806 485288 311862 485344
rect 307758 484472 307814 484528
rect 338026 485152 338082 485208
rect 335358 484608 335414 484664
rect 365626 485288 365682 485344
rect 361578 485152 361634 485208
rect 391846 485152 391902 485208
rect 389178 484472 389234 484528
rect 419446 485288 419502 485344
rect 415398 484608 415454 484664
rect 442998 484472 443054 484528
rect 445666 485152 445722 485208
rect 473266 485696 473322 485752
rect 469218 485152 469274 485208
rect 500866 485288 500922 485344
rect 496818 484472 496874 484528
rect 526442 485288 526498 485344
rect 523038 484608 523094 484664
rect 550638 484608 550694 484664
rect 148966 458360 149022 458416
rect 41326 431296 41382 431352
rect 37922 430888 37978 430944
rect 13726 377168 13782 377224
rect 13726 350240 13782 350296
rect 68926 431568 68982 431624
rect 64878 430616 64934 430672
rect 95146 431296 95202 431352
rect 91098 430616 91154 430672
rect 122746 431296 122802 431352
rect 118698 430616 118754 430672
rect 146298 431160 146354 431216
rect 41326 404232 41382 404288
rect 37922 403008 37978 403064
rect 68926 403688 68982 403744
rect 64878 403552 64934 403608
rect 95146 404232 95202 404288
rect 91098 403552 91154 403608
rect 122746 404232 122802 404288
rect 118698 403552 118754 403608
rect 146298 403280 146354 403336
rect 148966 431296 149022 431352
rect 176566 458904 176622 458960
rect 172518 457680 172574 457736
rect 200118 457680 200174 457736
rect 202786 458360 202842 458416
rect 230386 458360 230442 458416
rect 226338 457680 226394 457736
rect 256606 458360 256662 458416
rect 253938 458088 253994 458144
rect 284206 458904 284262 458960
rect 280158 457680 280214 457736
rect 311806 458360 311862 458416
rect 307758 457680 307814 457736
rect 335358 457680 335414 457736
rect 338026 458360 338082 458416
rect 365626 458360 365682 458416
rect 361578 458088 361634 458144
rect 391846 458904 391902 458960
rect 389178 457680 389234 457736
rect 419446 458360 419502 458416
rect 415398 457680 415454 457736
rect 445666 458360 445722 458416
rect 442998 458088 443054 458144
rect 473266 458904 473322 458960
rect 469218 458088 469274 458144
rect 500866 458904 500922 458960
rect 496818 457680 496874 457736
rect 526442 458360 526498 458416
rect 550638 458088 550694 458144
rect 523038 457680 523094 457736
rect 176566 431568 176622 431624
rect 172518 430616 172574 430672
rect 200118 430616 200174 430672
rect 202786 431296 202842 431352
rect 230386 431296 230442 431352
rect 226338 430616 226394 430672
rect 256606 431296 256662 431352
rect 253938 431160 253994 431216
rect 284206 431568 284262 431624
rect 280158 430616 280214 430672
rect 311806 431296 311862 431352
rect 307758 430616 307814 430672
rect 338026 431296 338082 431352
rect 335358 430616 335414 430672
rect 365626 431296 365682 431352
rect 361578 431160 361634 431216
rect 391846 431296 391902 431352
rect 389178 430616 389234 430672
rect 419446 431296 419502 431352
rect 415398 430616 415454 430672
rect 442998 430616 443054 430672
rect 445666 431296 445722 431352
rect 473266 431568 473322 431624
rect 469218 431160 469274 431216
rect 500866 431296 500922 431352
rect 496818 430616 496874 430672
rect 526442 431296 526498 431352
rect 523038 430616 523094 430672
rect 550638 430616 550694 430672
rect 148966 404232 149022 404288
rect 41326 377168 41382 377224
rect 37922 375944 37978 376000
rect 13726 323176 13782 323232
rect 13726 296248 13782 296304
rect 13726 269320 13782 269376
rect 68926 376760 68982 376816
rect 64878 376488 64934 376544
rect 95146 377168 95202 377224
rect 91098 376488 91154 376544
rect 122746 377168 122802 377224
rect 118698 376488 118754 376544
rect 144826 375944 144882 376000
rect 41326 350240 41382 350296
rect 37922 349152 37978 349208
rect 68926 349696 68982 349752
rect 64878 349560 64934 349616
rect 95146 350240 95202 350296
rect 91098 349560 91154 349616
rect 122746 350240 122802 350296
rect 118698 349560 118754 349616
rect 146298 349152 146354 349208
rect 148966 377168 149022 377224
rect 176566 403688 176622 403744
rect 172518 403552 172574 403608
rect 200118 403552 200174 403608
rect 202786 404232 202842 404288
rect 230386 404232 230442 404288
rect 226338 403552 226394 403608
rect 256606 404232 256662 404288
rect 253938 403280 253994 403336
rect 284206 403688 284262 403744
rect 280158 403552 280214 403608
rect 311806 404232 311862 404288
rect 307758 403552 307814 403608
rect 335358 403552 335414 403608
rect 338026 404232 338082 404288
rect 365626 404232 365682 404288
rect 361578 403280 361634 403336
rect 391846 404232 391902 404288
rect 389178 403552 389234 403608
rect 419446 404232 419502 404288
rect 415398 403552 415454 403608
rect 442998 403552 443054 403608
rect 445666 404232 445722 404288
rect 473266 403688 473322 403744
rect 469218 403280 469274 403336
rect 500866 404232 500922 404288
rect 496818 403552 496874 403608
rect 526442 404232 526498 404288
rect 523038 403552 523094 403608
rect 550638 403552 550694 403608
rect 176566 376760 176622 376816
rect 172518 376488 172574 376544
rect 200118 376488 200174 376544
rect 202786 377168 202842 377224
rect 230386 377168 230442 377224
rect 226338 376488 226394 376544
rect 256606 377168 256662 377224
rect 253938 375944 253994 376000
rect 284206 376760 284262 376816
rect 280158 376488 280214 376544
rect 311806 377168 311862 377224
rect 307758 376488 307814 376544
rect 335358 376488 335414 376544
rect 338026 377168 338082 377224
rect 365626 377168 365682 377224
rect 361578 375944 361634 376000
rect 391846 377168 391902 377224
rect 389178 376488 389234 376544
rect 419446 377168 419502 377224
rect 415398 376488 415454 376544
rect 445666 377168 445722 377224
rect 442998 376488 443054 376544
rect 473266 376760 473322 376816
rect 469218 375944 469274 376000
rect 500866 377168 500922 377224
rect 496818 376488 496874 376544
rect 526442 377304 526498 377360
rect 523038 376488 523094 376544
rect 550638 376488 550694 376544
rect 148966 350240 149022 350296
rect 41326 323176 41382 323232
rect 37922 321952 37978 322008
rect 68926 322904 68982 322960
rect 64878 322496 64934 322552
rect 95146 323176 95202 323232
rect 91098 322496 91154 322552
rect 122746 323176 122802 323232
rect 118698 322496 118754 322552
rect 146298 321952 146354 322008
rect 41326 296248 41382 296304
rect 37922 295296 37978 295352
rect 13726 242120 13782 242176
rect 13726 215192 13782 215248
rect 68926 295704 68982 295760
rect 64878 295568 64934 295624
rect 95146 296248 95202 296304
rect 91098 295568 91154 295624
rect 122746 296248 122802 296304
rect 118698 295568 118754 295624
rect 146298 295296 146354 295352
rect 148966 323176 149022 323232
rect 176566 349696 176622 349752
rect 172518 349560 172574 349616
rect 200118 349560 200174 349616
rect 202786 350240 202842 350296
rect 230386 350240 230442 350296
rect 226338 349560 226394 349616
rect 256606 350240 256662 350296
rect 253938 349152 253994 349208
rect 284206 349696 284262 349752
rect 280158 349560 280214 349616
rect 311806 350240 311862 350296
rect 307758 349560 307814 349616
rect 338026 350240 338082 350296
rect 335358 349560 335414 349616
rect 365626 350240 365682 350296
rect 361578 349152 361634 349208
rect 391846 350240 391902 350296
rect 389178 349560 389234 349616
rect 419446 350240 419502 350296
rect 415398 349560 415454 349616
rect 442998 349560 443054 349616
rect 445666 350240 445722 350296
rect 473266 349696 473322 349752
rect 469218 349152 469274 349208
rect 500866 350240 500922 350296
rect 496818 349560 496874 349616
rect 526442 350240 526498 350296
rect 523038 349560 523094 349616
rect 550638 349560 550694 349616
rect 176566 322904 176622 322960
rect 172518 322496 172574 322552
rect 200118 322496 200174 322552
rect 202786 323176 202842 323232
rect 230386 323176 230442 323232
rect 226338 322496 226394 322552
rect 256606 323176 256662 323232
rect 253938 321952 253994 322008
rect 284206 322904 284262 322960
rect 280158 322496 280214 322552
rect 311806 323176 311862 323232
rect 307758 322496 307814 322552
rect 335358 322496 335414 322552
rect 338026 323176 338082 323232
rect 365626 323176 365682 323232
rect 361578 321952 361634 322008
rect 391846 323176 391902 323232
rect 389178 322496 389234 322552
rect 419446 323176 419502 323232
rect 415398 322496 415454 322552
rect 445666 323176 445722 323232
rect 442998 322496 443054 322552
rect 473266 322904 473322 322960
rect 469218 321952 469274 322008
rect 500866 323176 500922 323232
rect 496818 322496 496874 322552
rect 526442 323312 526498 323368
rect 523038 322496 523094 322552
rect 550638 322496 550694 322552
rect 148966 296248 149022 296304
rect 41326 269320 41382 269376
rect 37922 267960 37978 268016
rect 68926 269864 68982 269920
rect 64878 268640 64934 268696
rect 95146 269320 95202 269376
rect 91098 268640 91154 268696
rect 122746 269320 122802 269376
rect 118698 268640 118754 268696
rect 146298 269048 146354 269104
rect 41326 242256 41382 242312
rect 37922 241848 37978 241904
rect 13726 188128 13782 188184
rect 13726 161200 13782 161256
rect 68926 242800 68982 242856
rect 64878 241576 64934 241632
rect 95146 242120 95202 242176
rect 91098 241576 91154 241632
rect 122746 242256 122802 242312
rect 118698 241576 118754 241632
rect 146298 241848 146354 241904
rect 148966 269320 149022 269376
rect 176566 295704 176622 295760
rect 172518 295568 172574 295624
rect 200118 295568 200174 295624
rect 202786 296248 202842 296304
rect 230386 296248 230442 296304
rect 226338 295568 226394 295624
rect 256606 296248 256662 296304
rect 253938 295296 253994 295352
rect 284206 295704 284262 295760
rect 280158 295568 280214 295624
rect 311806 296248 311862 296304
rect 307758 295568 307814 295624
rect 338026 296248 338082 296304
rect 335358 295568 335414 295624
rect 365626 296248 365682 296304
rect 361578 295296 361634 295352
rect 391846 296248 391902 296304
rect 389178 295568 389234 295624
rect 419446 296248 419502 296304
rect 415398 295568 415454 295624
rect 442998 295568 443054 295624
rect 445666 296248 445722 296304
rect 473266 295704 473322 295760
rect 469218 295296 469274 295352
rect 500866 296248 500922 296304
rect 496818 295568 496874 295624
rect 526442 296248 526498 296304
rect 523038 295568 523094 295624
rect 550638 295568 550694 295624
rect 176566 269864 176622 269920
rect 172518 268640 172574 268696
rect 200118 268640 200174 268696
rect 202786 269320 202842 269376
rect 230386 269320 230442 269376
rect 226338 268640 226394 268696
rect 256606 269320 256662 269376
rect 253938 269048 253994 269104
rect 284206 269864 284262 269920
rect 280158 268640 280214 268696
rect 311806 269320 311862 269376
rect 307758 268640 307814 268696
rect 335358 268640 335414 268696
rect 338026 269320 338082 269376
rect 365626 269320 365682 269376
rect 361578 269048 361634 269104
rect 391846 269320 391902 269376
rect 389178 268640 389234 268696
rect 419446 269320 419502 269376
rect 415398 268640 415454 268696
rect 445666 269320 445722 269376
rect 442998 268640 443054 268696
rect 473266 269864 473322 269920
rect 469218 269048 469274 269104
rect 500866 269320 500922 269376
rect 496818 268640 496874 268696
rect 526442 269320 526498 269376
rect 523038 268640 523094 268696
rect 550638 268640 550694 268696
rect 41326 215192 41382 215248
rect 37922 213968 37978 214024
rect 68926 214648 68982 214704
rect 64878 214512 64934 214568
rect 95146 215192 95202 215248
rect 91098 214512 91154 214568
rect 122746 215192 122802 215248
rect 118698 214512 118754 214568
rect 146298 213968 146354 214024
rect 41326 188128 41382 188184
rect 37922 186904 37978 186960
rect 13726 134136 13782 134192
rect 13726 107208 13782 107264
rect 68926 187720 68982 187776
rect 64878 187448 64934 187504
rect 95146 188128 95202 188184
rect 91098 187448 91154 187504
rect 122746 188128 122802 188184
rect 118698 187448 118754 187504
rect 146298 186904 146354 186960
rect 148966 242256 149022 242312
rect 172518 241576 172574 241632
rect 176566 241576 176622 241632
rect 200118 241576 200174 241632
rect 202786 242256 202842 242312
rect 230386 242256 230442 242312
rect 226338 241576 226394 241632
rect 253938 242120 253994 242176
rect 256606 242120 256662 242176
rect 284206 242800 284262 242856
rect 280158 241576 280214 241632
rect 311806 242256 311862 242312
rect 307758 241576 307814 241632
rect 338026 242120 338082 242176
rect 335358 241576 335414 241632
rect 365626 242256 365682 242312
rect 361578 242120 361634 242176
rect 391846 241848 391902 241904
rect 389178 241576 389234 241632
rect 419446 242256 419502 242312
rect 415398 241576 415454 241632
rect 442998 241576 443054 241632
rect 445666 242120 445722 242176
rect 473266 242800 473322 242856
rect 469218 242120 469274 242176
rect 500866 242256 500922 242312
rect 496818 241576 496874 241632
rect 526442 242256 526498 242312
rect 523038 241576 523094 241632
rect 550638 241576 550694 241632
rect 148966 215192 149022 215248
rect 176566 214648 176622 214704
rect 172518 214512 172574 214568
rect 200118 214512 200174 214568
rect 202786 215192 202842 215248
rect 230386 215192 230442 215248
rect 226338 214512 226394 214568
rect 256606 215192 256662 215248
rect 253938 213968 253994 214024
rect 284206 214648 284262 214704
rect 280158 214512 280214 214568
rect 311806 215192 311862 215248
rect 307758 214512 307814 214568
rect 335358 214512 335414 214568
rect 338026 215192 338082 215248
rect 365626 215192 365682 215248
rect 361578 213968 361634 214024
rect 391846 215192 391902 215248
rect 389178 214512 389234 214568
rect 419446 215192 419502 215248
rect 415398 214512 415454 214568
rect 442998 214512 443054 214568
rect 445666 215192 445722 215248
rect 473266 214648 473322 214704
rect 469218 213968 469274 214024
rect 500866 215192 500922 215248
rect 496818 214512 496874 214568
rect 526442 215192 526498 215248
rect 523038 214512 523094 214568
rect 550638 214512 550694 214568
rect 148966 188128 149022 188184
rect 41326 161200 41382 161256
rect 37922 160112 37978 160168
rect 68926 160656 68982 160712
rect 64878 160520 64934 160576
rect 95146 161200 95202 161256
rect 91098 160520 91154 160576
rect 122746 161200 122802 161256
rect 118698 160520 118754 160576
rect 146298 160112 146354 160168
rect 41326 134136 41382 134192
rect 37922 132912 37978 132968
rect 13726 80280 13782 80336
rect 13726 53216 13782 53272
rect 13726 26288 13782 26344
rect 68926 133864 68982 133920
rect 64878 133456 64934 133512
rect 95146 134136 95202 134192
rect 91098 133456 91154 133512
rect 122746 134136 122802 134192
rect 118698 133456 118754 133512
rect 146298 132912 146354 132968
rect 148966 161200 149022 161256
rect 176566 187720 176622 187776
rect 172518 187448 172574 187504
rect 200118 187448 200174 187504
rect 202786 188128 202842 188184
rect 230386 188128 230442 188184
rect 226338 187448 226394 187504
rect 256606 188128 256662 188184
rect 253938 186904 253994 186960
rect 284206 187720 284262 187776
rect 280158 187448 280214 187504
rect 311806 188128 311862 188184
rect 307758 187448 307814 187504
rect 335358 187448 335414 187504
rect 338026 188128 338082 188184
rect 365626 188128 365682 188184
rect 361578 186904 361634 186960
rect 391846 187720 391902 187776
rect 389178 187448 389234 187504
rect 419446 188128 419502 188184
rect 415398 187448 415454 187504
rect 445666 188128 445722 188184
rect 442998 186904 443054 186960
rect 473266 187720 473322 187776
rect 469218 186904 469274 186960
rect 500866 187720 500922 187776
rect 496818 187448 496874 187504
rect 526442 188264 526498 188320
rect 523038 187448 523094 187504
rect 550638 186904 550694 186960
rect 176566 160656 176622 160712
rect 172518 160520 172574 160576
rect 200118 160520 200174 160576
rect 202786 161200 202842 161256
rect 230386 161200 230442 161256
rect 226338 160520 226394 160576
rect 256606 161200 256662 161256
rect 253938 160112 253994 160168
rect 284206 160656 284262 160712
rect 280158 160520 280214 160576
rect 311806 161200 311862 161256
rect 307758 160520 307814 160576
rect 338026 161200 338082 161256
rect 335358 160520 335414 160576
rect 365626 161200 365682 161256
rect 361578 160112 361634 160168
rect 391846 161200 391902 161256
rect 389178 160520 389234 160576
rect 419446 161200 419502 161256
rect 415398 160520 415454 160576
rect 442998 160520 443054 160576
rect 445666 161200 445722 161256
rect 473266 160656 473322 160712
rect 469218 160112 469274 160168
rect 500866 161200 500922 161256
rect 496818 160520 496874 160576
rect 526442 161336 526498 161392
rect 523038 160520 523094 160576
rect 550638 160520 550694 160576
rect 148966 134136 149022 134192
rect 41326 107208 41382 107264
rect 37922 106528 37978 106584
rect 68926 106664 68982 106720
rect 64878 106528 64934 106584
rect 95146 107208 95202 107264
rect 91098 106528 91154 106584
rect 122746 107208 122802 107264
rect 118698 106528 118754 106584
rect 146298 106256 146354 106312
rect 41326 80280 41382 80336
rect 37922 78920 37978 78976
rect 68926 80824 68982 80880
rect 64878 79600 64934 79656
rect 95146 80280 95202 80336
rect 91098 79600 91154 79656
rect 122746 80280 122802 80336
rect 118698 79600 118754 79656
rect 146298 80008 146354 80064
rect 148966 107208 149022 107264
rect 176566 133864 176622 133920
rect 172518 133456 172574 133512
rect 200118 133456 200174 133512
rect 202786 134136 202842 134192
rect 230386 134136 230442 134192
rect 226338 133456 226394 133512
rect 256606 134136 256662 134192
rect 253938 132912 253994 132968
rect 284206 133864 284262 133920
rect 280158 133456 280214 133512
rect 311806 134136 311862 134192
rect 307758 133456 307814 133512
rect 335358 133456 335414 133512
rect 338026 134136 338082 134192
rect 365626 134136 365682 134192
rect 361578 132912 361634 132968
rect 391846 133864 391902 133920
rect 389178 133456 389234 133512
rect 419446 134136 419502 134192
rect 415398 133456 415454 133512
rect 442998 133456 443054 133512
rect 445666 134136 445722 134192
rect 473266 133864 473322 133920
rect 469218 132912 469274 132968
rect 500866 134136 500922 134192
rect 496818 133456 496874 133512
rect 526442 134272 526498 134328
rect 523038 133456 523094 133512
rect 550638 132912 550694 132968
rect 176566 106664 176622 106720
rect 172518 106528 172574 106584
rect 200118 106528 200174 106584
rect 202786 107208 202842 107264
rect 230386 107208 230442 107264
rect 226338 106528 226394 106584
rect 256606 107208 256662 107264
rect 253938 106256 253994 106312
rect 284206 106664 284262 106720
rect 280158 106528 280214 106584
rect 311806 107208 311862 107264
rect 307758 106528 307814 106584
rect 338026 107208 338082 107264
rect 335358 106528 335414 106584
rect 365626 107208 365682 107264
rect 361578 106256 361634 106312
rect 391846 107208 391902 107264
rect 389178 106528 389234 106584
rect 419446 107208 419502 107264
rect 415398 106528 415454 106584
rect 442998 106528 443054 106584
rect 445666 107208 445722 107264
rect 473266 106664 473322 106720
rect 469218 106256 469274 106312
rect 500866 107208 500922 107264
rect 496818 106528 496874 106584
rect 526442 107344 526498 107400
rect 523038 106528 523094 106584
rect 550638 106528 550694 106584
rect 148966 80280 149022 80336
rect 41326 53352 41382 53408
rect 37922 52808 37978 52864
rect 68926 53760 68982 53816
rect 64878 52536 64934 52592
rect 95146 53216 95202 53272
rect 91098 52672 91154 52728
rect 122746 53352 122802 53408
rect 118698 52672 118754 52728
rect 146298 52808 146354 52864
rect 41326 26288 41382 26344
rect 38014 26152 38070 26208
rect 68926 26832 68982 26888
rect 64878 25608 64934 25664
rect 95146 26288 95202 26344
rect 91098 25608 91154 25664
rect 122746 26288 122802 26344
rect 118698 25608 118754 25664
rect 146298 25880 146354 25936
rect 148966 53352 149022 53408
rect 176566 80824 176622 80880
rect 172518 79600 172574 79656
rect 200118 79600 200174 79656
rect 202786 80280 202842 80336
rect 230386 80280 230442 80336
rect 226338 79600 226394 79656
rect 256606 80280 256662 80336
rect 253938 80008 253994 80064
rect 284206 80824 284262 80880
rect 280158 79600 280214 79656
rect 311806 80280 311862 80336
rect 307758 79600 307814 79656
rect 338026 80280 338082 80336
rect 335358 79600 335414 79656
rect 365626 80280 365682 80336
rect 361578 80008 361634 80064
rect 391846 80280 391902 80336
rect 389178 79600 389234 79656
rect 419446 80280 419502 80336
rect 415398 79600 415454 79656
rect 442998 79600 443054 79656
rect 445666 80280 445722 80336
rect 473266 80824 473322 80880
rect 469218 80008 469274 80064
rect 500866 80280 500922 80336
rect 496818 79600 496874 79656
rect 526442 80280 526498 80336
rect 523038 79600 523094 79656
rect 550638 79600 550694 79656
rect 172518 52672 172574 52728
rect 176566 52672 176622 52728
rect 200118 52672 200174 52728
rect 202786 53352 202842 53408
rect 230386 53352 230442 53408
rect 226338 52536 226394 52592
rect 253938 53216 253994 53272
rect 256606 53216 256662 53272
rect 284206 53760 284262 53816
rect 280158 52672 280214 52728
rect 311806 53352 311862 53408
rect 307758 52536 307814 52592
rect 338026 53216 338082 53272
rect 335358 52672 335414 52728
rect 365626 53352 365682 53408
rect 361578 53216 361634 53272
rect 391846 53216 391902 53272
rect 389178 52536 389234 52592
rect 419446 53352 419502 53408
rect 415398 52672 415454 52728
rect 442998 52536 443054 52592
rect 445666 53216 445722 53272
rect 473266 53760 473322 53816
rect 469218 53216 469274 53272
rect 500866 53760 500922 53816
rect 496818 52536 496874 52592
rect 526442 53352 526498 53408
rect 550638 53216 550694 53272
rect 523038 52672 523094 52728
rect 148966 26288 149022 26344
rect 176566 26832 176622 26888
rect 172518 25608 172574 25664
rect 200118 25608 200174 25664
rect 202786 26288 202842 26344
rect 230386 26288 230442 26344
rect 226338 25608 226394 25664
rect 256606 26288 256662 26344
rect 253938 25880 253994 25936
rect 284206 26832 284262 26888
rect 280158 25608 280214 25664
rect 311806 26288 311862 26344
rect 307758 25608 307814 25664
rect 335358 25608 335414 25664
rect 338026 26288 338082 26344
rect 365626 26288 365682 26344
rect 361578 25880 361634 25936
rect 391846 26288 391902 26344
rect 389178 25608 389234 25664
rect 419446 26288 419502 26344
rect 415398 25608 415454 25664
rect 445666 26288 445722 26344
rect 442998 25608 443054 25664
rect 473266 26832 473322 26888
rect 469218 25880 469274 25936
rect 500866 26288 500922 26344
rect 496818 25608 496874 25664
rect 526442 26288 526498 26344
rect 523038 25608 523094 25664
rect 550638 25608 550694 25664
rect 580354 458088 580410 458144
rect 580446 404912 580502 404968
rect 580538 351872 580594 351928
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect 68921 674794 68987 674797
rect 284201 674794 284267 674797
rect 473261 674794 473327 674797
rect 68921 674792 70226 674794
rect 68921 674736 68926 674792
rect 68982 674736 70226 674792
rect 68921 674734 70226 674736
rect 68921 674731 68987 674734
rect 41321 674386 41387 674389
rect 41321 674384 43148 674386
rect 41321 674328 41326 674384
rect 41382 674328 43148 674384
rect 70166 674356 70226 674734
rect 284201 674792 286242 674794
rect 284201 674736 284206 674792
rect 284262 674736 286242 674792
rect 284201 674734 286242 674736
rect 284201 674731 284267 674734
rect 122741 674386 122807 674389
rect 148961 674386 149027 674389
rect 202781 674386 202847 674389
rect 230381 674386 230447 674389
rect 122741 674384 124108 674386
rect 41321 674326 43148 674328
rect 122741 674328 122746 674384
rect 122802 674328 124108 674384
rect 122741 674326 124108 674328
rect 148961 674384 151156 674386
rect 148961 674328 148966 674384
rect 149022 674328 151156 674384
rect 148961 674326 151156 674328
rect 202781 674384 205068 674386
rect 202781 674328 202786 674384
rect 202842 674328 205068 674384
rect 202781 674326 205068 674328
rect 230381 674384 232116 674386
rect 230381 674328 230386 674384
rect 230442 674328 232116 674384
rect 286182 674356 286242 674734
rect 473261 674792 475210 674794
rect 473261 674736 473266 674792
rect 473322 674736 475210 674792
rect 473261 674734 475210 674736
rect 473261 674731 473327 674734
rect 311801 674386 311867 674389
rect 365621 674386 365687 674389
rect 419441 674386 419507 674389
rect 311801 674384 313076 674386
rect 230381 674326 232116 674328
rect 311801 674328 311806 674384
rect 311862 674328 313076 674384
rect 311801 674326 313076 674328
rect 365621 674384 367172 674386
rect 365621 674328 365626 674384
rect 365682 674328 367172 674384
rect 365621 674326 367172 674328
rect 419441 674384 421084 674386
rect 419441 674328 419446 674384
rect 419502 674328 421084 674384
rect 475150 674356 475210 674734
rect 500861 674386 500927 674389
rect 500861 674384 502044 674386
rect 419441 674326 421084 674328
rect 500861 674328 500866 674384
rect 500922 674328 502044 674384
rect 500861 674326 502044 674328
rect 41321 674323 41387 674326
rect 122741 674323 122807 674326
rect 148961 674323 149027 674326
rect 202781 674323 202847 674326
rect 230381 674323 230447 674326
rect 311801 674323 311867 674326
rect 365621 674323 365687 674326
rect 419441 674323 419507 674326
rect 500861 674323 500927 674326
rect 13721 674250 13787 674253
rect 95141 674250 95207 674253
rect 253933 674250 253999 674253
rect 13721 674248 16100 674250
rect 13721 674192 13726 674248
rect 13782 674192 16100 674248
rect 13721 674190 16100 674192
rect 95141 674248 97060 674250
rect 95141 674192 95146 674248
rect 95202 674192 97060 674248
rect 251774 674248 253999 674250
rect 95141 674190 97060 674192
rect 13721 674187 13787 674190
rect 95141 674187 95207 674190
rect 37917 673842 37983 673845
rect 35758 673840 37983 673842
rect 35758 673784 37922 673840
rect 37978 673784 37983 673840
rect 35758 673782 37983 673784
rect 35758 673676 35818 673782
rect 37917 673779 37983 673782
rect 176561 673842 176627 673845
rect 178174 673842 178234 674220
rect 176561 673840 178234 673842
rect 176561 673784 176566 673840
rect 176622 673784 178234 673840
rect 176561 673782 178234 673784
rect 251774 674192 253938 674248
rect 253994 674192 253999 674248
rect 251774 674190 253999 674192
rect 176561 673779 176627 673782
rect 91093 673706 91159 673709
rect 118693 673706 118759 673709
rect 172513 673706 172579 673709
rect 200113 673706 200179 673709
rect 89884 673704 91159 673706
rect 89884 673648 91098 673704
rect 91154 673648 91159 673704
rect 89884 673646 91159 673648
rect 116932 673704 118759 673706
rect 116932 673648 118698 673704
rect 118754 673648 118759 673704
rect 116932 673646 118759 673648
rect 170844 673704 172579 673706
rect 170844 673648 172518 673704
rect 172574 673648 172579 673704
rect 170844 673646 172579 673648
rect 197892 673704 200179 673706
rect 197892 673648 200118 673704
rect 200174 673648 200179 673704
rect 251774 673676 251834 674190
rect 253933 674187 253999 674190
rect 256601 674250 256667 674253
rect 338021 674250 338087 674253
rect 361573 674250 361639 674253
rect 256601 674248 259164 674250
rect 256601 674192 256606 674248
rect 256662 674192 259164 674248
rect 256601 674190 259164 674192
rect 338021 674248 340124 674250
rect 338021 674192 338026 674248
rect 338082 674192 340124 674248
rect 338021 674190 340124 674192
rect 359782 674248 361639 674250
rect 359782 674192 361578 674248
rect 361634 674192 361639 674248
rect 359782 674190 361639 674192
rect 256601 674187 256667 674190
rect 338021 674187 338087 674190
rect 280153 673706 280219 673709
rect 335353 673706 335419 673709
rect 278852 673704 280219 673706
rect 197892 673646 200179 673648
rect 278852 673648 280158 673704
rect 280214 673648 280219 673704
rect 278852 673646 280219 673648
rect 332948 673704 335419 673706
rect 332948 673648 335358 673704
rect 335414 673648 335419 673704
rect 359782 673676 359842 674190
rect 361573 674187 361639 674190
rect 391841 674250 391907 674253
rect 445661 674250 445727 674253
rect 469213 674250 469279 674253
rect 391841 674248 394036 674250
rect 391841 674192 391846 674248
rect 391902 674192 394036 674248
rect 391841 674190 394036 674192
rect 445661 674248 448132 674250
rect 445661 674192 445666 674248
rect 445722 674192 448132 674248
rect 445661 674190 448132 674192
rect 467790 674248 469279 674250
rect 467790 674192 469218 674248
rect 469274 674192 469279 674248
rect 467790 674190 469279 674192
rect 391841 674187 391907 674190
rect 445661 674187 445727 674190
rect 415393 673706 415459 673709
rect 413908 673704 415459 673706
rect 332948 673646 335419 673648
rect 413908 673648 415398 673704
rect 415454 673648 415459 673704
rect 467790 673676 467850 674190
rect 469213 674187 469279 674190
rect 527081 674250 527147 674253
rect 527081 674248 529092 674250
rect 527081 674192 527086 674248
rect 527142 674192 529092 674248
rect 527081 674190 529092 674192
rect 527081 674187 527147 674190
rect 523033 673706 523099 673709
rect 550633 673706 550699 673709
rect 521916 673704 523099 673706
rect 413908 673646 415459 673648
rect 521916 673648 523038 673704
rect 523094 673648 523099 673704
rect 521916 673646 523099 673648
rect 548964 673704 550699 673706
rect 548964 673648 550638 673704
rect 550694 673648 550699 673704
rect 548964 673646 550699 673648
rect 91093 673643 91159 673646
rect 118693 673643 118759 673646
rect 172513 673643 172579 673646
rect 200113 673643 200179 673646
rect 280153 673643 280219 673646
rect 335353 673643 335419 673646
rect 415393 673643 415459 673646
rect 523033 673643 523099 673646
rect 550633 673643 550699 673646
rect 64873 673570 64939 673573
rect 146293 673570 146359 673573
rect 226333 673570 226399 673573
rect 307753 673570 307819 673573
rect 389173 673570 389239 673573
rect 442993 673570 443059 673573
rect 496813 673570 496879 673573
rect 62836 673568 64939 673570
rect 62836 673512 64878 673568
rect 64934 673512 64939 673568
rect 143950 673568 146359 673570
rect 62836 673510 64939 673512
rect 64873 673507 64939 673510
rect 143766 673470 143826 673540
rect 143950 673512 146298 673568
rect 146354 673512 146359 673568
rect 143950 673510 146359 673512
rect 224940 673568 226399 673570
rect 224940 673512 226338 673568
rect 226394 673512 226399 673568
rect 224940 673510 226399 673512
rect 305900 673568 307819 673570
rect 305900 673512 307758 673568
rect 307814 673512 307819 673568
rect 305900 673510 307819 673512
rect 386860 673568 389239 673570
rect 386860 673512 389178 673568
rect 389234 673512 389239 673568
rect 386860 673510 389239 673512
rect 440956 673568 443059 673570
rect 440956 673512 442998 673568
rect 443054 673512 443059 673568
rect 440956 673510 443059 673512
rect 494868 673568 496879 673570
rect 494868 673512 496818 673568
rect 496874 673512 496879 673568
rect 494868 673510 496879 673512
rect 143950 673470 144010 673510
rect 146293 673507 146359 673510
rect 226333 673507 226399 673510
rect 307753 673507 307819 673510
rect 389173 673507 389239 673510
rect 442993 673507 443059 673510
rect 496813 673507 496879 673510
rect 143766 673410 144010 673470
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect 68921 647866 68987 647869
rect 176561 647866 176627 647869
rect 284201 647866 284267 647869
rect 473261 647866 473327 647869
rect 68921 647864 70226 647866
rect 68921 647808 68926 647864
rect 68982 647808 70226 647864
rect 68921 647806 70226 647808
rect 68921 647803 68987 647806
rect 13721 647322 13787 647325
rect 41321 647322 41387 647325
rect 13721 647320 16100 647322
rect 13721 647264 13726 647320
rect 13782 647264 16100 647320
rect 13721 647262 16100 647264
rect 41321 647320 43148 647322
rect 41321 647264 41326 647320
rect 41382 647264 43148 647320
rect 70166 647292 70226 647806
rect 176561 647864 178234 647866
rect 176561 647808 176566 647864
rect 176622 647808 178234 647864
rect 176561 647806 178234 647808
rect 176561 647803 176627 647806
rect 95141 647322 95207 647325
rect 122741 647322 122807 647325
rect 148961 647322 149027 647325
rect 95141 647320 97060 647322
rect 41321 647262 43148 647264
rect 95141 647264 95146 647320
rect 95202 647264 97060 647320
rect 95141 647262 97060 647264
rect 122741 647320 124108 647322
rect 122741 647264 122746 647320
rect 122802 647264 124108 647320
rect 122741 647262 124108 647264
rect 148961 647320 151156 647322
rect 148961 647264 148966 647320
rect 149022 647264 151156 647320
rect 178174 647292 178234 647806
rect 284201 647864 286242 647866
rect 284201 647808 284206 647864
rect 284262 647808 286242 647864
rect 284201 647806 286242 647808
rect 284201 647803 284267 647806
rect 202781 647322 202847 647325
rect 230381 647322 230447 647325
rect 256601 647322 256667 647325
rect 202781 647320 205068 647322
rect 148961 647262 151156 647264
rect 202781 647264 202786 647320
rect 202842 647264 205068 647320
rect 202781 647262 205068 647264
rect 230381 647320 232116 647322
rect 230381 647264 230386 647320
rect 230442 647264 232116 647320
rect 230381 647262 232116 647264
rect 256601 647320 259164 647322
rect 256601 647264 256606 647320
rect 256662 647264 259164 647320
rect 286182 647292 286242 647806
rect 473261 647864 475210 647866
rect 473261 647808 473266 647864
rect 473322 647808 475210 647864
rect 473261 647806 475210 647808
rect 473261 647803 473327 647806
rect 311801 647322 311867 647325
rect 338021 647322 338087 647325
rect 365621 647322 365687 647325
rect 391841 647322 391907 647325
rect 419441 647322 419507 647325
rect 445661 647322 445727 647325
rect 311801 647320 313076 647322
rect 256601 647262 259164 647264
rect 311801 647264 311806 647320
rect 311862 647264 313076 647320
rect 311801 647262 313076 647264
rect 338021 647320 340124 647322
rect 338021 647264 338026 647320
rect 338082 647264 340124 647320
rect 338021 647262 340124 647264
rect 365621 647320 367172 647322
rect 365621 647264 365626 647320
rect 365682 647264 367172 647320
rect 365621 647262 367172 647264
rect 391841 647320 394036 647322
rect 391841 647264 391846 647320
rect 391902 647264 394036 647320
rect 391841 647262 394036 647264
rect 419441 647320 421084 647322
rect 419441 647264 419446 647320
rect 419502 647264 421084 647320
rect 419441 647262 421084 647264
rect 445661 647320 448132 647322
rect 445661 647264 445666 647320
rect 445722 647264 448132 647320
rect 475150 647292 475210 647806
rect 500861 647322 500927 647325
rect 526437 647322 526503 647325
rect 500861 647320 502044 647322
rect 445661 647262 448132 647264
rect 500861 647264 500866 647320
rect 500922 647264 502044 647320
rect 500861 647262 502044 647264
rect 526437 647320 529092 647322
rect 526437 647264 526442 647320
rect 526498 647264 529092 647320
rect 526437 647262 529092 647264
rect 13721 647259 13787 647262
rect 41321 647259 41387 647262
rect 95141 647259 95207 647262
rect 122741 647259 122807 647262
rect 148961 647259 149027 647262
rect 202781 647259 202847 647262
rect 230381 647259 230447 647262
rect 256601 647259 256667 647262
rect 311801 647259 311867 647262
rect 338021 647259 338087 647262
rect 365621 647259 365687 647262
rect 391841 647259 391907 647262
rect 419441 647259 419507 647262
rect 445661 647259 445727 647262
rect 500861 647259 500927 647262
rect 526437 647259 526503 647262
rect 146293 647186 146359 647189
rect 253933 647186 253999 647189
rect 361573 647186 361639 647189
rect 469213 647186 469279 647189
rect 143766 647184 146359 647186
rect 143766 647128 146298 647184
rect 146354 647128 146359 647184
rect 143766 647126 146359 647128
rect 64873 646642 64939 646645
rect 91093 646642 91159 646645
rect 118693 646642 118759 646645
rect 62836 646640 64939 646642
rect 62836 646584 64878 646640
rect 64934 646584 64939 646640
rect 62836 646582 64939 646584
rect 89884 646640 91159 646642
rect 89884 646584 91098 646640
rect 91154 646584 91159 646640
rect 89884 646582 91159 646584
rect 116932 646640 118759 646642
rect 116932 646584 118698 646640
rect 118754 646584 118759 646640
rect 143766 646612 143826 647126
rect 146293 647123 146359 647126
rect 251774 647184 253999 647186
rect 251774 647128 253938 647184
rect 253994 647128 253999 647184
rect 251774 647126 253999 647128
rect 172513 646642 172579 646645
rect 200113 646642 200179 646645
rect 226333 646642 226399 646645
rect 170844 646640 172579 646642
rect 116932 646582 118759 646584
rect 170844 646584 172518 646640
rect 172574 646584 172579 646640
rect 170844 646582 172579 646584
rect 197892 646640 200179 646642
rect 197892 646584 200118 646640
rect 200174 646584 200179 646640
rect 197892 646582 200179 646584
rect 224940 646640 226399 646642
rect 224940 646584 226338 646640
rect 226394 646584 226399 646640
rect 251774 646612 251834 647126
rect 253933 647123 253999 647126
rect 359782 647184 361639 647186
rect 359782 647128 361578 647184
rect 361634 647128 361639 647184
rect 359782 647126 361639 647128
rect 280153 646642 280219 646645
rect 307753 646642 307819 646645
rect 335353 646642 335419 646645
rect 278852 646640 280219 646642
rect 224940 646582 226399 646584
rect 278852 646584 280158 646640
rect 280214 646584 280219 646640
rect 278852 646582 280219 646584
rect 305900 646640 307819 646642
rect 305900 646584 307758 646640
rect 307814 646584 307819 646640
rect 305900 646582 307819 646584
rect 332948 646640 335419 646642
rect 332948 646584 335358 646640
rect 335414 646584 335419 646640
rect 359782 646612 359842 647126
rect 361573 647123 361639 647126
rect 467790 647184 469279 647186
rect 467790 647128 469218 647184
rect 469274 647128 469279 647184
rect 467790 647126 469279 647128
rect 389173 646642 389239 646645
rect 415393 646642 415459 646645
rect 442993 646642 443059 646645
rect 386860 646640 389239 646642
rect 332948 646582 335419 646584
rect 386860 646584 389178 646640
rect 389234 646584 389239 646640
rect 386860 646582 389239 646584
rect 413908 646640 415459 646642
rect 413908 646584 415398 646640
rect 415454 646584 415459 646640
rect 413908 646582 415459 646584
rect 440956 646640 443059 646642
rect 440956 646584 442998 646640
rect 443054 646584 443059 646640
rect 467790 646612 467850 647126
rect 469213 647123 469279 647126
rect 496813 646642 496879 646645
rect 523033 646642 523099 646645
rect 550633 646642 550699 646645
rect 494868 646640 496879 646642
rect 440956 646582 443059 646584
rect 494868 646584 496818 646640
rect 496874 646584 496879 646640
rect 494868 646582 496879 646584
rect 521916 646640 523099 646642
rect 521916 646584 523038 646640
rect 523094 646584 523099 646640
rect 521916 646582 523099 646584
rect 548964 646640 550699 646642
rect 548964 646584 550638 646640
rect 550694 646584 550699 646640
rect 548964 646582 550699 646584
rect 64873 646579 64939 646582
rect 91093 646579 91159 646582
rect 118693 646579 118759 646582
rect 172513 646579 172579 646582
rect 200113 646579 200179 646582
rect 226333 646579 226399 646582
rect 280153 646579 280219 646582
rect 307753 646579 307819 646582
rect 335353 646579 335419 646582
rect 389173 646579 389239 646582
rect 415393 646579 415459 646582
rect 442993 646579 443059 646582
rect 496813 646579 496879 646582
rect 523033 646579 523099 646582
rect 550633 646579 550699 646582
rect 35758 645962 35818 646476
rect 37917 645962 37983 645965
rect 35758 645960 37983 645962
rect 35758 645904 37922 645960
rect 37978 645904 37983 645960
rect 35758 645902 37983 645904
rect 37917 645899 37983 645902
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect 526437 620394 526503 620397
rect 526437 620392 529092 620394
rect 526437 620336 526442 620392
rect 526498 620336 529092 620392
rect 526437 620334 529092 620336
rect 526437 620331 526503 620334
rect 13721 620258 13787 620261
rect 41321 620258 41387 620261
rect 95141 620258 95207 620261
rect 122741 620258 122807 620261
rect 148961 620258 149027 620261
rect 202781 620258 202847 620261
rect 230381 620258 230447 620261
rect 256601 620258 256667 620261
rect 311801 620258 311867 620261
rect 338021 620258 338087 620261
rect 365621 620258 365687 620261
rect 391841 620258 391907 620261
rect 419441 620258 419507 620261
rect 445661 620258 445727 620261
rect 500861 620258 500927 620261
rect 13721 620256 16100 620258
rect 13721 620200 13726 620256
rect 13782 620200 16100 620256
rect 13721 620198 16100 620200
rect 41321 620256 43148 620258
rect 41321 620200 41326 620256
rect 41382 620200 43148 620256
rect 95141 620256 97060 620258
rect 41321 620198 43148 620200
rect 13721 620195 13787 620198
rect 41321 620195 41387 620198
rect 68921 619714 68987 619717
rect 70166 619714 70226 620228
rect 95141 620200 95146 620256
rect 95202 620200 97060 620256
rect 95141 620198 97060 620200
rect 122741 620256 124108 620258
rect 122741 620200 122746 620256
rect 122802 620200 124108 620256
rect 122741 620198 124108 620200
rect 148961 620256 151156 620258
rect 148961 620200 148966 620256
rect 149022 620200 151156 620256
rect 202781 620256 205068 620258
rect 148961 620198 151156 620200
rect 95141 620195 95207 620198
rect 122741 620195 122807 620198
rect 148961 620195 149027 620198
rect 68921 619712 70226 619714
rect 68921 619656 68926 619712
rect 68982 619656 70226 619712
rect 68921 619654 70226 619656
rect 176561 619714 176627 619717
rect 178174 619714 178234 620228
rect 202781 620200 202786 620256
rect 202842 620200 205068 620256
rect 202781 620198 205068 620200
rect 230381 620256 232116 620258
rect 230381 620200 230386 620256
rect 230442 620200 232116 620256
rect 230381 620198 232116 620200
rect 256601 620256 259164 620258
rect 256601 620200 256606 620256
rect 256662 620200 259164 620256
rect 311801 620256 313076 620258
rect 256601 620198 259164 620200
rect 202781 620195 202847 620198
rect 230381 620195 230447 620198
rect 256601 620195 256667 620198
rect 176561 619712 178234 619714
rect 176561 619656 176566 619712
rect 176622 619656 178234 619712
rect 176561 619654 178234 619656
rect 284201 619714 284267 619717
rect 286182 619714 286242 620228
rect 311801 620200 311806 620256
rect 311862 620200 313076 620256
rect 311801 620198 313076 620200
rect 338021 620256 340124 620258
rect 338021 620200 338026 620256
rect 338082 620200 340124 620256
rect 338021 620198 340124 620200
rect 365621 620256 367172 620258
rect 365621 620200 365626 620256
rect 365682 620200 367172 620256
rect 365621 620198 367172 620200
rect 391841 620256 394036 620258
rect 391841 620200 391846 620256
rect 391902 620200 394036 620256
rect 391841 620198 394036 620200
rect 419441 620256 421084 620258
rect 419441 620200 419446 620256
rect 419502 620200 421084 620256
rect 419441 620198 421084 620200
rect 445661 620256 448132 620258
rect 445661 620200 445666 620256
rect 445722 620200 448132 620256
rect 500861 620256 502044 620258
rect 445661 620198 448132 620200
rect 311801 620195 311867 620198
rect 338021 620195 338087 620198
rect 365621 620195 365687 620198
rect 391841 620195 391907 620198
rect 419441 620195 419507 620198
rect 445661 620195 445727 620198
rect 284201 619712 286242 619714
rect 284201 619656 284206 619712
rect 284262 619656 286242 619712
rect 284201 619654 286242 619656
rect 473261 619714 473327 619717
rect 475150 619714 475210 620228
rect 500861 620200 500866 620256
rect 500922 620200 502044 620256
rect 500861 620198 502044 620200
rect 500861 620195 500927 620198
rect 473261 619712 475210 619714
rect 473261 619656 473266 619712
rect 473322 619656 475210 619712
rect 473261 619654 475210 619656
rect 68921 619651 68987 619654
rect 176561 619651 176627 619654
rect 284201 619651 284267 619654
rect 473261 619651 473327 619654
rect 64873 619578 64939 619581
rect 91093 619578 91159 619581
rect 118693 619578 118759 619581
rect 172513 619578 172579 619581
rect 200113 619578 200179 619581
rect 226333 619578 226399 619581
rect 280153 619578 280219 619581
rect 307753 619578 307819 619581
rect 335353 619578 335419 619581
rect 389173 619578 389239 619581
rect 415393 619578 415459 619581
rect 442993 619578 443059 619581
rect 496813 619578 496879 619581
rect 523033 619578 523099 619581
rect 550633 619578 550699 619581
rect 62836 619576 64939 619578
rect -960 619020 480 619260
rect 35758 619034 35818 619548
rect 62836 619520 64878 619576
rect 64934 619520 64939 619576
rect 62836 619518 64939 619520
rect 89884 619576 91159 619578
rect 89884 619520 91098 619576
rect 91154 619520 91159 619576
rect 89884 619518 91159 619520
rect 116932 619576 118759 619578
rect 116932 619520 118698 619576
rect 118754 619520 118759 619576
rect 170844 619576 172579 619578
rect 116932 619518 118759 619520
rect 64873 619515 64939 619518
rect 91093 619515 91159 619518
rect 118693 619515 118759 619518
rect 37917 619034 37983 619037
rect 35758 619032 37983 619034
rect 35758 618976 37922 619032
rect 37978 618976 37983 619032
rect 35758 618974 37983 618976
rect 143766 619034 143826 619548
rect 170844 619520 172518 619576
rect 172574 619520 172579 619576
rect 170844 619518 172579 619520
rect 197892 619576 200179 619578
rect 197892 619520 200118 619576
rect 200174 619520 200179 619576
rect 197892 619518 200179 619520
rect 224940 619576 226399 619578
rect 224940 619520 226338 619576
rect 226394 619520 226399 619576
rect 278852 619576 280219 619578
rect 224940 619518 226399 619520
rect 172513 619515 172579 619518
rect 200113 619515 200179 619518
rect 226333 619515 226399 619518
rect 146293 619034 146359 619037
rect 143766 619032 146359 619034
rect 143766 618976 146298 619032
rect 146354 618976 146359 619032
rect 143766 618974 146359 618976
rect 251774 619034 251834 619548
rect 278852 619520 280158 619576
rect 280214 619520 280219 619576
rect 278852 619518 280219 619520
rect 305900 619576 307819 619578
rect 305900 619520 307758 619576
rect 307814 619520 307819 619576
rect 305900 619518 307819 619520
rect 332948 619576 335419 619578
rect 332948 619520 335358 619576
rect 335414 619520 335419 619576
rect 386860 619576 389239 619578
rect 332948 619518 335419 619520
rect 280153 619515 280219 619518
rect 307753 619515 307819 619518
rect 335353 619515 335419 619518
rect 253933 619034 253999 619037
rect 251774 619032 253999 619034
rect 251774 618976 253938 619032
rect 253994 618976 253999 619032
rect 251774 618974 253999 618976
rect 359782 619034 359842 619548
rect 386860 619520 389178 619576
rect 389234 619520 389239 619576
rect 386860 619518 389239 619520
rect 413908 619576 415459 619578
rect 413908 619520 415398 619576
rect 415454 619520 415459 619576
rect 413908 619518 415459 619520
rect 440956 619576 443059 619578
rect 440956 619520 442998 619576
rect 443054 619520 443059 619576
rect 494868 619576 496879 619578
rect 440956 619518 443059 619520
rect 389173 619515 389239 619518
rect 415393 619515 415459 619518
rect 442993 619515 443059 619518
rect 361573 619034 361639 619037
rect 359782 619032 361639 619034
rect 359782 618976 361578 619032
rect 361634 618976 361639 619032
rect 359782 618974 361639 618976
rect 467790 619034 467850 619548
rect 494868 619520 496818 619576
rect 496874 619520 496879 619576
rect 494868 619518 496879 619520
rect 521916 619576 523099 619578
rect 521916 619520 523038 619576
rect 523094 619520 523099 619576
rect 521916 619518 523099 619520
rect 548964 619576 550699 619578
rect 548964 619520 550638 619576
rect 550694 619520 550699 619576
rect 548964 619518 550699 619520
rect 496813 619515 496879 619518
rect 523033 619515 523099 619518
rect 550633 619515 550699 619518
rect 469213 619034 469279 619037
rect 467790 619032 469279 619034
rect 467790 618976 469218 619032
rect 469274 618976 469279 619032
rect 467790 618974 469279 618976
rect 37917 618971 37983 618974
rect 146293 618971 146359 618974
rect 253933 618971 253999 618974
rect 361573 618971 361639 618974
rect 469213 618971 469279 618974
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect 526437 593330 526503 593333
rect 526437 593328 529092 593330
rect 526437 593272 526442 593328
rect 526498 593272 529092 593328
rect 526437 593270 529092 593272
rect 526437 593267 526503 593270
rect 13721 593194 13787 593197
rect 41321 593194 41387 593197
rect 95141 593194 95207 593197
rect 122741 593194 122807 593197
rect 148961 593194 149027 593197
rect 202781 593194 202847 593197
rect 230381 593194 230447 593197
rect 256601 593194 256667 593197
rect 311801 593194 311867 593197
rect 338021 593194 338087 593197
rect 365621 593194 365687 593197
rect 419441 593194 419507 593197
rect 445661 593194 445727 593197
rect 500861 593194 500927 593197
rect 13721 593192 16100 593194
rect -960 592908 480 593148
rect 13721 593136 13726 593192
rect 13782 593136 16100 593192
rect 13721 593134 16100 593136
rect 41321 593192 43148 593194
rect 41321 593136 41326 593192
rect 41382 593136 43148 593192
rect 95141 593192 97060 593194
rect 41321 593134 43148 593136
rect 13721 593131 13787 593134
rect 41321 593131 41387 593134
rect 68921 592650 68987 592653
rect 70166 592650 70226 593164
rect 95141 593136 95146 593192
rect 95202 593136 97060 593192
rect 95141 593134 97060 593136
rect 122741 593192 124108 593194
rect 122741 593136 122746 593192
rect 122802 593136 124108 593192
rect 122741 593134 124108 593136
rect 148961 593192 151156 593194
rect 148961 593136 148966 593192
rect 149022 593136 151156 593192
rect 202781 593192 205068 593194
rect 148961 593134 151156 593136
rect 95141 593131 95207 593134
rect 122741 593131 122807 593134
rect 148961 593131 149027 593134
rect 68921 592648 70226 592650
rect 68921 592592 68926 592648
rect 68982 592592 70226 592648
rect 68921 592590 70226 592592
rect 176561 592650 176627 592653
rect 178174 592650 178234 593164
rect 202781 593136 202786 593192
rect 202842 593136 205068 593192
rect 202781 593134 205068 593136
rect 230381 593192 232116 593194
rect 230381 593136 230386 593192
rect 230442 593136 232116 593192
rect 230381 593134 232116 593136
rect 256601 593192 259164 593194
rect 256601 593136 256606 593192
rect 256662 593136 259164 593192
rect 311801 593192 313076 593194
rect 256601 593134 259164 593136
rect 202781 593131 202847 593134
rect 230381 593131 230447 593134
rect 256601 593131 256667 593134
rect 176561 592648 178234 592650
rect 176561 592592 176566 592648
rect 176622 592592 178234 592648
rect 176561 592590 178234 592592
rect 284201 592650 284267 592653
rect 286182 592650 286242 593164
rect 311801 593136 311806 593192
rect 311862 593136 313076 593192
rect 311801 593134 313076 593136
rect 338021 593192 340124 593194
rect 338021 593136 338026 593192
rect 338082 593136 340124 593192
rect 338021 593134 340124 593136
rect 365621 593192 367172 593194
rect 365621 593136 365626 593192
rect 365682 593136 367172 593192
rect 419441 593192 421084 593194
rect 365621 593134 367172 593136
rect 311801 593131 311867 593134
rect 338021 593131 338087 593134
rect 365621 593131 365687 593134
rect 284201 592648 286242 592650
rect 284201 592592 284206 592648
rect 284262 592592 286242 592648
rect 284201 592590 286242 592592
rect 391841 592650 391907 592653
rect 394006 592650 394066 593164
rect 419441 593136 419446 593192
rect 419502 593136 421084 593192
rect 419441 593134 421084 593136
rect 445661 593192 448132 593194
rect 445661 593136 445666 593192
rect 445722 593136 448132 593192
rect 500861 593192 502044 593194
rect 445661 593134 448132 593136
rect 419441 593131 419507 593134
rect 445661 593131 445727 593134
rect 391841 592648 394066 592650
rect 391841 592592 391846 592648
rect 391902 592592 394066 592648
rect 391841 592590 394066 592592
rect 473261 592650 473327 592653
rect 475150 592650 475210 593164
rect 500861 593136 500866 593192
rect 500922 593136 502044 593192
rect 500861 593134 502044 593136
rect 500861 593131 500927 593134
rect 473261 592648 475210 592650
rect 473261 592592 473266 592648
rect 473322 592592 475210 592648
rect 473261 592590 475210 592592
rect 68921 592587 68987 592590
rect 176561 592587 176627 592590
rect 284201 592587 284267 592590
rect 391841 592587 391907 592590
rect 473261 592587 473327 592590
rect 64873 592514 64939 592517
rect 91093 592514 91159 592517
rect 118693 592514 118759 592517
rect 172513 592514 172579 592517
rect 200113 592514 200179 592517
rect 226333 592514 226399 592517
rect 280153 592514 280219 592517
rect 307753 592514 307819 592517
rect 335353 592514 335419 592517
rect 389173 592514 389239 592517
rect 415393 592514 415459 592517
rect 442993 592514 443059 592517
rect 496813 592514 496879 592517
rect 523033 592514 523099 592517
rect 62836 592512 64939 592514
rect 35758 592106 35818 592484
rect 62836 592456 64878 592512
rect 64934 592456 64939 592512
rect 62836 592454 64939 592456
rect 89884 592512 91159 592514
rect 89884 592456 91098 592512
rect 91154 592456 91159 592512
rect 89884 592454 91159 592456
rect 116932 592512 118759 592514
rect 116932 592456 118698 592512
rect 118754 592456 118759 592512
rect 170844 592512 172579 592514
rect 116932 592454 118759 592456
rect 64873 592451 64939 592454
rect 91093 592451 91159 592454
rect 118693 592451 118759 592454
rect 37917 592106 37983 592109
rect 35758 592104 37983 592106
rect 35758 592048 37922 592104
rect 37978 592048 37983 592104
rect 35758 592046 37983 592048
rect 143766 592106 143826 592484
rect 170844 592456 172518 592512
rect 172574 592456 172579 592512
rect 170844 592454 172579 592456
rect 197892 592512 200179 592514
rect 197892 592456 200118 592512
rect 200174 592456 200179 592512
rect 197892 592454 200179 592456
rect 224940 592512 226399 592514
rect 224940 592456 226338 592512
rect 226394 592456 226399 592512
rect 278852 592512 280219 592514
rect 224940 592454 226399 592456
rect 172513 592451 172579 592454
rect 200113 592451 200179 592454
rect 226333 592451 226399 592454
rect 146293 592106 146359 592109
rect 143766 592104 146359 592106
rect 143766 592048 146298 592104
rect 146354 592048 146359 592104
rect 143766 592046 146359 592048
rect 251774 592106 251834 592484
rect 278852 592456 280158 592512
rect 280214 592456 280219 592512
rect 278852 592454 280219 592456
rect 305900 592512 307819 592514
rect 305900 592456 307758 592512
rect 307814 592456 307819 592512
rect 305900 592454 307819 592456
rect 332948 592512 335419 592514
rect 332948 592456 335358 592512
rect 335414 592456 335419 592512
rect 386860 592512 389239 592514
rect 332948 592454 335419 592456
rect 280153 592451 280219 592454
rect 307753 592451 307819 592454
rect 335353 592451 335419 592454
rect 253933 592106 253999 592109
rect 251774 592104 253999 592106
rect 251774 592048 253938 592104
rect 253994 592048 253999 592104
rect 251774 592046 253999 592048
rect 359782 592106 359842 592484
rect 386860 592456 389178 592512
rect 389234 592456 389239 592512
rect 386860 592454 389239 592456
rect 413908 592512 415459 592514
rect 413908 592456 415398 592512
rect 415454 592456 415459 592512
rect 413908 592454 415459 592456
rect 440956 592512 443059 592514
rect 440956 592456 442998 592512
rect 443054 592456 443059 592512
rect 494868 592512 496879 592514
rect 440956 592454 443059 592456
rect 389173 592451 389239 592454
rect 415393 592451 415459 592454
rect 442993 592451 443059 592454
rect 361573 592106 361639 592109
rect 359782 592104 361639 592106
rect 359782 592048 361578 592104
rect 361634 592048 361639 592104
rect 359782 592046 361639 592048
rect 467790 592106 467850 592484
rect 494868 592456 496818 592512
rect 496874 592456 496879 592512
rect 494868 592454 496879 592456
rect 521916 592512 523099 592514
rect 521916 592456 523038 592512
rect 523094 592456 523099 592512
rect 521916 592454 523099 592456
rect 496813 592451 496879 592454
rect 523033 592451 523099 592454
rect 469213 592106 469279 592109
rect 467790 592104 469279 592106
rect 467790 592048 469218 592104
rect 469274 592048 469279 592104
rect 467790 592046 469279 592048
rect 548934 592106 548994 592484
rect 550633 592106 550699 592109
rect 548934 592104 550699 592106
rect 548934 592048 550638 592104
rect 550694 592048 550699 592104
rect 548934 592046 550699 592048
rect 37917 592043 37983 592046
rect 146293 592043 146359 592046
rect 253933 592043 253999 592046
rect 361573 592043 361639 592046
rect 469213 592043 469279 592046
rect 550633 592043 550699 592046
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 526437 566402 526503 566405
rect 526437 566400 529092 566402
rect 526437 566344 526442 566400
rect 526498 566344 529092 566400
rect 526437 566342 529092 566344
rect 526437 566339 526503 566342
rect 13721 566266 13787 566269
rect 41321 566266 41387 566269
rect 95141 566266 95207 566269
rect 122741 566266 122807 566269
rect 148961 566266 149027 566269
rect 202781 566266 202847 566269
rect 230381 566266 230447 566269
rect 256601 566266 256667 566269
rect 311801 566266 311867 566269
rect 338021 566266 338087 566269
rect 365621 566266 365687 566269
rect 391841 566266 391907 566269
rect 419441 566266 419507 566269
rect 445661 566266 445727 566269
rect 500861 566266 500927 566269
rect 13721 566264 16100 566266
rect 13721 566208 13726 566264
rect 13782 566208 16100 566264
rect 13721 566206 16100 566208
rect 41321 566264 43148 566266
rect 41321 566208 41326 566264
rect 41382 566208 43148 566264
rect 95141 566264 97060 566266
rect 41321 566206 43148 566208
rect 13721 566203 13787 566206
rect 41321 566203 41387 566206
rect 68921 565858 68987 565861
rect 70166 565858 70226 566236
rect 95141 566208 95146 566264
rect 95202 566208 97060 566264
rect 95141 566206 97060 566208
rect 122741 566264 124108 566266
rect 122741 566208 122746 566264
rect 122802 566208 124108 566264
rect 122741 566206 124108 566208
rect 148961 566264 151156 566266
rect 148961 566208 148966 566264
rect 149022 566208 151156 566264
rect 202781 566264 205068 566266
rect 148961 566206 151156 566208
rect 95141 566203 95207 566206
rect 122741 566203 122807 566206
rect 148961 566203 149027 566206
rect 68921 565856 70226 565858
rect 68921 565800 68926 565856
rect 68982 565800 70226 565856
rect 68921 565798 70226 565800
rect 176561 565858 176627 565861
rect 178174 565858 178234 566236
rect 202781 566208 202786 566264
rect 202842 566208 205068 566264
rect 202781 566206 205068 566208
rect 230381 566264 232116 566266
rect 230381 566208 230386 566264
rect 230442 566208 232116 566264
rect 230381 566206 232116 566208
rect 256601 566264 259164 566266
rect 256601 566208 256606 566264
rect 256662 566208 259164 566264
rect 311801 566264 313076 566266
rect 256601 566206 259164 566208
rect 202781 566203 202847 566206
rect 230381 566203 230447 566206
rect 256601 566203 256667 566206
rect 176561 565856 178234 565858
rect 176561 565800 176566 565856
rect 176622 565800 178234 565856
rect 176561 565798 178234 565800
rect 284201 565858 284267 565861
rect 286182 565858 286242 566236
rect 311801 566208 311806 566264
rect 311862 566208 313076 566264
rect 311801 566206 313076 566208
rect 338021 566264 340124 566266
rect 338021 566208 338026 566264
rect 338082 566208 340124 566264
rect 338021 566206 340124 566208
rect 365621 566264 367172 566266
rect 365621 566208 365626 566264
rect 365682 566208 367172 566264
rect 365621 566206 367172 566208
rect 391841 566264 394036 566266
rect 391841 566208 391846 566264
rect 391902 566208 394036 566264
rect 391841 566206 394036 566208
rect 419441 566264 421084 566266
rect 419441 566208 419446 566264
rect 419502 566208 421084 566264
rect 419441 566206 421084 566208
rect 445661 566264 448132 566266
rect 445661 566208 445666 566264
rect 445722 566208 448132 566264
rect 500861 566264 502044 566266
rect 445661 566206 448132 566208
rect 311801 566203 311867 566206
rect 338021 566203 338087 566206
rect 365621 566203 365687 566206
rect 391841 566203 391907 566206
rect 419441 566203 419507 566206
rect 445661 566203 445727 566206
rect 284201 565856 286242 565858
rect 284201 565800 284206 565856
rect 284262 565800 286242 565856
rect 284201 565798 286242 565800
rect 473261 565858 473327 565861
rect 475150 565858 475210 566236
rect 500861 566208 500866 566264
rect 500922 566208 502044 566264
rect 500861 566206 502044 566208
rect 500861 566203 500927 566206
rect 473261 565856 475210 565858
rect 473261 565800 473266 565856
rect 473322 565800 475210 565856
rect 473261 565798 475210 565800
rect 68921 565795 68987 565798
rect 176561 565795 176627 565798
rect 284201 565795 284267 565798
rect 473261 565795 473327 565798
rect 64873 565586 64939 565589
rect 91093 565586 91159 565589
rect 118693 565586 118759 565589
rect 172513 565586 172579 565589
rect 200113 565586 200179 565589
rect 226333 565586 226399 565589
rect 280153 565586 280219 565589
rect 307753 565586 307819 565589
rect 335353 565586 335419 565589
rect 389173 565586 389239 565589
rect 415393 565586 415459 565589
rect 442993 565586 443059 565589
rect 496813 565586 496879 565589
rect 523033 565586 523099 565589
rect 550633 565586 550699 565589
rect 62836 565584 64939 565586
rect 35758 565042 35818 565556
rect 62836 565528 64878 565584
rect 64934 565528 64939 565584
rect 62836 565526 64939 565528
rect 89884 565584 91159 565586
rect 89884 565528 91098 565584
rect 91154 565528 91159 565584
rect 89884 565526 91159 565528
rect 116932 565584 118759 565586
rect 116932 565528 118698 565584
rect 118754 565528 118759 565584
rect 170844 565584 172579 565586
rect 116932 565526 118759 565528
rect 64873 565523 64939 565526
rect 91093 565523 91159 565526
rect 118693 565523 118759 565526
rect 37917 565042 37983 565045
rect 35758 565040 37983 565042
rect 35758 564984 37922 565040
rect 37978 564984 37983 565040
rect 35758 564982 37983 564984
rect 143766 565042 143826 565556
rect 170844 565528 172518 565584
rect 172574 565528 172579 565584
rect 170844 565526 172579 565528
rect 197892 565584 200179 565586
rect 197892 565528 200118 565584
rect 200174 565528 200179 565584
rect 197892 565526 200179 565528
rect 224940 565584 226399 565586
rect 224940 565528 226338 565584
rect 226394 565528 226399 565584
rect 278852 565584 280219 565586
rect 224940 565526 226399 565528
rect 172513 565523 172579 565526
rect 200113 565523 200179 565526
rect 226333 565523 226399 565526
rect 146293 565042 146359 565045
rect 143766 565040 146359 565042
rect 143766 564984 146298 565040
rect 146354 564984 146359 565040
rect 143766 564982 146359 564984
rect 251774 565042 251834 565556
rect 278852 565528 280158 565584
rect 280214 565528 280219 565584
rect 278852 565526 280219 565528
rect 305900 565584 307819 565586
rect 305900 565528 307758 565584
rect 307814 565528 307819 565584
rect 305900 565526 307819 565528
rect 332948 565584 335419 565586
rect 332948 565528 335358 565584
rect 335414 565528 335419 565584
rect 386860 565584 389239 565586
rect 332948 565526 335419 565528
rect 280153 565523 280219 565526
rect 307753 565523 307819 565526
rect 335353 565523 335419 565526
rect 253933 565042 253999 565045
rect 251774 565040 253999 565042
rect 251774 564984 253938 565040
rect 253994 564984 253999 565040
rect 251774 564982 253999 564984
rect 359782 565042 359842 565556
rect 386860 565528 389178 565584
rect 389234 565528 389239 565584
rect 386860 565526 389239 565528
rect 413908 565584 415459 565586
rect 413908 565528 415398 565584
rect 415454 565528 415459 565584
rect 413908 565526 415459 565528
rect 440956 565584 443059 565586
rect 440956 565528 442998 565584
rect 443054 565528 443059 565584
rect 494868 565584 496879 565586
rect 440956 565526 443059 565528
rect 389173 565523 389239 565526
rect 415393 565523 415459 565526
rect 442993 565523 443059 565526
rect 361573 565042 361639 565045
rect 359782 565040 361639 565042
rect 359782 564984 361578 565040
rect 361634 564984 361639 565040
rect 359782 564982 361639 564984
rect 467790 565042 467850 565556
rect 494868 565528 496818 565584
rect 496874 565528 496879 565584
rect 494868 565526 496879 565528
rect 521916 565584 523099 565586
rect 521916 565528 523038 565584
rect 523094 565528 523099 565584
rect 521916 565526 523099 565528
rect 548964 565584 550699 565586
rect 548964 565528 550638 565584
rect 550694 565528 550699 565584
rect 548964 565526 550699 565528
rect 496813 565523 496879 565526
rect 523033 565523 523099 565526
rect 550633 565523 550699 565526
rect 469213 565042 469279 565045
rect 467790 565040 469279 565042
rect 467790 564984 469218 565040
rect 469274 564984 469279 565040
rect 467790 564982 469279 564984
rect 37917 564979 37983 564982
rect 146293 564979 146359 564982
rect 253933 564979 253999 564982
rect 361573 564979 361639 564982
rect 469213 564979 469279 564982
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 526437 539338 526503 539341
rect 526437 539336 529092 539338
rect 526437 539280 526442 539336
rect 526498 539280 529092 539336
rect 526437 539278 529092 539280
rect 526437 539275 526503 539278
rect 13721 539202 13787 539205
rect 41321 539202 41387 539205
rect 95141 539202 95207 539205
rect 122741 539202 122807 539205
rect 148961 539202 149027 539205
rect 202781 539202 202847 539205
rect 230381 539202 230447 539205
rect 256601 539202 256667 539205
rect 311801 539202 311867 539205
rect 338021 539202 338087 539205
rect 365621 539202 365687 539205
rect 391841 539202 391907 539205
rect 419441 539202 419507 539205
rect 445661 539202 445727 539205
rect 500861 539202 500927 539205
rect 13721 539200 16100 539202
rect 13721 539144 13726 539200
rect 13782 539144 16100 539200
rect 13721 539142 16100 539144
rect 41321 539200 43148 539202
rect 41321 539144 41326 539200
rect 41382 539144 43148 539200
rect 95141 539200 97060 539202
rect 41321 539142 43148 539144
rect 13721 539139 13787 539142
rect 41321 539139 41387 539142
rect 68921 538658 68987 538661
rect 70166 538658 70226 539172
rect 95141 539144 95146 539200
rect 95202 539144 97060 539200
rect 95141 539142 97060 539144
rect 122741 539200 124108 539202
rect 122741 539144 122746 539200
rect 122802 539144 124108 539200
rect 122741 539142 124108 539144
rect 148961 539200 151156 539202
rect 148961 539144 148966 539200
rect 149022 539144 151156 539200
rect 202781 539200 205068 539202
rect 148961 539142 151156 539144
rect 95141 539139 95207 539142
rect 122741 539139 122807 539142
rect 148961 539139 149027 539142
rect 68921 538656 70226 538658
rect 68921 538600 68926 538656
rect 68982 538600 70226 538656
rect 68921 538598 70226 538600
rect 176561 538658 176627 538661
rect 178174 538658 178234 539172
rect 202781 539144 202786 539200
rect 202842 539144 205068 539200
rect 202781 539142 205068 539144
rect 230381 539200 232116 539202
rect 230381 539144 230386 539200
rect 230442 539144 232116 539200
rect 230381 539142 232116 539144
rect 256601 539200 259164 539202
rect 256601 539144 256606 539200
rect 256662 539144 259164 539200
rect 311801 539200 313076 539202
rect 256601 539142 259164 539144
rect 202781 539139 202847 539142
rect 230381 539139 230447 539142
rect 256601 539139 256667 539142
rect 176561 538656 178234 538658
rect 176561 538600 176566 538656
rect 176622 538600 178234 538656
rect 176561 538598 178234 538600
rect 284201 538658 284267 538661
rect 286182 538658 286242 539172
rect 311801 539144 311806 539200
rect 311862 539144 313076 539200
rect 311801 539142 313076 539144
rect 338021 539200 340124 539202
rect 338021 539144 338026 539200
rect 338082 539144 340124 539200
rect 338021 539142 340124 539144
rect 365621 539200 367172 539202
rect 365621 539144 365626 539200
rect 365682 539144 367172 539200
rect 365621 539142 367172 539144
rect 391841 539200 394036 539202
rect 391841 539144 391846 539200
rect 391902 539144 394036 539200
rect 391841 539142 394036 539144
rect 419441 539200 421084 539202
rect 419441 539144 419446 539200
rect 419502 539144 421084 539200
rect 419441 539142 421084 539144
rect 445661 539200 448132 539202
rect 445661 539144 445666 539200
rect 445722 539144 448132 539200
rect 500861 539200 502044 539202
rect 445661 539142 448132 539144
rect 311801 539139 311867 539142
rect 338021 539139 338087 539142
rect 365621 539139 365687 539142
rect 391841 539139 391907 539142
rect 419441 539139 419507 539142
rect 445661 539139 445727 539142
rect 284201 538656 286242 538658
rect 284201 538600 284206 538656
rect 284262 538600 286242 538656
rect 284201 538598 286242 538600
rect 473261 538658 473327 538661
rect 475150 538658 475210 539172
rect 500861 539144 500866 539200
rect 500922 539144 502044 539200
rect 500861 539142 502044 539144
rect 500861 539139 500927 539142
rect 473261 538656 475210 538658
rect 473261 538600 473266 538656
rect 473322 538600 475210 538656
rect 473261 538598 475210 538600
rect 68921 538595 68987 538598
rect 176561 538595 176627 538598
rect 284201 538595 284267 538598
rect 473261 538595 473327 538598
rect 64873 538522 64939 538525
rect 91093 538522 91159 538525
rect 118693 538522 118759 538525
rect 172513 538522 172579 538525
rect 200113 538522 200179 538525
rect 226333 538522 226399 538525
rect 280153 538522 280219 538525
rect 307753 538522 307819 538525
rect 335353 538522 335419 538525
rect 389173 538522 389239 538525
rect 415393 538522 415459 538525
rect 442993 538522 443059 538525
rect 496813 538522 496879 538525
rect 523033 538522 523099 538525
rect 550633 538522 550699 538525
rect 62836 538520 64939 538522
rect 35758 538250 35818 538492
rect 62836 538464 64878 538520
rect 64934 538464 64939 538520
rect 62836 538462 64939 538464
rect 89884 538520 91159 538522
rect 89884 538464 91098 538520
rect 91154 538464 91159 538520
rect 89884 538462 91159 538464
rect 116932 538520 118759 538522
rect 116932 538464 118698 538520
rect 118754 538464 118759 538520
rect 170844 538520 172579 538522
rect 116932 538462 118759 538464
rect 64873 538459 64939 538462
rect 91093 538459 91159 538462
rect 118693 538459 118759 538462
rect 143766 538386 143826 538492
rect 170844 538464 172518 538520
rect 172574 538464 172579 538520
rect 170844 538462 172579 538464
rect 197892 538520 200179 538522
rect 197892 538464 200118 538520
rect 200174 538464 200179 538520
rect 197892 538462 200179 538464
rect 224940 538520 226399 538522
rect 224940 538464 226338 538520
rect 226394 538464 226399 538520
rect 278852 538520 280219 538522
rect 224940 538462 226399 538464
rect 172513 538459 172579 538462
rect 200113 538459 200179 538462
rect 226333 538459 226399 538462
rect 146293 538386 146359 538389
rect 143766 538384 146359 538386
rect 143766 538328 146298 538384
rect 146354 538328 146359 538384
rect 143766 538326 146359 538328
rect 251774 538386 251834 538492
rect 278852 538464 280158 538520
rect 280214 538464 280219 538520
rect 278852 538462 280219 538464
rect 305900 538520 307819 538522
rect 305900 538464 307758 538520
rect 307814 538464 307819 538520
rect 305900 538462 307819 538464
rect 332948 538520 335419 538522
rect 332948 538464 335358 538520
rect 335414 538464 335419 538520
rect 386860 538520 389239 538522
rect 332948 538462 335419 538464
rect 280153 538459 280219 538462
rect 307753 538459 307819 538462
rect 335353 538459 335419 538462
rect 253933 538386 253999 538389
rect 251774 538384 253999 538386
rect 251774 538328 253938 538384
rect 253994 538328 253999 538384
rect 251774 538326 253999 538328
rect 359782 538386 359842 538492
rect 386860 538464 389178 538520
rect 389234 538464 389239 538520
rect 386860 538462 389239 538464
rect 413908 538520 415459 538522
rect 413908 538464 415398 538520
rect 415454 538464 415459 538520
rect 413908 538462 415459 538464
rect 440956 538520 443059 538522
rect 440956 538464 442998 538520
rect 443054 538464 443059 538520
rect 494868 538520 496879 538522
rect 440956 538462 443059 538464
rect 389173 538459 389239 538462
rect 415393 538459 415459 538462
rect 442993 538459 443059 538462
rect 361573 538386 361639 538389
rect 359782 538384 361639 538386
rect 359782 538328 361578 538384
rect 361634 538328 361639 538384
rect 359782 538326 361639 538328
rect 467790 538386 467850 538492
rect 494868 538464 496818 538520
rect 496874 538464 496879 538520
rect 494868 538462 496879 538464
rect 521916 538520 523099 538522
rect 521916 538464 523038 538520
rect 523094 538464 523099 538520
rect 521916 538462 523099 538464
rect 548964 538520 550699 538522
rect 548964 538464 550638 538520
rect 550694 538464 550699 538520
rect 548964 538462 550699 538464
rect 496813 538459 496879 538462
rect 523033 538459 523099 538462
rect 550633 538459 550699 538462
rect 469213 538386 469279 538389
rect 467790 538384 469279 538386
rect 467790 538328 469218 538384
rect 469274 538328 469279 538384
rect 467790 538326 469279 538328
rect 146293 538323 146359 538326
rect 253933 538323 253999 538326
rect 361573 538323 361639 538326
rect 469213 538323 469279 538326
rect 37917 538250 37983 538253
rect 35758 538248 37983 538250
rect 35758 538192 37922 538248
rect 37978 538192 37983 538248
rect 35758 538190 37983 538192
rect 37917 538187 37983 538190
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 579797 524514 579863 524517
rect 583520 524514 584960 524604
rect 579797 524512 584960 524514
rect 579797 524456 579802 524512
rect 579858 524456 584960 524512
rect 579797 524454 584960 524456
rect 579797 524451 579863 524454
rect 583520 524364 584960 524454
rect -960 514708 480 514948
rect 68921 512954 68987 512957
rect 96889 512954 96955 512957
rect 176561 512954 176627 512957
rect 204897 512954 204963 512957
rect 284201 512954 284267 512957
rect 339861 512954 339927 512957
rect 391841 512954 391907 512957
rect 473261 512954 473327 512957
rect 500861 512954 500927 512957
rect 68921 512952 70226 512954
rect 68921 512896 68926 512952
rect 68982 512896 70226 512952
rect 68921 512894 70226 512896
rect 68921 512891 68987 512894
rect 13721 512410 13787 512413
rect 41321 512410 41387 512413
rect 13721 512408 16100 512410
rect 13721 512352 13726 512408
rect 13782 512352 16100 512408
rect 13721 512350 16100 512352
rect 41321 512408 43148 512410
rect 41321 512352 41326 512408
rect 41382 512352 43148 512408
rect 70166 512380 70226 512894
rect 96889 512952 97090 512954
rect 96889 512896 96894 512952
rect 96950 512896 97090 512952
rect 96889 512894 97090 512896
rect 96889 512891 96955 512894
rect 97030 512380 97090 512894
rect 176561 512952 178234 512954
rect 176561 512896 176566 512952
rect 176622 512896 178234 512952
rect 176561 512894 178234 512896
rect 176561 512891 176627 512894
rect 122741 512410 122807 512413
rect 148961 512410 149027 512413
rect 122741 512408 124108 512410
rect 41321 512350 43148 512352
rect 122741 512352 122746 512408
rect 122802 512352 124108 512408
rect 122741 512350 124108 512352
rect 148961 512408 151156 512410
rect 148961 512352 148966 512408
rect 149022 512352 151156 512408
rect 178174 512380 178234 512894
rect 204897 512952 205098 512954
rect 204897 512896 204902 512952
rect 204958 512896 205098 512952
rect 204897 512894 205098 512896
rect 204897 512891 204963 512894
rect 205038 512380 205098 512894
rect 284201 512952 286242 512954
rect 284201 512896 284206 512952
rect 284262 512896 286242 512952
rect 284201 512894 286242 512896
rect 284201 512891 284267 512894
rect 230381 512410 230447 512413
rect 256601 512410 256667 512413
rect 230381 512408 232116 512410
rect 148961 512350 151156 512352
rect 230381 512352 230386 512408
rect 230442 512352 232116 512408
rect 230381 512350 232116 512352
rect 256601 512408 259164 512410
rect 256601 512352 256606 512408
rect 256662 512352 259164 512408
rect 286182 512380 286242 512894
rect 339861 512952 340154 512954
rect 339861 512896 339866 512952
rect 339922 512896 340154 512952
rect 339861 512894 340154 512896
rect 339861 512891 339927 512894
rect 311801 512410 311867 512413
rect 311801 512408 313076 512410
rect 256601 512350 259164 512352
rect 311801 512352 311806 512408
rect 311862 512352 313076 512408
rect 340094 512380 340154 512894
rect 391841 512952 394066 512954
rect 391841 512896 391846 512952
rect 391902 512896 394066 512952
rect 391841 512894 394066 512896
rect 391841 512891 391907 512894
rect 365621 512410 365687 512413
rect 365621 512408 367172 512410
rect 311801 512350 313076 512352
rect 365621 512352 365626 512408
rect 365682 512352 367172 512408
rect 394006 512380 394066 512894
rect 473261 512952 475210 512954
rect 473261 512896 473266 512952
rect 473322 512896 475210 512952
rect 473261 512894 475210 512896
rect 473261 512891 473327 512894
rect 419441 512410 419507 512413
rect 445661 512410 445727 512413
rect 419441 512408 421084 512410
rect 365621 512350 367172 512352
rect 419441 512352 419446 512408
rect 419502 512352 421084 512408
rect 419441 512350 421084 512352
rect 445661 512408 448132 512410
rect 445661 512352 445666 512408
rect 445722 512352 448132 512408
rect 475150 512380 475210 512894
rect 500861 512952 502074 512954
rect 500861 512896 500866 512952
rect 500922 512896 502074 512952
rect 500861 512894 502074 512896
rect 500861 512891 500927 512894
rect 502014 512380 502074 512894
rect 526437 512410 526503 512413
rect 526437 512408 529092 512410
rect 445661 512350 448132 512352
rect 526437 512352 526442 512408
rect 526498 512352 529092 512408
rect 526437 512350 529092 512352
rect 13721 512347 13787 512350
rect 41321 512347 41387 512350
rect 122741 512347 122807 512350
rect 148961 512347 149027 512350
rect 230381 512347 230447 512350
rect 256601 512347 256667 512350
rect 311801 512347 311867 512350
rect 365621 512347 365687 512350
rect 419441 512347 419507 512350
rect 445661 512347 445727 512350
rect 526437 512347 526503 512350
rect 146293 512002 146359 512005
rect 253933 512002 253999 512005
rect 361573 512002 361639 512005
rect 469213 512002 469279 512005
rect 550633 512002 550699 512005
rect 143766 512000 146359 512002
rect 143766 511944 146298 512000
rect 146354 511944 146359 512000
rect 143766 511942 146359 511944
rect 64873 511730 64939 511733
rect 91093 511730 91159 511733
rect 118693 511730 118759 511733
rect 62836 511728 64939 511730
rect 62836 511672 64878 511728
rect 64934 511672 64939 511728
rect 62836 511670 64939 511672
rect 89884 511728 91159 511730
rect 89884 511672 91098 511728
rect 91154 511672 91159 511728
rect 89884 511670 91159 511672
rect 116932 511728 118759 511730
rect 116932 511672 118698 511728
rect 118754 511672 118759 511728
rect 143766 511700 143826 511942
rect 146293 511939 146359 511942
rect 251774 512000 253999 512002
rect 251774 511944 253938 512000
rect 253994 511944 253999 512000
rect 251774 511942 253999 511944
rect 172513 511730 172579 511733
rect 200113 511730 200179 511733
rect 226333 511730 226399 511733
rect 170844 511728 172579 511730
rect 116932 511670 118759 511672
rect 170844 511672 172518 511728
rect 172574 511672 172579 511728
rect 170844 511670 172579 511672
rect 197892 511728 200179 511730
rect 197892 511672 200118 511728
rect 200174 511672 200179 511728
rect 197892 511670 200179 511672
rect 224940 511728 226399 511730
rect 224940 511672 226338 511728
rect 226394 511672 226399 511728
rect 251774 511700 251834 511942
rect 253933 511939 253999 511942
rect 359782 512000 361639 512002
rect 359782 511944 361578 512000
rect 361634 511944 361639 512000
rect 359782 511942 361639 511944
rect 280153 511730 280219 511733
rect 307753 511730 307819 511733
rect 335353 511730 335419 511733
rect 278852 511728 280219 511730
rect 224940 511670 226399 511672
rect 278852 511672 280158 511728
rect 280214 511672 280219 511728
rect 278852 511670 280219 511672
rect 305900 511728 307819 511730
rect 305900 511672 307758 511728
rect 307814 511672 307819 511728
rect 305900 511670 307819 511672
rect 332948 511728 335419 511730
rect 332948 511672 335358 511728
rect 335414 511672 335419 511728
rect 359782 511700 359842 511942
rect 361573 511939 361639 511942
rect 467790 512000 469279 512002
rect 467790 511944 469218 512000
rect 469274 511944 469279 512000
rect 467790 511942 469279 511944
rect 442993 511866 443059 511869
rect 440926 511864 443059 511866
rect 440926 511808 442998 511864
rect 443054 511808 443059 511864
rect 440926 511806 443059 511808
rect 389173 511730 389239 511733
rect 415393 511730 415459 511733
rect 386860 511728 389239 511730
rect 332948 511670 335419 511672
rect 386860 511672 389178 511728
rect 389234 511672 389239 511728
rect 386860 511670 389239 511672
rect 413908 511728 415459 511730
rect 413908 511672 415398 511728
rect 415454 511672 415459 511728
rect 440926 511700 440986 511806
rect 442993 511803 443059 511806
rect 467790 511700 467850 511942
rect 469213 511939 469279 511942
rect 548934 512000 550699 512002
rect 548934 511944 550638 512000
rect 550694 511944 550699 512000
rect 548934 511942 550699 511944
rect 496813 511730 496879 511733
rect 523033 511730 523099 511733
rect 494868 511728 496879 511730
rect 413908 511670 415459 511672
rect 494868 511672 496818 511728
rect 496874 511672 496879 511728
rect 494868 511670 496879 511672
rect 521916 511728 523099 511730
rect 521916 511672 523038 511728
rect 523094 511672 523099 511728
rect 548934 511700 548994 511942
rect 550633 511939 550699 511942
rect 521916 511670 523099 511672
rect 64873 511667 64939 511670
rect 91093 511667 91159 511670
rect 118693 511667 118759 511670
rect 172513 511667 172579 511670
rect 200113 511667 200179 511670
rect 226333 511667 226399 511670
rect 280153 511667 280219 511670
rect 307753 511667 307819 511670
rect 335353 511667 335419 511670
rect 389173 511667 389239 511670
rect 415393 511667 415459 511670
rect 496813 511667 496879 511670
rect 523033 511667 523099 511670
rect 35758 511050 35818 511564
rect 580257 511322 580323 511325
rect 583520 511322 584960 511412
rect 580257 511320 584960 511322
rect 580257 511264 580262 511320
rect 580318 511264 584960 511320
rect 580257 511262 584960 511264
rect 580257 511259 580323 511262
rect 583520 511172 584960 511262
rect 37917 511050 37983 511053
rect 35758 511048 37983 511050
rect 35758 510992 37922 511048
rect 37978 510992 37983 511048
rect 35758 510990 37983 510992
rect 37917 510987 37983 510990
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 68921 485754 68987 485757
rect 284201 485754 284267 485757
rect 473261 485754 473327 485757
rect 68921 485752 70226 485754
rect 68921 485696 68926 485752
rect 68982 485696 70226 485752
rect 68921 485694 70226 485696
rect 68921 485691 68987 485694
rect 41321 485346 41387 485349
rect 41321 485344 43148 485346
rect 41321 485288 41326 485344
rect 41382 485288 43148 485344
rect 70166 485316 70226 485694
rect 284201 485752 286242 485754
rect 284201 485696 284206 485752
rect 284262 485696 286242 485752
rect 284201 485694 286242 485696
rect 284201 485691 284267 485694
rect 122741 485346 122807 485349
rect 148961 485346 149027 485349
rect 202781 485346 202847 485349
rect 230381 485346 230447 485349
rect 122741 485344 124108 485346
rect 41321 485286 43148 485288
rect 122741 485288 122746 485344
rect 122802 485288 124108 485344
rect 122741 485286 124108 485288
rect 148961 485344 151156 485346
rect 148961 485288 148966 485344
rect 149022 485288 151156 485344
rect 148961 485286 151156 485288
rect 202781 485344 205068 485346
rect 202781 485288 202786 485344
rect 202842 485288 205068 485344
rect 202781 485286 205068 485288
rect 230381 485344 232116 485346
rect 230381 485288 230386 485344
rect 230442 485288 232116 485344
rect 286182 485316 286242 485694
rect 473261 485752 475210 485754
rect 473261 485696 473266 485752
rect 473322 485696 475210 485752
rect 473261 485694 475210 485696
rect 473261 485691 473327 485694
rect 311801 485346 311867 485349
rect 365621 485346 365687 485349
rect 419441 485346 419507 485349
rect 311801 485344 313076 485346
rect 230381 485286 232116 485288
rect 311801 485288 311806 485344
rect 311862 485288 313076 485344
rect 311801 485286 313076 485288
rect 365621 485344 367172 485346
rect 365621 485288 365626 485344
rect 365682 485288 367172 485344
rect 365621 485286 367172 485288
rect 419441 485344 421084 485346
rect 419441 485288 419446 485344
rect 419502 485288 421084 485344
rect 475150 485316 475210 485694
rect 500861 485346 500927 485349
rect 526437 485346 526503 485349
rect 500861 485344 502044 485346
rect 419441 485286 421084 485288
rect 500861 485288 500866 485344
rect 500922 485288 502044 485344
rect 500861 485286 502044 485288
rect 526437 485344 529092 485346
rect 526437 485288 526442 485344
rect 526498 485288 529092 485344
rect 526437 485286 529092 485288
rect 41321 485283 41387 485286
rect 122741 485283 122807 485286
rect 148961 485283 149027 485286
rect 202781 485283 202847 485286
rect 230381 485283 230447 485286
rect 311801 485283 311867 485286
rect 365621 485283 365687 485286
rect 419441 485283 419507 485286
rect 500861 485283 500927 485286
rect 526437 485283 526503 485286
rect 13721 485210 13787 485213
rect 95141 485210 95207 485213
rect 253933 485210 253999 485213
rect 13721 485208 16100 485210
rect 13721 485152 13726 485208
rect 13782 485152 16100 485208
rect 13721 485150 16100 485152
rect 95141 485208 97060 485210
rect 95141 485152 95146 485208
rect 95202 485152 97060 485208
rect 251774 485208 253999 485210
rect 95141 485150 97060 485152
rect 13721 485147 13787 485150
rect 95141 485147 95207 485150
rect 37917 484938 37983 484941
rect 35758 484936 37983 484938
rect 35758 484880 37922 484936
rect 37978 484880 37983 484936
rect 35758 484878 37983 484880
rect 35758 484636 35818 484878
rect 37917 484875 37983 484878
rect 91093 484666 91159 484669
rect 118693 484666 118759 484669
rect 172513 484666 172579 484669
rect 89884 484664 91159 484666
rect 89884 484608 91098 484664
rect 91154 484608 91159 484664
rect 89884 484606 91159 484608
rect 116932 484664 118759 484666
rect 116932 484608 118698 484664
rect 118754 484608 118759 484664
rect 116932 484606 118759 484608
rect 170844 484664 172579 484666
rect 170844 484608 172518 484664
rect 172574 484608 172579 484664
rect 170844 484606 172579 484608
rect 91093 484603 91159 484606
rect 118693 484603 118759 484606
rect 172513 484603 172579 484606
rect 176561 484666 176627 484669
rect 178174 484666 178234 485180
rect 251774 485152 253938 485208
rect 253994 485152 253999 485208
rect 251774 485150 253999 485152
rect 200113 484666 200179 484669
rect 176561 484664 178234 484666
rect 176561 484608 176566 484664
rect 176622 484608 178234 484664
rect 176561 484606 178234 484608
rect 197892 484664 200179 484666
rect 197892 484608 200118 484664
rect 200174 484608 200179 484664
rect 251774 484636 251834 485150
rect 253933 485147 253999 485150
rect 256601 485210 256667 485213
rect 338021 485210 338087 485213
rect 361573 485210 361639 485213
rect 256601 485208 259164 485210
rect 256601 485152 256606 485208
rect 256662 485152 259164 485208
rect 256601 485150 259164 485152
rect 338021 485208 340124 485210
rect 338021 485152 338026 485208
rect 338082 485152 340124 485208
rect 338021 485150 340124 485152
rect 359782 485208 361639 485210
rect 359782 485152 361578 485208
rect 361634 485152 361639 485208
rect 359782 485150 361639 485152
rect 256601 485147 256667 485150
rect 338021 485147 338087 485150
rect 280153 484666 280219 484669
rect 335353 484666 335419 484669
rect 278852 484664 280219 484666
rect 197892 484606 200179 484608
rect 278852 484608 280158 484664
rect 280214 484608 280219 484664
rect 278852 484606 280219 484608
rect 332948 484664 335419 484666
rect 332948 484608 335358 484664
rect 335414 484608 335419 484664
rect 359782 484636 359842 485150
rect 361573 485147 361639 485150
rect 391841 485210 391907 485213
rect 445661 485210 445727 485213
rect 469213 485210 469279 485213
rect 391841 485208 394036 485210
rect 391841 485152 391846 485208
rect 391902 485152 394036 485208
rect 391841 485150 394036 485152
rect 445661 485208 448132 485210
rect 445661 485152 445666 485208
rect 445722 485152 448132 485208
rect 445661 485150 448132 485152
rect 467790 485208 469279 485210
rect 467790 485152 469218 485208
rect 469274 485152 469279 485208
rect 467790 485150 469279 485152
rect 391841 485147 391907 485150
rect 445661 485147 445727 485150
rect 415393 484666 415459 484669
rect 413908 484664 415459 484666
rect 332948 484606 335419 484608
rect 413908 484608 415398 484664
rect 415454 484608 415459 484664
rect 467790 484636 467850 485150
rect 469213 485147 469279 485150
rect 523033 484666 523099 484669
rect 550633 484666 550699 484669
rect 521916 484664 523099 484666
rect 413908 484606 415459 484608
rect 521916 484608 523038 484664
rect 523094 484608 523099 484664
rect 521916 484606 523099 484608
rect 548964 484664 550699 484666
rect 548964 484608 550638 484664
rect 550694 484608 550699 484664
rect 548964 484606 550699 484608
rect 176561 484603 176627 484606
rect 200113 484603 200179 484606
rect 280153 484603 280219 484606
rect 335353 484603 335419 484606
rect 415393 484603 415459 484606
rect 523033 484603 523099 484606
rect 550633 484603 550699 484606
rect 64873 484530 64939 484533
rect 146293 484530 146359 484533
rect 226333 484530 226399 484533
rect 307753 484530 307819 484533
rect 389173 484530 389239 484533
rect 442993 484530 443059 484533
rect 496813 484530 496879 484533
rect 62836 484528 64939 484530
rect 62836 484472 64878 484528
rect 64934 484472 64939 484528
rect 143950 484528 146359 484530
rect 62836 484470 64939 484472
rect 64873 484467 64939 484470
rect 143766 484394 143826 484500
rect 143950 484472 146298 484528
rect 146354 484472 146359 484528
rect 143950 484470 146359 484472
rect 224940 484528 226399 484530
rect 224940 484472 226338 484528
rect 226394 484472 226399 484528
rect 224940 484470 226399 484472
rect 305900 484528 307819 484530
rect 305900 484472 307758 484528
rect 307814 484472 307819 484528
rect 305900 484470 307819 484472
rect 386860 484528 389239 484530
rect 386860 484472 389178 484528
rect 389234 484472 389239 484528
rect 386860 484470 389239 484472
rect 440956 484528 443059 484530
rect 440956 484472 442998 484528
rect 443054 484472 443059 484528
rect 440956 484470 443059 484472
rect 494868 484528 496879 484530
rect 494868 484472 496818 484528
rect 496874 484472 496879 484528
rect 583520 484516 584960 484756
rect 494868 484470 496879 484472
rect 143950 484394 144010 484470
rect 146293 484467 146359 484470
rect 226333 484467 226399 484470
rect 307753 484467 307819 484470
rect 389173 484467 389239 484470
rect 442993 484467 443059 484470
rect 496813 484467 496879 484470
rect 143766 484334 144010 484394
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 68921 458962 68987 458965
rect 176561 458962 176627 458965
rect 284201 458962 284267 458965
rect 391841 458962 391907 458965
rect 473261 458962 473327 458965
rect 500861 458962 500927 458965
rect 68921 458960 70226 458962
rect 68921 458904 68926 458960
rect 68982 458904 70226 458960
rect 68921 458902 70226 458904
rect 68921 458899 68987 458902
rect 13721 458418 13787 458421
rect 41321 458418 41387 458421
rect 13721 458416 16100 458418
rect 13721 458360 13726 458416
rect 13782 458360 16100 458416
rect 13721 458358 16100 458360
rect 41321 458416 43148 458418
rect 41321 458360 41326 458416
rect 41382 458360 43148 458416
rect 70166 458388 70226 458902
rect 176561 458960 178234 458962
rect 176561 458904 176566 458960
rect 176622 458904 178234 458960
rect 176561 458902 178234 458904
rect 176561 458899 176627 458902
rect 95141 458418 95207 458421
rect 122741 458418 122807 458421
rect 148961 458418 149027 458421
rect 95141 458416 97060 458418
rect 41321 458358 43148 458360
rect 95141 458360 95146 458416
rect 95202 458360 97060 458416
rect 95141 458358 97060 458360
rect 122741 458416 124108 458418
rect 122741 458360 122746 458416
rect 122802 458360 124108 458416
rect 122741 458358 124108 458360
rect 148961 458416 151156 458418
rect 148961 458360 148966 458416
rect 149022 458360 151156 458416
rect 178174 458388 178234 458902
rect 284201 458960 286242 458962
rect 284201 458904 284206 458960
rect 284262 458904 286242 458960
rect 284201 458902 286242 458904
rect 284201 458899 284267 458902
rect 202781 458418 202847 458421
rect 230381 458418 230447 458421
rect 256601 458418 256667 458421
rect 202781 458416 205068 458418
rect 148961 458358 151156 458360
rect 202781 458360 202786 458416
rect 202842 458360 205068 458416
rect 202781 458358 205068 458360
rect 230381 458416 232116 458418
rect 230381 458360 230386 458416
rect 230442 458360 232116 458416
rect 230381 458358 232116 458360
rect 256601 458416 259164 458418
rect 256601 458360 256606 458416
rect 256662 458360 259164 458416
rect 286182 458388 286242 458902
rect 391841 458960 394066 458962
rect 391841 458904 391846 458960
rect 391902 458904 394066 458960
rect 391841 458902 394066 458904
rect 391841 458899 391907 458902
rect 311801 458418 311867 458421
rect 338021 458418 338087 458421
rect 365621 458418 365687 458421
rect 311801 458416 313076 458418
rect 256601 458358 259164 458360
rect 311801 458360 311806 458416
rect 311862 458360 313076 458416
rect 311801 458358 313076 458360
rect 338021 458416 340124 458418
rect 338021 458360 338026 458416
rect 338082 458360 340124 458416
rect 338021 458358 340124 458360
rect 365621 458416 367172 458418
rect 365621 458360 365626 458416
rect 365682 458360 367172 458416
rect 394006 458388 394066 458902
rect 473261 458960 475210 458962
rect 473261 458904 473266 458960
rect 473322 458904 475210 458960
rect 473261 458902 475210 458904
rect 473261 458899 473327 458902
rect 419441 458418 419507 458421
rect 445661 458418 445727 458421
rect 419441 458416 421084 458418
rect 365621 458358 367172 458360
rect 419441 458360 419446 458416
rect 419502 458360 421084 458416
rect 419441 458358 421084 458360
rect 445661 458416 448132 458418
rect 445661 458360 445666 458416
rect 445722 458360 448132 458416
rect 475150 458388 475210 458902
rect 500861 458960 502074 458962
rect 500861 458904 500866 458960
rect 500922 458904 502074 458960
rect 500861 458902 502074 458904
rect 500861 458899 500927 458902
rect 502014 458388 502074 458902
rect 526437 458418 526503 458421
rect 526437 458416 529092 458418
rect 445661 458358 448132 458360
rect 526437 458360 526442 458416
rect 526498 458360 529092 458416
rect 526437 458358 529092 458360
rect 13721 458355 13787 458358
rect 41321 458355 41387 458358
rect 95141 458355 95207 458358
rect 122741 458355 122807 458358
rect 148961 458355 149027 458358
rect 202781 458355 202847 458358
rect 230381 458355 230447 458358
rect 256601 458355 256667 458358
rect 311801 458355 311867 458358
rect 338021 458355 338087 458358
rect 365621 458355 365687 458358
rect 419441 458355 419507 458358
rect 445661 458355 445727 458358
rect 526437 458355 526503 458358
rect 146293 458146 146359 458149
rect 253933 458146 253999 458149
rect 361573 458146 361639 458149
rect 442993 458146 443059 458149
rect 469213 458146 469279 458149
rect 550633 458146 550699 458149
rect 143766 458144 146359 458146
rect 143766 458088 146298 458144
rect 146354 458088 146359 458144
rect 143766 458086 146359 458088
rect 64873 457738 64939 457741
rect 91093 457738 91159 457741
rect 118693 457738 118759 457741
rect 62836 457736 64939 457738
rect 62836 457680 64878 457736
rect 64934 457680 64939 457736
rect 62836 457678 64939 457680
rect 89884 457736 91159 457738
rect 89884 457680 91098 457736
rect 91154 457680 91159 457736
rect 89884 457678 91159 457680
rect 116932 457736 118759 457738
rect 116932 457680 118698 457736
rect 118754 457680 118759 457736
rect 143766 457708 143826 458086
rect 146293 458083 146359 458086
rect 251774 458144 253999 458146
rect 251774 458088 253938 458144
rect 253994 458088 253999 458144
rect 251774 458086 253999 458088
rect 172513 457738 172579 457741
rect 200113 457738 200179 457741
rect 226333 457738 226399 457741
rect 170844 457736 172579 457738
rect 116932 457678 118759 457680
rect 170844 457680 172518 457736
rect 172574 457680 172579 457736
rect 170844 457678 172579 457680
rect 197892 457736 200179 457738
rect 197892 457680 200118 457736
rect 200174 457680 200179 457736
rect 197892 457678 200179 457680
rect 224940 457736 226399 457738
rect 224940 457680 226338 457736
rect 226394 457680 226399 457736
rect 251774 457708 251834 458086
rect 253933 458083 253999 458086
rect 359782 458144 361639 458146
rect 359782 458088 361578 458144
rect 361634 458088 361639 458144
rect 359782 458086 361639 458088
rect 280153 457738 280219 457741
rect 307753 457738 307819 457741
rect 335353 457738 335419 457741
rect 278852 457736 280219 457738
rect 224940 457678 226399 457680
rect 278852 457680 280158 457736
rect 280214 457680 280219 457736
rect 278852 457678 280219 457680
rect 305900 457736 307819 457738
rect 305900 457680 307758 457736
rect 307814 457680 307819 457736
rect 305900 457678 307819 457680
rect 332948 457736 335419 457738
rect 332948 457680 335358 457736
rect 335414 457680 335419 457736
rect 359782 457708 359842 458086
rect 361573 458083 361639 458086
rect 440926 458144 443059 458146
rect 440926 458088 442998 458144
rect 443054 458088 443059 458144
rect 440926 458086 443059 458088
rect 389173 457738 389239 457741
rect 415393 457738 415459 457741
rect 386860 457736 389239 457738
rect 332948 457678 335419 457680
rect 386860 457680 389178 457736
rect 389234 457680 389239 457736
rect 386860 457678 389239 457680
rect 413908 457736 415459 457738
rect 413908 457680 415398 457736
rect 415454 457680 415459 457736
rect 440926 457708 440986 458086
rect 442993 458083 443059 458086
rect 467790 458144 469279 458146
rect 467790 458088 469218 458144
rect 469274 458088 469279 458144
rect 467790 458086 469279 458088
rect 467790 457708 467850 458086
rect 469213 458083 469279 458086
rect 548934 458144 550699 458146
rect 548934 458088 550638 458144
rect 550694 458088 550699 458144
rect 548934 458086 550699 458088
rect 496813 457738 496879 457741
rect 523033 457738 523099 457741
rect 494868 457736 496879 457738
rect 413908 457678 415459 457680
rect 494868 457680 496818 457736
rect 496874 457680 496879 457736
rect 494868 457678 496879 457680
rect 521916 457736 523099 457738
rect 521916 457680 523038 457736
rect 523094 457680 523099 457736
rect 548934 457708 548994 458086
rect 550633 458083 550699 458086
rect 580349 458146 580415 458149
rect 583520 458146 584960 458236
rect 580349 458144 584960 458146
rect 580349 458088 580354 458144
rect 580410 458088 584960 458144
rect 580349 458086 584960 458088
rect 580349 458083 580415 458086
rect 583520 457996 584960 458086
rect 521916 457678 523099 457680
rect 64873 457675 64939 457678
rect 91093 457675 91159 457678
rect 118693 457675 118759 457678
rect 172513 457675 172579 457678
rect 200113 457675 200179 457678
rect 226333 457675 226399 457678
rect 280153 457675 280219 457678
rect 307753 457675 307819 457678
rect 335353 457675 335419 457678
rect 389173 457675 389239 457678
rect 415393 457675 415459 457678
rect 496813 457675 496879 457678
rect 523033 457675 523099 457678
rect 35758 457058 35818 457572
rect 37917 457058 37983 457061
rect 35758 457056 37983 457058
rect 35758 457000 37922 457056
rect 37978 457000 37983 457056
rect 35758 456998 37983 457000
rect 37917 456995 37983 456998
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 68921 431626 68987 431629
rect 176561 431626 176627 431629
rect 284201 431626 284267 431629
rect 473261 431626 473327 431629
rect 68921 431624 70226 431626
rect 68921 431568 68926 431624
rect 68982 431568 70226 431624
rect 68921 431566 70226 431568
rect 68921 431563 68987 431566
rect 13721 431354 13787 431357
rect 41321 431354 41387 431357
rect 13721 431352 16100 431354
rect 13721 431296 13726 431352
rect 13782 431296 16100 431352
rect 13721 431294 16100 431296
rect 41321 431352 43148 431354
rect 41321 431296 41326 431352
rect 41382 431296 43148 431352
rect 70166 431324 70226 431566
rect 176561 431624 178234 431626
rect 176561 431568 176566 431624
rect 176622 431568 178234 431624
rect 176561 431566 178234 431568
rect 176561 431563 176627 431566
rect 95141 431354 95207 431357
rect 122741 431354 122807 431357
rect 148961 431354 149027 431357
rect 95141 431352 97060 431354
rect 41321 431294 43148 431296
rect 95141 431296 95146 431352
rect 95202 431296 97060 431352
rect 95141 431294 97060 431296
rect 122741 431352 124108 431354
rect 122741 431296 122746 431352
rect 122802 431296 124108 431352
rect 122741 431294 124108 431296
rect 148961 431352 151156 431354
rect 148961 431296 148966 431352
rect 149022 431296 151156 431352
rect 178174 431324 178234 431566
rect 284201 431624 286242 431626
rect 284201 431568 284206 431624
rect 284262 431568 286242 431624
rect 284201 431566 286242 431568
rect 284201 431563 284267 431566
rect 202781 431354 202847 431357
rect 230381 431354 230447 431357
rect 256601 431354 256667 431357
rect 202781 431352 205068 431354
rect 148961 431294 151156 431296
rect 202781 431296 202786 431352
rect 202842 431296 205068 431352
rect 202781 431294 205068 431296
rect 230381 431352 232116 431354
rect 230381 431296 230386 431352
rect 230442 431296 232116 431352
rect 230381 431294 232116 431296
rect 256601 431352 259164 431354
rect 256601 431296 256606 431352
rect 256662 431296 259164 431352
rect 286182 431324 286242 431566
rect 473261 431624 475210 431626
rect 473261 431568 473266 431624
rect 473322 431568 475210 431624
rect 473261 431566 475210 431568
rect 473261 431563 473327 431566
rect 311801 431354 311867 431357
rect 338021 431354 338087 431357
rect 365621 431354 365687 431357
rect 391841 431354 391907 431357
rect 419441 431354 419507 431357
rect 445661 431354 445727 431357
rect 311801 431352 313076 431354
rect 256601 431294 259164 431296
rect 311801 431296 311806 431352
rect 311862 431296 313076 431352
rect 311801 431294 313076 431296
rect 338021 431352 340124 431354
rect 338021 431296 338026 431352
rect 338082 431296 340124 431352
rect 338021 431294 340124 431296
rect 365621 431352 367172 431354
rect 365621 431296 365626 431352
rect 365682 431296 367172 431352
rect 365621 431294 367172 431296
rect 391841 431352 394036 431354
rect 391841 431296 391846 431352
rect 391902 431296 394036 431352
rect 391841 431294 394036 431296
rect 419441 431352 421084 431354
rect 419441 431296 419446 431352
rect 419502 431296 421084 431352
rect 419441 431294 421084 431296
rect 445661 431352 448132 431354
rect 445661 431296 445666 431352
rect 445722 431296 448132 431352
rect 475150 431324 475210 431566
rect 583520 431476 584960 431716
rect 500861 431354 500927 431357
rect 526437 431354 526503 431357
rect 500861 431352 502044 431354
rect 445661 431294 448132 431296
rect 500861 431296 500866 431352
rect 500922 431296 502044 431352
rect 500861 431294 502044 431296
rect 526437 431352 529092 431354
rect 526437 431296 526442 431352
rect 526498 431296 529092 431352
rect 526437 431294 529092 431296
rect 13721 431291 13787 431294
rect 41321 431291 41387 431294
rect 95141 431291 95207 431294
rect 122741 431291 122807 431294
rect 148961 431291 149027 431294
rect 202781 431291 202847 431294
rect 230381 431291 230447 431294
rect 256601 431291 256667 431294
rect 311801 431291 311867 431294
rect 338021 431291 338087 431294
rect 365621 431291 365687 431294
rect 391841 431291 391907 431294
rect 419441 431291 419507 431294
rect 445661 431291 445727 431294
rect 500861 431291 500927 431294
rect 526437 431291 526503 431294
rect 146293 431218 146359 431221
rect 253933 431218 253999 431221
rect 361573 431218 361639 431221
rect 469213 431218 469279 431221
rect 143766 431216 146359 431218
rect 143766 431160 146298 431216
rect 146354 431160 146359 431216
rect 143766 431158 146359 431160
rect 37917 430946 37983 430949
rect 35758 430944 37983 430946
rect 35758 430888 37922 430944
rect 37978 430888 37983 430944
rect 35758 430886 37983 430888
rect 35758 430644 35818 430886
rect 37917 430883 37983 430886
rect 64873 430674 64939 430677
rect 91093 430674 91159 430677
rect 118693 430674 118759 430677
rect 62836 430672 64939 430674
rect 62836 430616 64878 430672
rect 64934 430616 64939 430672
rect 62836 430614 64939 430616
rect 89884 430672 91159 430674
rect 89884 430616 91098 430672
rect 91154 430616 91159 430672
rect 89884 430614 91159 430616
rect 116932 430672 118759 430674
rect 116932 430616 118698 430672
rect 118754 430616 118759 430672
rect 143766 430644 143826 431158
rect 146293 431155 146359 431158
rect 251774 431216 253999 431218
rect 251774 431160 253938 431216
rect 253994 431160 253999 431216
rect 251774 431158 253999 431160
rect 172513 430674 172579 430677
rect 200113 430674 200179 430677
rect 226333 430674 226399 430677
rect 170844 430672 172579 430674
rect 116932 430614 118759 430616
rect 170844 430616 172518 430672
rect 172574 430616 172579 430672
rect 170844 430614 172579 430616
rect 197892 430672 200179 430674
rect 197892 430616 200118 430672
rect 200174 430616 200179 430672
rect 197892 430614 200179 430616
rect 224940 430672 226399 430674
rect 224940 430616 226338 430672
rect 226394 430616 226399 430672
rect 251774 430644 251834 431158
rect 253933 431155 253999 431158
rect 359782 431216 361639 431218
rect 359782 431160 361578 431216
rect 361634 431160 361639 431216
rect 359782 431158 361639 431160
rect 280153 430674 280219 430677
rect 307753 430674 307819 430677
rect 335353 430674 335419 430677
rect 278852 430672 280219 430674
rect 224940 430614 226399 430616
rect 278852 430616 280158 430672
rect 280214 430616 280219 430672
rect 278852 430614 280219 430616
rect 305900 430672 307819 430674
rect 305900 430616 307758 430672
rect 307814 430616 307819 430672
rect 305900 430614 307819 430616
rect 332948 430672 335419 430674
rect 332948 430616 335358 430672
rect 335414 430616 335419 430672
rect 359782 430644 359842 431158
rect 361573 431155 361639 431158
rect 467790 431216 469279 431218
rect 467790 431160 469218 431216
rect 469274 431160 469279 431216
rect 467790 431158 469279 431160
rect 389173 430674 389239 430677
rect 415393 430674 415459 430677
rect 442993 430674 443059 430677
rect 386860 430672 389239 430674
rect 332948 430614 335419 430616
rect 386860 430616 389178 430672
rect 389234 430616 389239 430672
rect 386860 430614 389239 430616
rect 413908 430672 415459 430674
rect 413908 430616 415398 430672
rect 415454 430616 415459 430672
rect 413908 430614 415459 430616
rect 440956 430672 443059 430674
rect 440956 430616 442998 430672
rect 443054 430616 443059 430672
rect 467790 430644 467850 431158
rect 469213 431155 469279 431158
rect 496813 430674 496879 430677
rect 523033 430674 523099 430677
rect 550633 430674 550699 430677
rect 494868 430672 496879 430674
rect 440956 430614 443059 430616
rect 494868 430616 496818 430672
rect 496874 430616 496879 430672
rect 494868 430614 496879 430616
rect 521916 430672 523099 430674
rect 521916 430616 523038 430672
rect 523094 430616 523099 430672
rect 521916 430614 523099 430616
rect 548964 430672 550699 430674
rect 548964 430616 550638 430672
rect 550694 430616 550699 430672
rect 548964 430614 550699 430616
rect 64873 430611 64939 430614
rect 91093 430611 91159 430614
rect 118693 430611 118759 430614
rect 172513 430611 172579 430614
rect 200113 430611 200179 430614
rect 226333 430611 226399 430614
rect 280153 430611 280219 430614
rect 307753 430611 307819 430614
rect 335353 430611 335419 430614
rect 389173 430611 389239 430614
rect 415393 430611 415459 430614
rect 442993 430611 443059 430614
rect 496813 430611 496879 430614
rect 523033 430611 523099 430614
rect 550633 430611 550699 430614
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 580441 404970 580507 404973
rect 583520 404970 584960 405060
rect 580441 404968 584960 404970
rect 580441 404912 580446 404968
rect 580502 404912 584960 404968
rect 580441 404910 584960 404912
rect 580441 404907 580507 404910
rect 583520 404820 584960 404910
rect 13721 404290 13787 404293
rect 41321 404290 41387 404293
rect 95141 404290 95207 404293
rect 122741 404290 122807 404293
rect 148961 404290 149027 404293
rect 202781 404290 202847 404293
rect 230381 404290 230447 404293
rect 256601 404290 256667 404293
rect 311801 404290 311867 404293
rect 338021 404290 338087 404293
rect 365621 404290 365687 404293
rect 391841 404290 391907 404293
rect 419441 404290 419507 404293
rect 445661 404290 445727 404293
rect 500861 404290 500927 404293
rect 526437 404290 526503 404293
rect 13721 404288 16100 404290
rect 13721 404232 13726 404288
rect 13782 404232 16100 404288
rect 13721 404230 16100 404232
rect 41321 404288 43148 404290
rect 41321 404232 41326 404288
rect 41382 404232 43148 404288
rect 95141 404288 97060 404290
rect 41321 404230 43148 404232
rect 13721 404227 13787 404230
rect 41321 404227 41387 404230
rect 68921 403746 68987 403749
rect 70166 403746 70226 404260
rect 95141 404232 95146 404288
rect 95202 404232 97060 404288
rect 95141 404230 97060 404232
rect 122741 404288 124108 404290
rect 122741 404232 122746 404288
rect 122802 404232 124108 404288
rect 122741 404230 124108 404232
rect 148961 404288 151156 404290
rect 148961 404232 148966 404288
rect 149022 404232 151156 404288
rect 202781 404288 205068 404290
rect 148961 404230 151156 404232
rect 95141 404227 95207 404230
rect 122741 404227 122807 404230
rect 148961 404227 149027 404230
rect 68921 403744 70226 403746
rect 68921 403688 68926 403744
rect 68982 403688 70226 403744
rect 68921 403686 70226 403688
rect 176561 403746 176627 403749
rect 178174 403746 178234 404260
rect 202781 404232 202786 404288
rect 202842 404232 205068 404288
rect 202781 404230 205068 404232
rect 230381 404288 232116 404290
rect 230381 404232 230386 404288
rect 230442 404232 232116 404288
rect 230381 404230 232116 404232
rect 256601 404288 259164 404290
rect 256601 404232 256606 404288
rect 256662 404232 259164 404288
rect 311801 404288 313076 404290
rect 256601 404230 259164 404232
rect 202781 404227 202847 404230
rect 230381 404227 230447 404230
rect 256601 404227 256667 404230
rect 176561 403744 178234 403746
rect 176561 403688 176566 403744
rect 176622 403688 178234 403744
rect 176561 403686 178234 403688
rect 284201 403746 284267 403749
rect 286182 403746 286242 404260
rect 311801 404232 311806 404288
rect 311862 404232 313076 404288
rect 311801 404230 313076 404232
rect 338021 404288 340124 404290
rect 338021 404232 338026 404288
rect 338082 404232 340124 404288
rect 338021 404230 340124 404232
rect 365621 404288 367172 404290
rect 365621 404232 365626 404288
rect 365682 404232 367172 404288
rect 365621 404230 367172 404232
rect 391841 404288 394036 404290
rect 391841 404232 391846 404288
rect 391902 404232 394036 404288
rect 391841 404230 394036 404232
rect 419441 404288 421084 404290
rect 419441 404232 419446 404288
rect 419502 404232 421084 404288
rect 419441 404230 421084 404232
rect 445661 404288 448132 404290
rect 445661 404232 445666 404288
rect 445722 404232 448132 404288
rect 500861 404288 502044 404290
rect 445661 404230 448132 404232
rect 311801 404227 311867 404230
rect 338021 404227 338087 404230
rect 365621 404227 365687 404230
rect 391841 404227 391907 404230
rect 419441 404227 419507 404230
rect 445661 404227 445727 404230
rect 284201 403744 286242 403746
rect 284201 403688 284206 403744
rect 284262 403688 286242 403744
rect 284201 403686 286242 403688
rect 473261 403746 473327 403749
rect 475150 403746 475210 404260
rect 500861 404232 500866 404288
rect 500922 404232 502044 404288
rect 500861 404230 502044 404232
rect 526437 404288 529092 404290
rect 526437 404232 526442 404288
rect 526498 404232 529092 404288
rect 526437 404230 529092 404232
rect 500861 404227 500927 404230
rect 526437 404227 526503 404230
rect 473261 403744 475210 403746
rect 473261 403688 473266 403744
rect 473322 403688 475210 403744
rect 473261 403686 475210 403688
rect 68921 403683 68987 403686
rect 176561 403683 176627 403686
rect 284201 403683 284267 403686
rect 473261 403683 473327 403686
rect 64873 403610 64939 403613
rect 91093 403610 91159 403613
rect 118693 403610 118759 403613
rect 172513 403610 172579 403613
rect 200113 403610 200179 403613
rect 226333 403610 226399 403613
rect 280153 403610 280219 403613
rect 307753 403610 307819 403613
rect 335353 403610 335419 403613
rect 389173 403610 389239 403613
rect 415393 403610 415459 403613
rect 442993 403610 443059 403613
rect 496813 403610 496879 403613
rect 523033 403610 523099 403613
rect 550633 403610 550699 403613
rect 62836 403608 64939 403610
rect 35758 403066 35818 403580
rect 62836 403552 64878 403608
rect 64934 403552 64939 403608
rect 62836 403550 64939 403552
rect 89884 403608 91159 403610
rect 89884 403552 91098 403608
rect 91154 403552 91159 403608
rect 89884 403550 91159 403552
rect 116932 403608 118759 403610
rect 116932 403552 118698 403608
rect 118754 403552 118759 403608
rect 170844 403608 172579 403610
rect 116932 403550 118759 403552
rect 64873 403547 64939 403550
rect 91093 403547 91159 403550
rect 118693 403547 118759 403550
rect 143766 403338 143826 403580
rect 170844 403552 172518 403608
rect 172574 403552 172579 403608
rect 170844 403550 172579 403552
rect 197892 403608 200179 403610
rect 197892 403552 200118 403608
rect 200174 403552 200179 403608
rect 197892 403550 200179 403552
rect 224940 403608 226399 403610
rect 224940 403552 226338 403608
rect 226394 403552 226399 403608
rect 278852 403608 280219 403610
rect 224940 403550 226399 403552
rect 172513 403547 172579 403550
rect 200113 403547 200179 403550
rect 226333 403547 226399 403550
rect 146293 403338 146359 403341
rect 143766 403336 146359 403338
rect 143766 403280 146298 403336
rect 146354 403280 146359 403336
rect 143766 403278 146359 403280
rect 251774 403338 251834 403580
rect 278852 403552 280158 403608
rect 280214 403552 280219 403608
rect 278852 403550 280219 403552
rect 305900 403608 307819 403610
rect 305900 403552 307758 403608
rect 307814 403552 307819 403608
rect 305900 403550 307819 403552
rect 332948 403608 335419 403610
rect 332948 403552 335358 403608
rect 335414 403552 335419 403608
rect 386860 403608 389239 403610
rect 332948 403550 335419 403552
rect 280153 403547 280219 403550
rect 307753 403547 307819 403550
rect 335353 403547 335419 403550
rect 253933 403338 253999 403341
rect 251774 403336 253999 403338
rect 251774 403280 253938 403336
rect 253994 403280 253999 403336
rect 251774 403278 253999 403280
rect 359782 403338 359842 403580
rect 386860 403552 389178 403608
rect 389234 403552 389239 403608
rect 386860 403550 389239 403552
rect 413908 403608 415459 403610
rect 413908 403552 415398 403608
rect 415454 403552 415459 403608
rect 413908 403550 415459 403552
rect 440956 403608 443059 403610
rect 440956 403552 442998 403608
rect 443054 403552 443059 403608
rect 494868 403608 496879 403610
rect 440956 403550 443059 403552
rect 389173 403547 389239 403550
rect 415393 403547 415459 403550
rect 442993 403547 443059 403550
rect 361573 403338 361639 403341
rect 359782 403336 361639 403338
rect 359782 403280 361578 403336
rect 361634 403280 361639 403336
rect 359782 403278 361639 403280
rect 467790 403338 467850 403580
rect 494868 403552 496818 403608
rect 496874 403552 496879 403608
rect 494868 403550 496879 403552
rect 521916 403608 523099 403610
rect 521916 403552 523038 403608
rect 523094 403552 523099 403608
rect 521916 403550 523099 403552
rect 548964 403608 550699 403610
rect 548964 403552 550638 403608
rect 550694 403552 550699 403608
rect 548964 403550 550699 403552
rect 496813 403547 496879 403550
rect 523033 403547 523099 403550
rect 550633 403547 550699 403550
rect 469213 403338 469279 403341
rect 467790 403336 469279 403338
rect 467790 403280 469218 403336
rect 469274 403280 469279 403336
rect 467790 403278 469279 403280
rect 146293 403275 146359 403278
rect 253933 403275 253999 403278
rect 361573 403275 361639 403278
rect 469213 403275 469279 403278
rect 37917 403066 37983 403069
rect 35758 403064 37983 403066
rect 35758 403008 37922 403064
rect 37978 403008 37983 403064
rect 35758 403006 37983 403008
rect 37917 403003 37983 403006
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect 526437 377362 526503 377365
rect 526437 377360 529092 377362
rect 526437 377304 526442 377360
rect 526498 377304 529092 377360
rect 526437 377302 529092 377304
rect 526437 377299 526503 377302
rect 13721 377226 13787 377229
rect 41321 377226 41387 377229
rect 95141 377226 95207 377229
rect 122741 377226 122807 377229
rect 148961 377226 149027 377229
rect 202781 377226 202847 377229
rect 230381 377226 230447 377229
rect 256601 377226 256667 377229
rect 311801 377226 311867 377229
rect 338021 377226 338087 377229
rect 365621 377226 365687 377229
rect 391841 377226 391907 377229
rect 419441 377226 419507 377229
rect 445661 377226 445727 377229
rect 500861 377226 500927 377229
rect 13721 377224 16100 377226
rect 13721 377168 13726 377224
rect 13782 377168 16100 377224
rect 13721 377166 16100 377168
rect 41321 377224 43148 377226
rect 41321 377168 41326 377224
rect 41382 377168 43148 377224
rect 95141 377224 97060 377226
rect 41321 377166 43148 377168
rect 13721 377163 13787 377166
rect 41321 377163 41387 377166
rect 68921 376818 68987 376821
rect 70166 376818 70226 377196
rect 95141 377168 95146 377224
rect 95202 377168 97060 377224
rect 95141 377166 97060 377168
rect 122741 377224 124108 377226
rect 122741 377168 122746 377224
rect 122802 377168 124108 377224
rect 122741 377166 124108 377168
rect 148961 377224 151156 377226
rect 148961 377168 148966 377224
rect 149022 377168 151156 377224
rect 202781 377224 205068 377226
rect 148961 377166 151156 377168
rect 95141 377163 95207 377166
rect 122741 377163 122807 377166
rect 148961 377163 149027 377166
rect 68921 376816 70226 376818
rect 68921 376760 68926 376816
rect 68982 376760 70226 376816
rect 68921 376758 70226 376760
rect 176561 376818 176627 376821
rect 178174 376818 178234 377196
rect 202781 377168 202786 377224
rect 202842 377168 205068 377224
rect 202781 377166 205068 377168
rect 230381 377224 232116 377226
rect 230381 377168 230386 377224
rect 230442 377168 232116 377224
rect 230381 377166 232116 377168
rect 256601 377224 259164 377226
rect 256601 377168 256606 377224
rect 256662 377168 259164 377224
rect 311801 377224 313076 377226
rect 256601 377166 259164 377168
rect 202781 377163 202847 377166
rect 230381 377163 230447 377166
rect 256601 377163 256667 377166
rect 176561 376816 178234 376818
rect 176561 376760 176566 376816
rect 176622 376760 178234 376816
rect 176561 376758 178234 376760
rect 284201 376818 284267 376821
rect 286182 376818 286242 377196
rect 311801 377168 311806 377224
rect 311862 377168 313076 377224
rect 311801 377166 313076 377168
rect 338021 377224 340124 377226
rect 338021 377168 338026 377224
rect 338082 377168 340124 377224
rect 338021 377166 340124 377168
rect 365621 377224 367172 377226
rect 365621 377168 365626 377224
rect 365682 377168 367172 377224
rect 365621 377166 367172 377168
rect 391841 377224 394036 377226
rect 391841 377168 391846 377224
rect 391902 377168 394036 377224
rect 391841 377166 394036 377168
rect 419441 377224 421084 377226
rect 419441 377168 419446 377224
rect 419502 377168 421084 377224
rect 419441 377166 421084 377168
rect 445661 377224 448132 377226
rect 445661 377168 445666 377224
rect 445722 377168 448132 377224
rect 500861 377224 502044 377226
rect 445661 377166 448132 377168
rect 311801 377163 311867 377166
rect 338021 377163 338087 377166
rect 365621 377163 365687 377166
rect 391841 377163 391907 377166
rect 419441 377163 419507 377166
rect 445661 377163 445727 377166
rect 284201 376816 286242 376818
rect 284201 376760 284206 376816
rect 284262 376760 286242 376816
rect 284201 376758 286242 376760
rect 473261 376818 473327 376821
rect 475150 376818 475210 377196
rect 500861 377168 500866 377224
rect 500922 377168 502044 377224
rect 500861 377166 502044 377168
rect 500861 377163 500927 377166
rect 473261 376816 475210 376818
rect 473261 376760 473266 376816
rect 473322 376760 475210 376816
rect 473261 376758 475210 376760
rect 68921 376755 68987 376758
rect 176561 376755 176627 376758
rect 284201 376755 284267 376758
rect 473261 376755 473327 376758
rect 64873 376546 64939 376549
rect 91093 376546 91159 376549
rect 118693 376546 118759 376549
rect 172513 376546 172579 376549
rect 200113 376546 200179 376549
rect 226333 376546 226399 376549
rect 280153 376546 280219 376549
rect 307753 376546 307819 376549
rect 335353 376546 335419 376549
rect 389173 376546 389239 376549
rect 415393 376546 415459 376549
rect 442993 376546 443059 376549
rect 496813 376546 496879 376549
rect 523033 376546 523099 376549
rect 550633 376546 550699 376549
rect 62836 376544 64939 376546
rect 35758 376002 35818 376516
rect 62836 376488 64878 376544
rect 64934 376488 64939 376544
rect 62836 376486 64939 376488
rect 89884 376544 91159 376546
rect 89884 376488 91098 376544
rect 91154 376488 91159 376544
rect 89884 376486 91159 376488
rect 116932 376544 118759 376546
rect 116932 376488 118698 376544
rect 118754 376488 118759 376544
rect 170844 376544 172579 376546
rect 116932 376486 118759 376488
rect 64873 376483 64939 376486
rect 91093 376483 91159 376486
rect 118693 376483 118759 376486
rect 37917 376002 37983 376005
rect 35758 376000 37983 376002
rect 35758 375944 37922 376000
rect 37978 375944 37983 376000
rect 35758 375942 37983 375944
rect 143766 376002 143826 376516
rect 170844 376488 172518 376544
rect 172574 376488 172579 376544
rect 170844 376486 172579 376488
rect 197892 376544 200179 376546
rect 197892 376488 200118 376544
rect 200174 376488 200179 376544
rect 197892 376486 200179 376488
rect 224940 376544 226399 376546
rect 224940 376488 226338 376544
rect 226394 376488 226399 376544
rect 278852 376544 280219 376546
rect 224940 376486 226399 376488
rect 172513 376483 172579 376486
rect 200113 376483 200179 376486
rect 226333 376483 226399 376486
rect 144821 376002 144887 376005
rect 143766 376000 144887 376002
rect 143766 375944 144826 376000
rect 144882 375944 144887 376000
rect 143766 375942 144887 375944
rect 251774 376002 251834 376516
rect 278852 376488 280158 376544
rect 280214 376488 280219 376544
rect 278852 376486 280219 376488
rect 305900 376544 307819 376546
rect 305900 376488 307758 376544
rect 307814 376488 307819 376544
rect 305900 376486 307819 376488
rect 332948 376544 335419 376546
rect 332948 376488 335358 376544
rect 335414 376488 335419 376544
rect 386860 376544 389239 376546
rect 332948 376486 335419 376488
rect 280153 376483 280219 376486
rect 307753 376483 307819 376486
rect 335353 376483 335419 376486
rect 253933 376002 253999 376005
rect 251774 376000 253999 376002
rect 251774 375944 253938 376000
rect 253994 375944 253999 376000
rect 251774 375942 253999 375944
rect 359782 376002 359842 376516
rect 386860 376488 389178 376544
rect 389234 376488 389239 376544
rect 386860 376486 389239 376488
rect 413908 376544 415459 376546
rect 413908 376488 415398 376544
rect 415454 376488 415459 376544
rect 413908 376486 415459 376488
rect 440956 376544 443059 376546
rect 440956 376488 442998 376544
rect 443054 376488 443059 376544
rect 494868 376544 496879 376546
rect 440956 376486 443059 376488
rect 389173 376483 389239 376486
rect 415393 376483 415459 376486
rect 442993 376483 443059 376486
rect 361573 376002 361639 376005
rect 359782 376000 361639 376002
rect 359782 375944 361578 376000
rect 361634 375944 361639 376000
rect 359782 375942 361639 375944
rect 467790 376002 467850 376516
rect 494868 376488 496818 376544
rect 496874 376488 496879 376544
rect 494868 376486 496879 376488
rect 521916 376544 523099 376546
rect 521916 376488 523038 376544
rect 523094 376488 523099 376544
rect 521916 376486 523099 376488
rect 548964 376544 550699 376546
rect 548964 376488 550638 376544
rect 550694 376488 550699 376544
rect 548964 376486 550699 376488
rect 496813 376483 496879 376486
rect 523033 376483 523099 376486
rect 550633 376483 550699 376486
rect 469213 376002 469279 376005
rect 467790 376000 469279 376002
rect 467790 375944 469218 376000
rect 469274 375944 469279 376000
rect 467790 375942 469279 375944
rect 37917 375939 37983 375942
rect 144821 375939 144887 375942
rect 253933 375939 253999 375942
rect 361573 375939 361639 375942
rect 469213 375939 469279 375942
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 580533 351930 580599 351933
rect 583520 351930 584960 352020
rect 580533 351928 584960 351930
rect 580533 351872 580538 351928
rect 580594 351872 584960 351928
rect 580533 351870 584960 351872
rect 580533 351867 580599 351870
rect 583520 351780 584960 351870
rect 13721 350298 13787 350301
rect 41321 350298 41387 350301
rect 95141 350298 95207 350301
rect 122741 350298 122807 350301
rect 148961 350298 149027 350301
rect 202781 350298 202847 350301
rect 230381 350298 230447 350301
rect 256601 350298 256667 350301
rect 311801 350298 311867 350301
rect 338021 350298 338087 350301
rect 365621 350298 365687 350301
rect 391841 350298 391907 350301
rect 419441 350298 419507 350301
rect 445661 350298 445727 350301
rect 500861 350298 500927 350301
rect 526437 350298 526503 350301
rect 13721 350296 16100 350298
rect 13721 350240 13726 350296
rect 13782 350240 16100 350296
rect 13721 350238 16100 350240
rect 41321 350296 43148 350298
rect 41321 350240 41326 350296
rect 41382 350240 43148 350296
rect 95141 350296 97060 350298
rect 41321 350238 43148 350240
rect 13721 350235 13787 350238
rect 41321 350235 41387 350238
rect 68921 349754 68987 349757
rect 70166 349754 70226 350268
rect 95141 350240 95146 350296
rect 95202 350240 97060 350296
rect 95141 350238 97060 350240
rect 122741 350296 124108 350298
rect 122741 350240 122746 350296
rect 122802 350240 124108 350296
rect 122741 350238 124108 350240
rect 148961 350296 151156 350298
rect 148961 350240 148966 350296
rect 149022 350240 151156 350296
rect 202781 350296 205068 350298
rect 148961 350238 151156 350240
rect 95141 350235 95207 350238
rect 122741 350235 122807 350238
rect 148961 350235 149027 350238
rect 68921 349752 70226 349754
rect 68921 349696 68926 349752
rect 68982 349696 70226 349752
rect 68921 349694 70226 349696
rect 176561 349754 176627 349757
rect 178174 349754 178234 350268
rect 202781 350240 202786 350296
rect 202842 350240 205068 350296
rect 202781 350238 205068 350240
rect 230381 350296 232116 350298
rect 230381 350240 230386 350296
rect 230442 350240 232116 350296
rect 230381 350238 232116 350240
rect 256601 350296 259164 350298
rect 256601 350240 256606 350296
rect 256662 350240 259164 350296
rect 311801 350296 313076 350298
rect 256601 350238 259164 350240
rect 202781 350235 202847 350238
rect 230381 350235 230447 350238
rect 256601 350235 256667 350238
rect 176561 349752 178234 349754
rect 176561 349696 176566 349752
rect 176622 349696 178234 349752
rect 176561 349694 178234 349696
rect 284201 349754 284267 349757
rect 286182 349754 286242 350268
rect 311801 350240 311806 350296
rect 311862 350240 313076 350296
rect 311801 350238 313076 350240
rect 338021 350296 340124 350298
rect 338021 350240 338026 350296
rect 338082 350240 340124 350296
rect 338021 350238 340124 350240
rect 365621 350296 367172 350298
rect 365621 350240 365626 350296
rect 365682 350240 367172 350296
rect 365621 350238 367172 350240
rect 391841 350296 394036 350298
rect 391841 350240 391846 350296
rect 391902 350240 394036 350296
rect 391841 350238 394036 350240
rect 419441 350296 421084 350298
rect 419441 350240 419446 350296
rect 419502 350240 421084 350296
rect 419441 350238 421084 350240
rect 445661 350296 448132 350298
rect 445661 350240 445666 350296
rect 445722 350240 448132 350296
rect 500861 350296 502044 350298
rect 445661 350238 448132 350240
rect 311801 350235 311867 350238
rect 338021 350235 338087 350238
rect 365621 350235 365687 350238
rect 391841 350235 391907 350238
rect 419441 350235 419507 350238
rect 445661 350235 445727 350238
rect 284201 349752 286242 349754
rect 284201 349696 284206 349752
rect 284262 349696 286242 349752
rect 284201 349694 286242 349696
rect 473261 349754 473327 349757
rect 475150 349754 475210 350268
rect 500861 350240 500866 350296
rect 500922 350240 502044 350296
rect 500861 350238 502044 350240
rect 526437 350296 529092 350298
rect 526437 350240 526442 350296
rect 526498 350240 529092 350296
rect 526437 350238 529092 350240
rect 500861 350235 500927 350238
rect 526437 350235 526503 350238
rect 473261 349752 475210 349754
rect 473261 349696 473266 349752
rect 473322 349696 475210 349752
rect 473261 349694 475210 349696
rect 68921 349691 68987 349694
rect 176561 349691 176627 349694
rect 284201 349691 284267 349694
rect 473261 349691 473327 349694
rect 64873 349618 64939 349621
rect 91093 349618 91159 349621
rect 118693 349618 118759 349621
rect 172513 349618 172579 349621
rect 200113 349618 200179 349621
rect 226333 349618 226399 349621
rect 280153 349618 280219 349621
rect 307753 349618 307819 349621
rect 335353 349618 335419 349621
rect 389173 349618 389239 349621
rect 415393 349618 415459 349621
rect 442993 349618 443059 349621
rect 496813 349618 496879 349621
rect 523033 349618 523099 349621
rect 550633 349618 550699 349621
rect 62836 349616 64939 349618
rect 35758 349210 35818 349588
rect 62836 349560 64878 349616
rect 64934 349560 64939 349616
rect 62836 349558 64939 349560
rect 89884 349616 91159 349618
rect 89884 349560 91098 349616
rect 91154 349560 91159 349616
rect 89884 349558 91159 349560
rect 116932 349616 118759 349618
rect 116932 349560 118698 349616
rect 118754 349560 118759 349616
rect 170844 349616 172579 349618
rect 116932 349558 118759 349560
rect 64873 349555 64939 349558
rect 91093 349555 91159 349558
rect 118693 349555 118759 349558
rect 37917 349210 37983 349213
rect 35758 349208 37983 349210
rect 35758 349152 37922 349208
rect 37978 349152 37983 349208
rect 35758 349150 37983 349152
rect 143766 349210 143826 349588
rect 170844 349560 172518 349616
rect 172574 349560 172579 349616
rect 170844 349558 172579 349560
rect 197892 349616 200179 349618
rect 197892 349560 200118 349616
rect 200174 349560 200179 349616
rect 197892 349558 200179 349560
rect 224940 349616 226399 349618
rect 224940 349560 226338 349616
rect 226394 349560 226399 349616
rect 278852 349616 280219 349618
rect 224940 349558 226399 349560
rect 172513 349555 172579 349558
rect 200113 349555 200179 349558
rect 226333 349555 226399 349558
rect 146293 349210 146359 349213
rect 143766 349208 146359 349210
rect 143766 349152 146298 349208
rect 146354 349152 146359 349208
rect 143766 349150 146359 349152
rect 251774 349210 251834 349588
rect 278852 349560 280158 349616
rect 280214 349560 280219 349616
rect 278852 349558 280219 349560
rect 305900 349616 307819 349618
rect 305900 349560 307758 349616
rect 307814 349560 307819 349616
rect 305900 349558 307819 349560
rect 332948 349616 335419 349618
rect 332948 349560 335358 349616
rect 335414 349560 335419 349616
rect 386860 349616 389239 349618
rect 332948 349558 335419 349560
rect 280153 349555 280219 349558
rect 307753 349555 307819 349558
rect 335353 349555 335419 349558
rect 253933 349210 253999 349213
rect 251774 349208 253999 349210
rect 251774 349152 253938 349208
rect 253994 349152 253999 349208
rect 251774 349150 253999 349152
rect 359782 349210 359842 349588
rect 386860 349560 389178 349616
rect 389234 349560 389239 349616
rect 386860 349558 389239 349560
rect 413908 349616 415459 349618
rect 413908 349560 415398 349616
rect 415454 349560 415459 349616
rect 413908 349558 415459 349560
rect 440956 349616 443059 349618
rect 440956 349560 442998 349616
rect 443054 349560 443059 349616
rect 494868 349616 496879 349618
rect 440956 349558 443059 349560
rect 389173 349555 389239 349558
rect 415393 349555 415459 349558
rect 442993 349555 443059 349558
rect 361573 349210 361639 349213
rect 359782 349208 361639 349210
rect 359782 349152 361578 349208
rect 361634 349152 361639 349208
rect 359782 349150 361639 349152
rect 467790 349210 467850 349588
rect 494868 349560 496818 349616
rect 496874 349560 496879 349616
rect 494868 349558 496879 349560
rect 521916 349616 523099 349618
rect 521916 349560 523038 349616
rect 523094 349560 523099 349616
rect 521916 349558 523099 349560
rect 548964 349616 550699 349618
rect 548964 349560 550638 349616
rect 550694 349560 550699 349616
rect 548964 349558 550699 349560
rect 496813 349555 496879 349558
rect 523033 349555 523099 349558
rect 550633 349555 550699 349558
rect 469213 349210 469279 349213
rect 467790 349208 469279 349210
rect 467790 349152 469218 349208
rect 469274 349152 469279 349208
rect 467790 349150 469279 349152
rect 37917 349147 37983 349150
rect 146293 349147 146359 349150
rect 253933 349147 253999 349150
rect 361573 349147 361639 349150
rect 469213 349147 469279 349150
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect 526437 323370 526503 323373
rect 526437 323368 529092 323370
rect 526437 323312 526442 323368
rect 526498 323312 529092 323368
rect 526437 323310 529092 323312
rect 526437 323307 526503 323310
rect 13721 323234 13787 323237
rect 41321 323234 41387 323237
rect 95141 323234 95207 323237
rect 122741 323234 122807 323237
rect 148961 323234 149027 323237
rect 202781 323234 202847 323237
rect 230381 323234 230447 323237
rect 256601 323234 256667 323237
rect 311801 323234 311867 323237
rect 338021 323234 338087 323237
rect 365621 323234 365687 323237
rect 391841 323234 391907 323237
rect 419441 323234 419507 323237
rect 445661 323234 445727 323237
rect 500861 323234 500927 323237
rect 13721 323232 16100 323234
rect 13721 323176 13726 323232
rect 13782 323176 16100 323232
rect 13721 323174 16100 323176
rect 41321 323232 43148 323234
rect 41321 323176 41326 323232
rect 41382 323176 43148 323232
rect 95141 323232 97060 323234
rect 41321 323174 43148 323176
rect 13721 323171 13787 323174
rect 41321 323171 41387 323174
rect 68921 322962 68987 322965
rect 70166 322962 70226 323204
rect 95141 323176 95146 323232
rect 95202 323176 97060 323232
rect 95141 323174 97060 323176
rect 122741 323232 124108 323234
rect 122741 323176 122746 323232
rect 122802 323176 124108 323232
rect 122741 323174 124108 323176
rect 148961 323232 151156 323234
rect 148961 323176 148966 323232
rect 149022 323176 151156 323232
rect 202781 323232 205068 323234
rect 148961 323174 151156 323176
rect 95141 323171 95207 323174
rect 122741 323171 122807 323174
rect 148961 323171 149027 323174
rect 68921 322960 70226 322962
rect 68921 322904 68926 322960
rect 68982 322904 70226 322960
rect 68921 322902 70226 322904
rect 176561 322962 176627 322965
rect 178174 322962 178234 323204
rect 202781 323176 202786 323232
rect 202842 323176 205068 323232
rect 202781 323174 205068 323176
rect 230381 323232 232116 323234
rect 230381 323176 230386 323232
rect 230442 323176 232116 323232
rect 230381 323174 232116 323176
rect 256601 323232 259164 323234
rect 256601 323176 256606 323232
rect 256662 323176 259164 323232
rect 311801 323232 313076 323234
rect 256601 323174 259164 323176
rect 202781 323171 202847 323174
rect 230381 323171 230447 323174
rect 256601 323171 256667 323174
rect 176561 322960 178234 322962
rect 176561 322904 176566 322960
rect 176622 322904 178234 322960
rect 176561 322902 178234 322904
rect 284201 322962 284267 322965
rect 286182 322962 286242 323204
rect 311801 323176 311806 323232
rect 311862 323176 313076 323232
rect 311801 323174 313076 323176
rect 338021 323232 340124 323234
rect 338021 323176 338026 323232
rect 338082 323176 340124 323232
rect 338021 323174 340124 323176
rect 365621 323232 367172 323234
rect 365621 323176 365626 323232
rect 365682 323176 367172 323232
rect 365621 323174 367172 323176
rect 391841 323232 394036 323234
rect 391841 323176 391846 323232
rect 391902 323176 394036 323232
rect 391841 323174 394036 323176
rect 419441 323232 421084 323234
rect 419441 323176 419446 323232
rect 419502 323176 421084 323232
rect 419441 323174 421084 323176
rect 445661 323232 448132 323234
rect 445661 323176 445666 323232
rect 445722 323176 448132 323232
rect 500861 323232 502044 323234
rect 445661 323174 448132 323176
rect 311801 323171 311867 323174
rect 338021 323171 338087 323174
rect 365621 323171 365687 323174
rect 391841 323171 391907 323174
rect 419441 323171 419507 323174
rect 445661 323171 445727 323174
rect 284201 322960 286242 322962
rect 284201 322904 284206 322960
rect 284262 322904 286242 322960
rect 284201 322902 286242 322904
rect 473261 322962 473327 322965
rect 475150 322962 475210 323204
rect 500861 323176 500866 323232
rect 500922 323176 502044 323232
rect 500861 323174 502044 323176
rect 500861 323171 500927 323174
rect 473261 322960 475210 322962
rect 473261 322904 473266 322960
rect 473322 322904 475210 322960
rect 473261 322902 475210 322904
rect 68921 322899 68987 322902
rect 176561 322899 176627 322902
rect 284201 322899 284267 322902
rect 473261 322899 473327 322902
rect 64873 322554 64939 322557
rect 91093 322554 91159 322557
rect 118693 322554 118759 322557
rect 172513 322554 172579 322557
rect 200113 322554 200179 322557
rect 226333 322554 226399 322557
rect 280153 322554 280219 322557
rect 307753 322554 307819 322557
rect 335353 322554 335419 322557
rect 389173 322554 389239 322557
rect 415393 322554 415459 322557
rect 442993 322554 443059 322557
rect 496813 322554 496879 322557
rect 523033 322554 523099 322557
rect 550633 322554 550699 322557
rect 62836 322552 64939 322554
rect 35758 322010 35818 322524
rect 62836 322496 64878 322552
rect 64934 322496 64939 322552
rect 62836 322494 64939 322496
rect 89884 322552 91159 322554
rect 89884 322496 91098 322552
rect 91154 322496 91159 322552
rect 89884 322494 91159 322496
rect 116932 322552 118759 322554
rect 116932 322496 118698 322552
rect 118754 322496 118759 322552
rect 170844 322552 172579 322554
rect 116932 322494 118759 322496
rect 64873 322491 64939 322494
rect 91093 322491 91159 322494
rect 118693 322491 118759 322494
rect 37917 322010 37983 322013
rect 35758 322008 37983 322010
rect 35758 321952 37922 322008
rect 37978 321952 37983 322008
rect 35758 321950 37983 321952
rect 143766 322010 143826 322524
rect 170844 322496 172518 322552
rect 172574 322496 172579 322552
rect 170844 322494 172579 322496
rect 197892 322552 200179 322554
rect 197892 322496 200118 322552
rect 200174 322496 200179 322552
rect 197892 322494 200179 322496
rect 224940 322552 226399 322554
rect 224940 322496 226338 322552
rect 226394 322496 226399 322552
rect 278852 322552 280219 322554
rect 224940 322494 226399 322496
rect 172513 322491 172579 322494
rect 200113 322491 200179 322494
rect 226333 322491 226399 322494
rect 146293 322010 146359 322013
rect 143766 322008 146359 322010
rect 143766 321952 146298 322008
rect 146354 321952 146359 322008
rect 143766 321950 146359 321952
rect 251774 322010 251834 322524
rect 278852 322496 280158 322552
rect 280214 322496 280219 322552
rect 278852 322494 280219 322496
rect 305900 322552 307819 322554
rect 305900 322496 307758 322552
rect 307814 322496 307819 322552
rect 305900 322494 307819 322496
rect 332948 322552 335419 322554
rect 332948 322496 335358 322552
rect 335414 322496 335419 322552
rect 386860 322552 389239 322554
rect 332948 322494 335419 322496
rect 280153 322491 280219 322494
rect 307753 322491 307819 322494
rect 335353 322491 335419 322494
rect 253933 322010 253999 322013
rect 251774 322008 253999 322010
rect 251774 321952 253938 322008
rect 253994 321952 253999 322008
rect 251774 321950 253999 321952
rect 359782 322010 359842 322524
rect 386860 322496 389178 322552
rect 389234 322496 389239 322552
rect 386860 322494 389239 322496
rect 413908 322552 415459 322554
rect 413908 322496 415398 322552
rect 415454 322496 415459 322552
rect 413908 322494 415459 322496
rect 440956 322552 443059 322554
rect 440956 322496 442998 322552
rect 443054 322496 443059 322552
rect 494868 322552 496879 322554
rect 440956 322494 443059 322496
rect 389173 322491 389239 322494
rect 415393 322491 415459 322494
rect 442993 322491 443059 322494
rect 361573 322010 361639 322013
rect 359782 322008 361639 322010
rect 359782 321952 361578 322008
rect 361634 321952 361639 322008
rect 359782 321950 361639 321952
rect 467790 322010 467850 322524
rect 494868 322496 496818 322552
rect 496874 322496 496879 322552
rect 494868 322494 496879 322496
rect 521916 322552 523099 322554
rect 521916 322496 523038 322552
rect 523094 322496 523099 322552
rect 521916 322494 523099 322496
rect 548964 322552 550699 322554
rect 548964 322496 550638 322552
rect 550694 322496 550699 322552
rect 548964 322494 550699 322496
rect 496813 322491 496879 322494
rect 523033 322491 523099 322494
rect 550633 322491 550699 322494
rect 469213 322010 469279 322013
rect 467790 322008 469279 322010
rect 467790 321952 469218 322008
rect 469274 321952 469279 322008
rect 467790 321950 469279 321952
rect 37917 321947 37983 321950
rect 146293 321947 146359 321950
rect 253933 321947 253999 321950
rect 361573 321947 361639 321950
rect 469213 321947 469279 321950
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 583520 298604 584960 298844
rect 13721 296306 13787 296309
rect 41321 296306 41387 296309
rect 95141 296306 95207 296309
rect 122741 296306 122807 296309
rect 148961 296306 149027 296309
rect 202781 296306 202847 296309
rect 230381 296306 230447 296309
rect 256601 296306 256667 296309
rect 311801 296306 311867 296309
rect 338021 296306 338087 296309
rect 365621 296306 365687 296309
rect 391841 296306 391907 296309
rect 419441 296306 419507 296309
rect 445661 296306 445727 296309
rect 500861 296306 500927 296309
rect 526437 296306 526503 296309
rect 13721 296304 16100 296306
rect 13721 296248 13726 296304
rect 13782 296248 16100 296304
rect 13721 296246 16100 296248
rect 41321 296304 43148 296306
rect 41321 296248 41326 296304
rect 41382 296248 43148 296304
rect 95141 296304 97060 296306
rect 41321 296246 43148 296248
rect 13721 296243 13787 296246
rect 41321 296243 41387 296246
rect 68921 295762 68987 295765
rect 70166 295762 70226 296276
rect 95141 296248 95146 296304
rect 95202 296248 97060 296304
rect 95141 296246 97060 296248
rect 122741 296304 124108 296306
rect 122741 296248 122746 296304
rect 122802 296248 124108 296304
rect 122741 296246 124108 296248
rect 148961 296304 151156 296306
rect 148961 296248 148966 296304
rect 149022 296248 151156 296304
rect 202781 296304 205068 296306
rect 148961 296246 151156 296248
rect 95141 296243 95207 296246
rect 122741 296243 122807 296246
rect 148961 296243 149027 296246
rect 68921 295760 70226 295762
rect 68921 295704 68926 295760
rect 68982 295704 70226 295760
rect 68921 295702 70226 295704
rect 176561 295762 176627 295765
rect 178174 295762 178234 296276
rect 202781 296248 202786 296304
rect 202842 296248 205068 296304
rect 202781 296246 205068 296248
rect 230381 296304 232116 296306
rect 230381 296248 230386 296304
rect 230442 296248 232116 296304
rect 230381 296246 232116 296248
rect 256601 296304 259164 296306
rect 256601 296248 256606 296304
rect 256662 296248 259164 296304
rect 311801 296304 313076 296306
rect 256601 296246 259164 296248
rect 202781 296243 202847 296246
rect 230381 296243 230447 296246
rect 256601 296243 256667 296246
rect 176561 295760 178234 295762
rect 176561 295704 176566 295760
rect 176622 295704 178234 295760
rect 176561 295702 178234 295704
rect 284201 295762 284267 295765
rect 286182 295762 286242 296276
rect 311801 296248 311806 296304
rect 311862 296248 313076 296304
rect 311801 296246 313076 296248
rect 338021 296304 340124 296306
rect 338021 296248 338026 296304
rect 338082 296248 340124 296304
rect 338021 296246 340124 296248
rect 365621 296304 367172 296306
rect 365621 296248 365626 296304
rect 365682 296248 367172 296304
rect 365621 296246 367172 296248
rect 391841 296304 394036 296306
rect 391841 296248 391846 296304
rect 391902 296248 394036 296304
rect 391841 296246 394036 296248
rect 419441 296304 421084 296306
rect 419441 296248 419446 296304
rect 419502 296248 421084 296304
rect 419441 296246 421084 296248
rect 445661 296304 448132 296306
rect 445661 296248 445666 296304
rect 445722 296248 448132 296304
rect 500861 296304 502044 296306
rect 445661 296246 448132 296248
rect 311801 296243 311867 296246
rect 338021 296243 338087 296246
rect 365621 296243 365687 296246
rect 391841 296243 391907 296246
rect 419441 296243 419507 296246
rect 445661 296243 445727 296246
rect 284201 295760 286242 295762
rect 284201 295704 284206 295760
rect 284262 295704 286242 295760
rect 284201 295702 286242 295704
rect 473261 295762 473327 295765
rect 475150 295762 475210 296276
rect 500861 296248 500866 296304
rect 500922 296248 502044 296304
rect 500861 296246 502044 296248
rect 526437 296304 529092 296306
rect 526437 296248 526442 296304
rect 526498 296248 529092 296304
rect 526437 296246 529092 296248
rect 500861 296243 500927 296246
rect 526437 296243 526503 296246
rect 473261 295760 475210 295762
rect 473261 295704 473266 295760
rect 473322 295704 475210 295760
rect 473261 295702 475210 295704
rect 68921 295699 68987 295702
rect 176561 295699 176627 295702
rect 284201 295699 284267 295702
rect 473261 295699 473327 295702
rect 64873 295626 64939 295629
rect 91093 295626 91159 295629
rect 118693 295626 118759 295629
rect 172513 295626 172579 295629
rect 200113 295626 200179 295629
rect 226333 295626 226399 295629
rect 280153 295626 280219 295629
rect 307753 295626 307819 295629
rect 335353 295626 335419 295629
rect 389173 295626 389239 295629
rect 415393 295626 415459 295629
rect 442993 295626 443059 295629
rect 496813 295626 496879 295629
rect 523033 295626 523099 295629
rect 550633 295626 550699 295629
rect 62836 295624 64939 295626
rect 35758 295354 35818 295596
rect 62836 295568 64878 295624
rect 64934 295568 64939 295624
rect 62836 295566 64939 295568
rect 89884 295624 91159 295626
rect 89884 295568 91098 295624
rect 91154 295568 91159 295624
rect 89884 295566 91159 295568
rect 116932 295624 118759 295626
rect 116932 295568 118698 295624
rect 118754 295568 118759 295624
rect 170844 295624 172579 295626
rect 116932 295566 118759 295568
rect 64873 295563 64939 295566
rect 91093 295563 91159 295566
rect 118693 295563 118759 295566
rect 37917 295354 37983 295357
rect 35758 295352 37983 295354
rect 35758 295296 37922 295352
rect 37978 295296 37983 295352
rect 35758 295294 37983 295296
rect 143766 295354 143826 295596
rect 170844 295568 172518 295624
rect 172574 295568 172579 295624
rect 170844 295566 172579 295568
rect 197892 295624 200179 295626
rect 197892 295568 200118 295624
rect 200174 295568 200179 295624
rect 197892 295566 200179 295568
rect 224940 295624 226399 295626
rect 224940 295568 226338 295624
rect 226394 295568 226399 295624
rect 278852 295624 280219 295626
rect 224940 295566 226399 295568
rect 172513 295563 172579 295566
rect 200113 295563 200179 295566
rect 226333 295563 226399 295566
rect 146293 295354 146359 295357
rect 143766 295352 146359 295354
rect 143766 295296 146298 295352
rect 146354 295296 146359 295352
rect 143766 295294 146359 295296
rect 251774 295354 251834 295596
rect 278852 295568 280158 295624
rect 280214 295568 280219 295624
rect 278852 295566 280219 295568
rect 305900 295624 307819 295626
rect 305900 295568 307758 295624
rect 307814 295568 307819 295624
rect 305900 295566 307819 295568
rect 332948 295624 335419 295626
rect 332948 295568 335358 295624
rect 335414 295568 335419 295624
rect 386860 295624 389239 295626
rect 332948 295566 335419 295568
rect 280153 295563 280219 295566
rect 307753 295563 307819 295566
rect 335353 295563 335419 295566
rect 253933 295354 253999 295357
rect 251774 295352 253999 295354
rect 251774 295296 253938 295352
rect 253994 295296 253999 295352
rect 251774 295294 253999 295296
rect 359782 295354 359842 295596
rect 386860 295568 389178 295624
rect 389234 295568 389239 295624
rect 386860 295566 389239 295568
rect 413908 295624 415459 295626
rect 413908 295568 415398 295624
rect 415454 295568 415459 295624
rect 413908 295566 415459 295568
rect 440956 295624 443059 295626
rect 440956 295568 442998 295624
rect 443054 295568 443059 295624
rect 494868 295624 496879 295626
rect 440956 295566 443059 295568
rect 389173 295563 389239 295566
rect 415393 295563 415459 295566
rect 442993 295563 443059 295566
rect 361573 295354 361639 295357
rect 359782 295352 361639 295354
rect 359782 295296 361578 295352
rect 361634 295296 361639 295352
rect 359782 295294 361639 295296
rect 467790 295354 467850 295596
rect 494868 295568 496818 295624
rect 496874 295568 496879 295624
rect 494868 295566 496879 295568
rect 521916 295624 523099 295626
rect 521916 295568 523038 295624
rect 523094 295568 523099 295624
rect 521916 295566 523099 295568
rect 548964 295624 550699 295626
rect 548964 295568 550638 295624
rect 550694 295568 550699 295624
rect 548964 295566 550699 295568
rect 496813 295563 496879 295566
rect 523033 295563 523099 295566
rect 550633 295563 550699 295566
rect 469213 295354 469279 295357
rect 467790 295352 469279 295354
rect 467790 295296 469218 295352
rect 469274 295296 469279 295352
rect 467790 295294 469279 295296
rect 37917 295291 37983 295294
rect 146293 295291 146359 295294
rect 253933 295291 253999 295294
rect 361573 295291 361639 295294
rect 469213 295291 469279 295294
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect 68921 269922 68987 269925
rect 176561 269922 176627 269925
rect 284201 269922 284267 269925
rect 473261 269922 473327 269925
rect 68921 269920 70226 269922
rect 68921 269864 68926 269920
rect 68982 269864 70226 269920
rect 68921 269862 70226 269864
rect 68921 269859 68987 269862
rect 13721 269378 13787 269381
rect 41321 269378 41387 269381
rect 13721 269376 16100 269378
rect 13721 269320 13726 269376
rect 13782 269320 16100 269376
rect 13721 269318 16100 269320
rect 41321 269376 43148 269378
rect 41321 269320 41326 269376
rect 41382 269320 43148 269376
rect 70166 269348 70226 269862
rect 176561 269920 178234 269922
rect 176561 269864 176566 269920
rect 176622 269864 178234 269920
rect 176561 269862 178234 269864
rect 176561 269859 176627 269862
rect 95141 269378 95207 269381
rect 122741 269378 122807 269381
rect 148961 269378 149027 269381
rect 95141 269376 97060 269378
rect 41321 269318 43148 269320
rect 95141 269320 95146 269376
rect 95202 269320 97060 269376
rect 95141 269318 97060 269320
rect 122741 269376 124108 269378
rect 122741 269320 122746 269376
rect 122802 269320 124108 269376
rect 122741 269318 124108 269320
rect 148961 269376 151156 269378
rect 148961 269320 148966 269376
rect 149022 269320 151156 269376
rect 178174 269348 178234 269862
rect 284201 269920 286242 269922
rect 284201 269864 284206 269920
rect 284262 269864 286242 269920
rect 284201 269862 286242 269864
rect 284201 269859 284267 269862
rect 202781 269378 202847 269381
rect 230381 269378 230447 269381
rect 256601 269378 256667 269381
rect 202781 269376 205068 269378
rect 148961 269318 151156 269320
rect 202781 269320 202786 269376
rect 202842 269320 205068 269376
rect 202781 269318 205068 269320
rect 230381 269376 232116 269378
rect 230381 269320 230386 269376
rect 230442 269320 232116 269376
rect 230381 269318 232116 269320
rect 256601 269376 259164 269378
rect 256601 269320 256606 269376
rect 256662 269320 259164 269376
rect 286182 269348 286242 269862
rect 473261 269920 475210 269922
rect 473261 269864 473266 269920
rect 473322 269864 475210 269920
rect 473261 269862 475210 269864
rect 473261 269859 473327 269862
rect 311801 269378 311867 269381
rect 338021 269378 338087 269381
rect 365621 269378 365687 269381
rect 391841 269378 391907 269381
rect 419441 269378 419507 269381
rect 445661 269378 445727 269381
rect 311801 269376 313076 269378
rect 256601 269318 259164 269320
rect 311801 269320 311806 269376
rect 311862 269320 313076 269376
rect 311801 269318 313076 269320
rect 338021 269376 340124 269378
rect 338021 269320 338026 269376
rect 338082 269320 340124 269376
rect 338021 269318 340124 269320
rect 365621 269376 367172 269378
rect 365621 269320 365626 269376
rect 365682 269320 367172 269376
rect 365621 269318 367172 269320
rect 391841 269376 394036 269378
rect 391841 269320 391846 269376
rect 391902 269320 394036 269376
rect 391841 269318 394036 269320
rect 419441 269376 421084 269378
rect 419441 269320 419446 269376
rect 419502 269320 421084 269376
rect 419441 269318 421084 269320
rect 445661 269376 448132 269378
rect 445661 269320 445666 269376
rect 445722 269320 448132 269376
rect 475150 269348 475210 269862
rect 500861 269378 500927 269381
rect 526437 269378 526503 269381
rect 500861 269376 502044 269378
rect 445661 269318 448132 269320
rect 500861 269320 500866 269376
rect 500922 269320 502044 269376
rect 500861 269318 502044 269320
rect 526437 269376 529092 269378
rect 526437 269320 526442 269376
rect 526498 269320 529092 269376
rect 526437 269318 529092 269320
rect 13721 269315 13787 269318
rect 41321 269315 41387 269318
rect 95141 269315 95207 269318
rect 122741 269315 122807 269318
rect 148961 269315 149027 269318
rect 202781 269315 202847 269318
rect 230381 269315 230447 269318
rect 256601 269315 256667 269318
rect 311801 269315 311867 269318
rect 338021 269315 338087 269318
rect 365621 269315 365687 269318
rect 391841 269315 391907 269318
rect 419441 269315 419507 269318
rect 445661 269315 445727 269318
rect 500861 269315 500927 269318
rect 526437 269315 526503 269318
rect 146293 269106 146359 269109
rect 253933 269106 253999 269109
rect 361573 269106 361639 269109
rect 469213 269106 469279 269109
rect 143766 269104 146359 269106
rect 143766 269048 146298 269104
rect 146354 269048 146359 269104
rect 143766 269046 146359 269048
rect 64873 268698 64939 268701
rect 91093 268698 91159 268701
rect 118693 268698 118759 268701
rect 62836 268696 64939 268698
rect 62836 268640 64878 268696
rect 64934 268640 64939 268696
rect 62836 268638 64939 268640
rect 89884 268696 91159 268698
rect 89884 268640 91098 268696
rect 91154 268640 91159 268696
rect 89884 268638 91159 268640
rect 116932 268696 118759 268698
rect 116932 268640 118698 268696
rect 118754 268640 118759 268696
rect 143766 268668 143826 269046
rect 146293 269043 146359 269046
rect 251774 269104 253999 269106
rect 251774 269048 253938 269104
rect 253994 269048 253999 269104
rect 251774 269046 253999 269048
rect 172513 268698 172579 268701
rect 200113 268698 200179 268701
rect 226333 268698 226399 268701
rect 170844 268696 172579 268698
rect 116932 268638 118759 268640
rect 170844 268640 172518 268696
rect 172574 268640 172579 268696
rect 170844 268638 172579 268640
rect 197892 268696 200179 268698
rect 197892 268640 200118 268696
rect 200174 268640 200179 268696
rect 197892 268638 200179 268640
rect 224940 268696 226399 268698
rect 224940 268640 226338 268696
rect 226394 268640 226399 268696
rect 251774 268668 251834 269046
rect 253933 269043 253999 269046
rect 359782 269104 361639 269106
rect 359782 269048 361578 269104
rect 361634 269048 361639 269104
rect 359782 269046 361639 269048
rect 280153 268698 280219 268701
rect 307753 268698 307819 268701
rect 335353 268698 335419 268701
rect 278852 268696 280219 268698
rect 224940 268638 226399 268640
rect 278852 268640 280158 268696
rect 280214 268640 280219 268696
rect 278852 268638 280219 268640
rect 305900 268696 307819 268698
rect 305900 268640 307758 268696
rect 307814 268640 307819 268696
rect 305900 268638 307819 268640
rect 332948 268696 335419 268698
rect 332948 268640 335358 268696
rect 335414 268640 335419 268696
rect 359782 268668 359842 269046
rect 361573 269043 361639 269046
rect 467790 269104 469279 269106
rect 467790 269048 469218 269104
rect 469274 269048 469279 269104
rect 467790 269046 469279 269048
rect 389173 268698 389239 268701
rect 415393 268698 415459 268701
rect 442993 268698 443059 268701
rect 386860 268696 389239 268698
rect 332948 268638 335419 268640
rect 386860 268640 389178 268696
rect 389234 268640 389239 268696
rect 386860 268638 389239 268640
rect 413908 268696 415459 268698
rect 413908 268640 415398 268696
rect 415454 268640 415459 268696
rect 413908 268638 415459 268640
rect 440956 268696 443059 268698
rect 440956 268640 442998 268696
rect 443054 268640 443059 268696
rect 467790 268668 467850 269046
rect 469213 269043 469279 269046
rect 496813 268698 496879 268701
rect 523033 268698 523099 268701
rect 550633 268698 550699 268701
rect 494868 268696 496879 268698
rect 440956 268638 443059 268640
rect 494868 268640 496818 268696
rect 496874 268640 496879 268696
rect 494868 268638 496879 268640
rect 521916 268696 523099 268698
rect 521916 268640 523038 268696
rect 523094 268640 523099 268696
rect 521916 268638 523099 268640
rect 548964 268696 550699 268698
rect 548964 268640 550638 268696
rect 550694 268640 550699 268696
rect 548964 268638 550699 268640
rect 64873 268635 64939 268638
rect 91093 268635 91159 268638
rect 118693 268635 118759 268638
rect 172513 268635 172579 268638
rect 200113 268635 200179 268638
rect 226333 268635 226399 268638
rect 280153 268635 280219 268638
rect 307753 268635 307819 268638
rect 335353 268635 335419 268638
rect 389173 268635 389239 268638
rect 415393 268635 415459 268638
rect 442993 268635 443059 268638
rect 496813 268635 496879 268638
rect 523033 268635 523099 268638
rect 550633 268635 550699 268638
rect 35758 268018 35818 268532
rect 37917 268018 37983 268021
rect 35758 268016 37983 268018
rect 35758 267960 37922 268016
rect 37978 267960 37983 268016
rect 35758 267958 37983 267960
rect 37917 267955 37983 267958
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect 68921 242858 68987 242861
rect 284201 242858 284267 242861
rect 473261 242858 473327 242861
rect 68921 242856 70226 242858
rect 68921 242800 68926 242856
rect 68982 242800 70226 242856
rect 68921 242798 70226 242800
rect 68921 242795 68987 242798
rect 41321 242314 41387 242317
rect 41321 242312 43148 242314
rect 41321 242256 41326 242312
rect 41382 242256 43148 242312
rect 70166 242284 70226 242798
rect 284201 242856 286242 242858
rect 284201 242800 284206 242856
rect 284262 242800 286242 242856
rect 284201 242798 286242 242800
rect 284201 242795 284267 242798
rect 122741 242314 122807 242317
rect 148961 242314 149027 242317
rect 202781 242314 202847 242317
rect 230381 242314 230447 242317
rect 122741 242312 124108 242314
rect 41321 242254 43148 242256
rect 122741 242256 122746 242312
rect 122802 242256 124108 242312
rect 122741 242254 124108 242256
rect 148961 242312 151156 242314
rect 148961 242256 148966 242312
rect 149022 242256 151156 242312
rect 148961 242254 151156 242256
rect 202781 242312 205068 242314
rect 202781 242256 202786 242312
rect 202842 242256 205068 242312
rect 202781 242254 205068 242256
rect 230381 242312 232116 242314
rect 230381 242256 230386 242312
rect 230442 242256 232116 242312
rect 286182 242284 286242 242798
rect 473261 242856 475210 242858
rect 473261 242800 473266 242856
rect 473322 242800 475210 242856
rect 473261 242798 475210 242800
rect 473261 242795 473327 242798
rect 311801 242314 311867 242317
rect 365621 242314 365687 242317
rect 419441 242314 419507 242317
rect 311801 242312 313076 242314
rect 230381 242254 232116 242256
rect 311801 242256 311806 242312
rect 311862 242256 313076 242312
rect 311801 242254 313076 242256
rect 365621 242312 367172 242314
rect 365621 242256 365626 242312
rect 365682 242256 367172 242312
rect 365621 242254 367172 242256
rect 419441 242312 421084 242314
rect 419441 242256 419446 242312
rect 419502 242256 421084 242312
rect 475150 242284 475210 242798
rect 500861 242314 500927 242317
rect 526437 242314 526503 242317
rect 500861 242312 502044 242314
rect 419441 242254 421084 242256
rect 500861 242256 500866 242312
rect 500922 242256 502044 242312
rect 500861 242254 502044 242256
rect 526437 242312 529092 242314
rect 526437 242256 526442 242312
rect 526498 242256 529092 242312
rect 526437 242254 529092 242256
rect 41321 242251 41387 242254
rect 122741 242251 122807 242254
rect 148961 242251 149027 242254
rect 202781 242251 202847 242254
rect 230381 242251 230447 242254
rect 311801 242251 311867 242254
rect 365621 242251 365687 242254
rect 419441 242251 419507 242254
rect 500861 242251 500927 242254
rect 526437 242251 526503 242254
rect 13721 242178 13787 242181
rect 95141 242178 95207 242181
rect 253933 242178 253999 242181
rect 13721 242176 16100 242178
rect 13721 242120 13726 242176
rect 13782 242120 16100 242176
rect 13721 242118 16100 242120
rect 95141 242176 97060 242178
rect 95141 242120 95146 242176
rect 95202 242120 97060 242176
rect 251774 242176 253999 242178
rect 95141 242118 97060 242120
rect 13721 242115 13787 242118
rect 95141 242115 95207 242118
rect 37917 241906 37983 241909
rect 146293 241906 146359 241909
rect 35758 241904 37983 241906
rect 35758 241848 37922 241904
rect 37978 241848 37983 241904
rect 35758 241846 37983 241848
rect 35758 241604 35818 241846
rect 37917 241843 37983 241846
rect 143582 241904 146359 241906
rect 143582 241848 146298 241904
rect 146354 241848 146359 241904
rect 143582 241846 146359 241848
rect 64873 241634 64939 241637
rect 91093 241634 91159 241637
rect 118693 241634 118759 241637
rect 62836 241632 64939 241634
rect 62836 241576 64878 241632
rect 64934 241576 64939 241632
rect 62836 241574 64939 241576
rect 89884 241632 91159 241634
rect 89884 241576 91098 241632
rect 91154 241576 91159 241632
rect 89884 241574 91159 241576
rect 116932 241632 118759 241634
rect 116932 241576 118698 241632
rect 118754 241576 118759 241632
rect 143582 241604 143642 241846
rect 146293 241843 146359 241846
rect 172513 241634 172579 241637
rect 170844 241632 172579 241634
rect 116932 241574 118759 241576
rect 170844 241576 172518 241632
rect 172574 241576 172579 241632
rect 170844 241574 172579 241576
rect 64873 241571 64939 241574
rect 91093 241571 91159 241574
rect 118693 241571 118759 241574
rect 172513 241571 172579 241574
rect 176561 241634 176627 241637
rect 178174 241634 178234 242148
rect 251774 242120 253938 242176
rect 253994 242120 253999 242176
rect 251774 242118 253999 242120
rect 200113 241634 200179 241637
rect 226333 241634 226399 241637
rect 176561 241632 178234 241634
rect 176561 241576 176566 241632
rect 176622 241576 178234 241632
rect 176561 241574 178234 241576
rect 197892 241632 200179 241634
rect 197892 241576 200118 241632
rect 200174 241576 200179 241632
rect 197892 241574 200179 241576
rect 224940 241632 226399 241634
rect 224940 241576 226338 241632
rect 226394 241576 226399 241632
rect 251774 241604 251834 242118
rect 253933 242115 253999 242118
rect 256601 242178 256667 242181
rect 338021 242178 338087 242181
rect 361573 242178 361639 242181
rect 256601 242176 259164 242178
rect 256601 242120 256606 242176
rect 256662 242120 259164 242176
rect 256601 242118 259164 242120
rect 338021 242176 340124 242178
rect 338021 242120 338026 242176
rect 338082 242120 340124 242176
rect 338021 242118 340124 242120
rect 359782 242176 361639 242178
rect 359782 242120 361578 242176
rect 361634 242120 361639 242176
rect 445661 242178 445727 242181
rect 469213 242178 469279 242181
rect 445661 242176 448132 242178
rect 359782 242118 361639 242120
rect 256601 242115 256667 242118
rect 338021 242115 338087 242118
rect 280153 241634 280219 241637
rect 307753 241634 307819 241637
rect 335353 241634 335419 241637
rect 278852 241632 280219 241634
rect 224940 241574 226399 241576
rect 278852 241576 280158 241632
rect 280214 241576 280219 241632
rect 278852 241574 280219 241576
rect 305900 241632 307819 241634
rect 305900 241576 307758 241632
rect 307814 241576 307819 241632
rect 305900 241574 307819 241576
rect 332948 241632 335419 241634
rect 332948 241576 335358 241632
rect 335414 241576 335419 241632
rect 359782 241604 359842 242118
rect 361573 242115 361639 242118
rect 391841 241906 391907 241909
rect 394006 241906 394066 242148
rect 445661 242120 445666 242176
rect 445722 242120 448132 242176
rect 445661 242118 448132 242120
rect 467790 242176 469279 242178
rect 467790 242120 469218 242176
rect 469274 242120 469279 242176
rect 467790 242118 469279 242120
rect 445661 242115 445727 242118
rect 391841 241904 394066 241906
rect 391841 241848 391846 241904
rect 391902 241848 394066 241904
rect 391841 241846 394066 241848
rect 391841 241843 391907 241846
rect 389173 241634 389239 241637
rect 415393 241634 415459 241637
rect 442993 241634 443059 241637
rect 386860 241632 389239 241634
rect 332948 241574 335419 241576
rect 386860 241576 389178 241632
rect 389234 241576 389239 241632
rect 386860 241574 389239 241576
rect 413908 241632 415459 241634
rect 413908 241576 415398 241632
rect 415454 241576 415459 241632
rect 413908 241574 415459 241576
rect 440956 241632 443059 241634
rect 440956 241576 442998 241632
rect 443054 241576 443059 241632
rect 467790 241604 467850 242118
rect 469213 242115 469279 242118
rect 496813 241634 496879 241637
rect 523033 241634 523099 241637
rect 550633 241634 550699 241637
rect 494868 241632 496879 241634
rect 440956 241574 443059 241576
rect 494868 241576 496818 241632
rect 496874 241576 496879 241632
rect 494868 241574 496879 241576
rect 521916 241632 523099 241634
rect 521916 241576 523038 241632
rect 523094 241576 523099 241632
rect 521916 241574 523099 241576
rect 548964 241632 550699 241634
rect 548964 241576 550638 241632
rect 550694 241576 550699 241632
rect 548964 241574 550699 241576
rect 176561 241571 176627 241574
rect 200113 241571 200179 241574
rect 226333 241571 226399 241574
rect 280153 241571 280219 241574
rect 307753 241571 307819 241574
rect 335353 241571 335419 241574
rect 389173 241571 389239 241574
rect 415393 241571 415459 241574
rect 442993 241571 443059 241574
rect 496813 241571 496879 241574
rect 523033 241571 523099 241574
rect 550633 241571 550699 241574
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect 13721 215250 13787 215253
rect 41321 215250 41387 215253
rect 95141 215250 95207 215253
rect 122741 215250 122807 215253
rect 148961 215250 149027 215253
rect 202781 215250 202847 215253
rect 230381 215250 230447 215253
rect 256601 215250 256667 215253
rect 311801 215250 311867 215253
rect 338021 215250 338087 215253
rect 365621 215250 365687 215253
rect 391841 215250 391907 215253
rect 419441 215250 419507 215253
rect 445661 215250 445727 215253
rect 500861 215250 500927 215253
rect 526437 215250 526503 215253
rect 13721 215248 16100 215250
rect 13721 215192 13726 215248
rect 13782 215192 16100 215248
rect 13721 215190 16100 215192
rect 41321 215248 43148 215250
rect 41321 215192 41326 215248
rect 41382 215192 43148 215248
rect 95141 215248 97060 215250
rect 41321 215190 43148 215192
rect 13721 215187 13787 215190
rect 41321 215187 41387 215190
rect -960 214828 480 215068
rect 68921 214706 68987 214709
rect 70166 214706 70226 215220
rect 95141 215192 95146 215248
rect 95202 215192 97060 215248
rect 95141 215190 97060 215192
rect 122741 215248 124108 215250
rect 122741 215192 122746 215248
rect 122802 215192 124108 215248
rect 122741 215190 124108 215192
rect 148961 215248 151156 215250
rect 148961 215192 148966 215248
rect 149022 215192 151156 215248
rect 202781 215248 205068 215250
rect 148961 215190 151156 215192
rect 95141 215187 95207 215190
rect 122741 215187 122807 215190
rect 148961 215187 149027 215190
rect 68921 214704 70226 214706
rect 68921 214648 68926 214704
rect 68982 214648 70226 214704
rect 68921 214646 70226 214648
rect 176561 214706 176627 214709
rect 178174 214706 178234 215220
rect 202781 215192 202786 215248
rect 202842 215192 205068 215248
rect 202781 215190 205068 215192
rect 230381 215248 232116 215250
rect 230381 215192 230386 215248
rect 230442 215192 232116 215248
rect 230381 215190 232116 215192
rect 256601 215248 259164 215250
rect 256601 215192 256606 215248
rect 256662 215192 259164 215248
rect 311801 215248 313076 215250
rect 256601 215190 259164 215192
rect 202781 215187 202847 215190
rect 230381 215187 230447 215190
rect 256601 215187 256667 215190
rect 176561 214704 178234 214706
rect 176561 214648 176566 214704
rect 176622 214648 178234 214704
rect 176561 214646 178234 214648
rect 284201 214706 284267 214709
rect 286182 214706 286242 215220
rect 311801 215192 311806 215248
rect 311862 215192 313076 215248
rect 311801 215190 313076 215192
rect 338021 215248 340124 215250
rect 338021 215192 338026 215248
rect 338082 215192 340124 215248
rect 338021 215190 340124 215192
rect 365621 215248 367172 215250
rect 365621 215192 365626 215248
rect 365682 215192 367172 215248
rect 365621 215190 367172 215192
rect 391841 215248 394036 215250
rect 391841 215192 391846 215248
rect 391902 215192 394036 215248
rect 391841 215190 394036 215192
rect 419441 215248 421084 215250
rect 419441 215192 419446 215248
rect 419502 215192 421084 215248
rect 419441 215190 421084 215192
rect 445661 215248 448132 215250
rect 445661 215192 445666 215248
rect 445722 215192 448132 215248
rect 500861 215248 502044 215250
rect 445661 215190 448132 215192
rect 311801 215187 311867 215190
rect 338021 215187 338087 215190
rect 365621 215187 365687 215190
rect 391841 215187 391907 215190
rect 419441 215187 419507 215190
rect 445661 215187 445727 215190
rect 284201 214704 286242 214706
rect 284201 214648 284206 214704
rect 284262 214648 286242 214704
rect 284201 214646 286242 214648
rect 473261 214706 473327 214709
rect 475150 214706 475210 215220
rect 500861 215192 500866 215248
rect 500922 215192 502044 215248
rect 500861 215190 502044 215192
rect 526437 215248 529092 215250
rect 526437 215192 526442 215248
rect 526498 215192 529092 215248
rect 526437 215190 529092 215192
rect 500861 215187 500927 215190
rect 526437 215187 526503 215190
rect 473261 214704 475210 214706
rect 473261 214648 473266 214704
rect 473322 214648 475210 214704
rect 473261 214646 475210 214648
rect 68921 214643 68987 214646
rect 176561 214643 176627 214646
rect 284201 214643 284267 214646
rect 473261 214643 473327 214646
rect 64873 214570 64939 214573
rect 91093 214570 91159 214573
rect 118693 214570 118759 214573
rect 172513 214570 172579 214573
rect 200113 214570 200179 214573
rect 226333 214570 226399 214573
rect 280153 214570 280219 214573
rect 307753 214570 307819 214573
rect 335353 214570 335419 214573
rect 389173 214570 389239 214573
rect 415393 214570 415459 214573
rect 442993 214570 443059 214573
rect 496813 214570 496879 214573
rect 523033 214570 523099 214573
rect 550633 214570 550699 214573
rect 62836 214568 64939 214570
rect 35758 214026 35818 214540
rect 62836 214512 64878 214568
rect 64934 214512 64939 214568
rect 62836 214510 64939 214512
rect 89884 214568 91159 214570
rect 89884 214512 91098 214568
rect 91154 214512 91159 214568
rect 89884 214510 91159 214512
rect 116932 214568 118759 214570
rect 116932 214512 118698 214568
rect 118754 214512 118759 214568
rect 170844 214568 172579 214570
rect 116932 214510 118759 214512
rect 64873 214507 64939 214510
rect 91093 214507 91159 214510
rect 118693 214507 118759 214510
rect 37917 214026 37983 214029
rect 35758 214024 37983 214026
rect 35758 213968 37922 214024
rect 37978 213968 37983 214024
rect 35758 213966 37983 213968
rect 143766 214026 143826 214540
rect 170844 214512 172518 214568
rect 172574 214512 172579 214568
rect 170844 214510 172579 214512
rect 197892 214568 200179 214570
rect 197892 214512 200118 214568
rect 200174 214512 200179 214568
rect 197892 214510 200179 214512
rect 224940 214568 226399 214570
rect 224940 214512 226338 214568
rect 226394 214512 226399 214568
rect 278852 214568 280219 214570
rect 224940 214510 226399 214512
rect 172513 214507 172579 214510
rect 200113 214507 200179 214510
rect 226333 214507 226399 214510
rect 146293 214026 146359 214029
rect 143766 214024 146359 214026
rect 143766 213968 146298 214024
rect 146354 213968 146359 214024
rect 143766 213966 146359 213968
rect 251774 214026 251834 214540
rect 278852 214512 280158 214568
rect 280214 214512 280219 214568
rect 278852 214510 280219 214512
rect 305900 214568 307819 214570
rect 305900 214512 307758 214568
rect 307814 214512 307819 214568
rect 305900 214510 307819 214512
rect 332948 214568 335419 214570
rect 332948 214512 335358 214568
rect 335414 214512 335419 214568
rect 386860 214568 389239 214570
rect 332948 214510 335419 214512
rect 280153 214507 280219 214510
rect 307753 214507 307819 214510
rect 335353 214507 335419 214510
rect 253933 214026 253999 214029
rect 251774 214024 253999 214026
rect 251774 213968 253938 214024
rect 253994 213968 253999 214024
rect 251774 213966 253999 213968
rect 359782 214026 359842 214540
rect 386860 214512 389178 214568
rect 389234 214512 389239 214568
rect 386860 214510 389239 214512
rect 413908 214568 415459 214570
rect 413908 214512 415398 214568
rect 415454 214512 415459 214568
rect 413908 214510 415459 214512
rect 440956 214568 443059 214570
rect 440956 214512 442998 214568
rect 443054 214512 443059 214568
rect 494868 214568 496879 214570
rect 440956 214510 443059 214512
rect 389173 214507 389239 214510
rect 415393 214507 415459 214510
rect 442993 214507 443059 214510
rect 361573 214026 361639 214029
rect 359782 214024 361639 214026
rect 359782 213968 361578 214024
rect 361634 213968 361639 214024
rect 359782 213966 361639 213968
rect 467790 214026 467850 214540
rect 494868 214512 496818 214568
rect 496874 214512 496879 214568
rect 494868 214510 496879 214512
rect 521916 214568 523099 214570
rect 521916 214512 523038 214568
rect 523094 214512 523099 214568
rect 521916 214510 523099 214512
rect 548964 214568 550699 214570
rect 548964 214512 550638 214568
rect 550694 214512 550699 214568
rect 548964 214510 550699 214512
rect 496813 214507 496879 214510
rect 523033 214507 523099 214510
rect 550633 214507 550699 214510
rect 469213 214026 469279 214029
rect 467790 214024 469279 214026
rect 467790 213968 469218 214024
rect 469274 213968 469279 214024
rect 467790 213966 469279 213968
rect 37917 213963 37983 213966
rect 146293 213963 146359 213966
rect 253933 213963 253999 213966
rect 361573 213963 361639 213966
rect 469213 213963 469279 213966
rect 583520 205580 584960 205820
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 526437 188322 526503 188325
rect 526437 188320 529092 188322
rect 526437 188264 526442 188320
rect 526498 188264 529092 188320
rect 526437 188262 529092 188264
rect 526437 188259 526503 188262
rect 13721 188186 13787 188189
rect 41321 188186 41387 188189
rect 95141 188186 95207 188189
rect 122741 188186 122807 188189
rect 148961 188186 149027 188189
rect 202781 188186 202847 188189
rect 230381 188186 230447 188189
rect 256601 188186 256667 188189
rect 311801 188186 311867 188189
rect 338021 188186 338087 188189
rect 365621 188186 365687 188189
rect 419441 188186 419507 188189
rect 445661 188186 445727 188189
rect 13721 188184 16100 188186
rect 13721 188128 13726 188184
rect 13782 188128 16100 188184
rect 13721 188126 16100 188128
rect 41321 188184 43148 188186
rect 41321 188128 41326 188184
rect 41382 188128 43148 188184
rect 95141 188184 97060 188186
rect 41321 188126 43148 188128
rect 13721 188123 13787 188126
rect 41321 188123 41387 188126
rect 68921 187778 68987 187781
rect 70166 187778 70226 188156
rect 95141 188128 95146 188184
rect 95202 188128 97060 188184
rect 95141 188126 97060 188128
rect 122741 188184 124108 188186
rect 122741 188128 122746 188184
rect 122802 188128 124108 188184
rect 122741 188126 124108 188128
rect 148961 188184 151156 188186
rect 148961 188128 148966 188184
rect 149022 188128 151156 188184
rect 202781 188184 205068 188186
rect 148961 188126 151156 188128
rect 95141 188123 95207 188126
rect 122741 188123 122807 188126
rect 148961 188123 149027 188126
rect 68921 187776 70226 187778
rect 68921 187720 68926 187776
rect 68982 187720 70226 187776
rect 68921 187718 70226 187720
rect 176561 187778 176627 187781
rect 178174 187778 178234 188156
rect 202781 188128 202786 188184
rect 202842 188128 205068 188184
rect 202781 188126 205068 188128
rect 230381 188184 232116 188186
rect 230381 188128 230386 188184
rect 230442 188128 232116 188184
rect 230381 188126 232116 188128
rect 256601 188184 259164 188186
rect 256601 188128 256606 188184
rect 256662 188128 259164 188184
rect 311801 188184 313076 188186
rect 256601 188126 259164 188128
rect 202781 188123 202847 188126
rect 230381 188123 230447 188126
rect 256601 188123 256667 188126
rect 176561 187776 178234 187778
rect 176561 187720 176566 187776
rect 176622 187720 178234 187776
rect 176561 187718 178234 187720
rect 284201 187778 284267 187781
rect 286182 187778 286242 188156
rect 311801 188128 311806 188184
rect 311862 188128 313076 188184
rect 311801 188126 313076 188128
rect 338021 188184 340124 188186
rect 338021 188128 338026 188184
rect 338082 188128 340124 188184
rect 338021 188126 340124 188128
rect 365621 188184 367172 188186
rect 365621 188128 365626 188184
rect 365682 188128 367172 188184
rect 419441 188184 421084 188186
rect 365621 188126 367172 188128
rect 311801 188123 311867 188126
rect 338021 188123 338087 188126
rect 365621 188123 365687 188126
rect 284201 187776 286242 187778
rect 284201 187720 284206 187776
rect 284262 187720 286242 187776
rect 284201 187718 286242 187720
rect 391841 187778 391907 187781
rect 394006 187778 394066 188156
rect 419441 188128 419446 188184
rect 419502 188128 421084 188184
rect 419441 188126 421084 188128
rect 445661 188184 448132 188186
rect 445661 188128 445666 188184
rect 445722 188128 448132 188184
rect 445661 188126 448132 188128
rect 419441 188123 419507 188126
rect 445661 188123 445727 188126
rect 391841 187776 394066 187778
rect 391841 187720 391846 187776
rect 391902 187720 394066 187776
rect 391841 187718 394066 187720
rect 473261 187778 473327 187781
rect 475150 187778 475210 188156
rect 473261 187776 475210 187778
rect 473261 187720 473266 187776
rect 473322 187720 475210 187776
rect 473261 187718 475210 187720
rect 500861 187778 500927 187781
rect 502014 187778 502074 188156
rect 500861 187776 502074 187778
rect 500861 187720 500866 187776
rect 500922 187720 502074 187776
rect 500861 187718 502074 187720
rect 68921 187715 68987 187718
rect 176561 187715 176627 187718
rect 284201 187715 284267 187718
rect 391841 187715 391907 187718
rect 473261 187715 473327 187718
rect 500861 187715 500927 187718
rect 64873 187506 64939 187509
rect 91093 187506 91159 187509
rect 118693 187506 118759 187509
rect 172513 187506 172579 187509
rect 200113 187506 200179 187509
rect 226333 187506 226399 187509
rect 280153 187506 280219 187509
rect 307753 187506 307819 187509
rect 335353 187506 335419 187509
rect 389173 187506 389239 187509
rect 415393 187506 415459 187509
rect 496813 187506 496879 187509
rect 523033 187506 523099 187509
rect 62836 187504 64939 187506
rect 35758 186962 35818 187476
rect 62836 187448 64878 187504
rect 64934 187448 64939 187504
rect 62836 187446 64939 187448
rect 89884 187504 91159 187506
rect 89884 187448 91098 187504
rect 91154 187448 91159 187504
rect 89884 187446 91159 187448
rect 116932 187504 118759 187506
rect 116932 187448 118698 187504
rect 118754 187448 118759 187504
rect 170844 187504 172579 187506
rect 116932 187446 118759 187448
rect 64873 187443 64939 187446
rect 91093 187443 91159 187446
rect 118693 187443 118759 187446
rect 37917 186962 37983 186965
rect 35758 186960 37983 186962
rect 35758 186904 37922 186960
rect 37978 186904 37983 186960
rect 35758 186902 37983 186904
rect 143766 186962 143826 187476
rect 170844 187448 172518 187504
rect 172574 187448 172579 187504
rect 170844 187446 172579 187448
rect 197892 187504 200179 187506
rect 197892 187448 200118 187504
rect 200174 187448 200179 187504
rect 197892 187446 200179 187448
rect 224940 187504 226399 187506
rect 224940 187448 226338 187504
rect 226394 187448 226399 187504
rect 278852 187504 280219 187506
rect 224940 187446 226399 187448
rect 172513 187443 172579 187446
rect 200113 187443 200179 187446
rect 226333 187443 226399 187446
rect 146293 186962 146359 186965
rect 143766 186960 146359 186962
rect 143766 186904 146298 186960
rect 146354 186904 146359 186960
rect 143766 186902 146359 186904
rect 251774 186962 251834 187476
rect 278852 187448 280158 187504
rect 280214 187448 280219 187504
rect 278852 187446 280219 187448
rect 305900 187504 307819 187506
rect 305900 187448 307758 187504
rect 307814 187448 307819 187504
rect 305900 187446 307819 187448
rect 332948 187504 335419 187506
rect 332948 187448 335358 187504
rect 335414 187448 335419 187504
rect 386860 187504 389239 187506
rect 332948 187446 335419 187448
rect 280153 187443 280219 187446
rect 307753 187443 307819 187446
rect 335353 187443 335419 187446
rect 253933 186962 253999 186965
rect 251774 186960 253999 186962
rect 251774 186904 253938 186960
rect 253994 186904 253999 186960
rect 251774 186902 253999 186904
rect 359782 186962 359842 187476
rect 386860 187448 389178 187504
rect 389234 187448 389239 187504
rect 386860 187446 389239 187448
rect 413908 187504 415459 187506
rect 413908 187448 415398 187504
rect 415454 187448 415459 187504
rect 494868 187504 496879 187506
rect 413908 187446 415459 187448
rect 389173 187443 389239 187446
rect 415393 187443 415459 187446
rect 361573 186962 361639 186965
rect 359782 186960 361639 186962
rect 359782 186904 361578 186960
rect 361634 186904 361639 186960
rect 359782 186902 361639 186904
rect 440926 186962 440986 187476
rect 442993 186962 443059 186965
rect 440926 186960 443059 186962
rect 440926 186904 442998 186960
rect 443054 186904 443059 186960
rect 440926 186902 443059 186904
rect 467790 186962 467850 187476
rect 494868 187448 496818 187504
rect 496874 187448 496879 187504
rect 494868 187446 496879 187448
rect 521916 187504 523099 187506
rect 521916 187448 523038 187504
rect 523094 187448 523099 187504
rect 521916 187446 523099 187448
rect 496813 187443 496879 187446
rect 523033 187443 523099 187446
rect 469213 186962 469279 186965
rect 467790 186960 469279 186962
rect 467790 186904 469218 186960
rect 469274 186904 469279 186960
rect 467790 186902 469279 186904
rect 548934 186962 548994 187476
rect 550633 186962 550699 186965
rect 548934 186960 550699 186962
rect 548934 186904 550638 186960
rect 550694 186904 550699 186960
rect 548934 186902 550699 186904
rect 37917 186899 37983 186902
rect 146293 186899 146359 186902
rect 253933 186899 253999 186902
rect 361573 186899 361639 186902
rect 442993 186899 443059 186902
rect 469213 186899 469279 186902
rect 550633 186899 550699 186902
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 526437 161394 526503 161397
rect 526437 161392 529092 161394
rect 526437 161336 526442 161392
rect 526498 161336 529092 161392
rect 526437 161334 529092 161336
rect 526437 161331 526503 161334
rect 13721 161258 13787 161261
rect 41321 161258 41387 161261
rect 95141 161258 95207 161261
rect 122741 161258 122807 161261
rect 148961 161258 149027 161261
rect 202781 161258 202847 161261
rect 230381 161258 230447 161261
rect 256601 161258 256667 161261
rect 311801 161258 311867 161261
rect 338021 161258 338087 161261
rect 365621 161258 365687 161261
rect 391841 161258 391907 161261
rect 419441 161258 419507 161261
rect 445661 161258 445727 161261
rect 500861 161258 500927 161261
rect 13721 161256 16100 161258
rect 13721 161200 13726 161256
rect 13782 161200 16100 161256
rect 13721 161198 16100 161200
rect 41321 161256 43148 161258
rect 41321 161200 41326 161256
rect 41382 161200 43148 161256
rect 95141 161256 97060 161258
rect 41321 161198 43148 161200
rect 13721 161195 13787 161198
rect 41321 161195 41387 161198
rect 68921 160714 68987 160717
rect 70166 160714 70226 161228
rect 95141 161200 95146 161256
rect 95202 161200 97060 161256
rect 95141 161198 97060 161200
rect 122741 161256 124108 161258
rect 122741 161200 122746 161256
rect 122802 161200 124108 161256
rect 122741 161198 124108 161200
rect 148961 161256 151156 161258
rect 148961 161200 148966 161256
rect 149022 161200 151156 161256
rect 202781 161256 205068 161258
rect 148961 161198 151156 161200
rect 95141 161195 95207 161198
rect 122741 161195 122807 161198
rect 148961 161195 149027 161198
rect 68921 160712 70226 160714
rect 68921 160656 68926 160712
rect 68982 160656 70226 160712
rect 68921 160654 70226 160656
rect 176561 160714 176627 160717
rect 178174 160714 178234 161228
rect 202781 161200 202786 161256
rect 202842 161200 205068 161256
rect 202781 161198 205068 161200
rect 230381 161256 232116 161258
rect 230381 161200 230386 161256
rect 230442 161200 232116 161256
rect 230381 161198 232116 161200
rect 256601 161256 259164 161258
rect 256601 161200 256606 161256
rect 256662 161200 259164 161256
rect 311801 161256 313076 161258
rect 256601 161198 259164 161200
rect 202781 161195 202847 161198
rect 230381 161195 230447 161198
rect 256601 161195 256667 161198
rect 176561 160712 178234 160714
rect 176561 160656 176566 160712
rect 176622 160656 178234 160712
rect 176561 160654 178234 160656
rect 284201 160714 284267 160717
rect 286182 160714 286242 161228
rect 311801 161200 311806 161256
rect 311862 161200 313076 161256
rect 311801 161198 313076 161200
rect 338021 161256 340124 161258
rect 338021 161200 338026 161256
rect 338082 161200 340124 161256
rect 338021 161198 340124 161200
rect 365621 161256 367172 161258
rect 365621 161200 365626 161256
rect 365682 161200 367172 161256
rect 365621 161198 367172 161200
rect 391841 161256 394036 161258
rect 391841 161200 391846 161256
rect 391902 161200 394036 161256
rect 391841 161198 394036 161200
rect 419441 161256 421084 161258
rect 419441 161200 419446 161256
rect 419502 161200 421084 161256
rect 419441 161198 421084 161200
rect 445661 161256 448132 161258
rect 445661 161200 445666 161256
rect 445722 161200 448132 161256
rect 500861 161256 502044 161258
rect 445661 161198 448132 161200
rect 311801 161195 311867 161198
rect 338021 161195 338087 161198
rect 365621 161195 365687 161198
rect 391841 161195 391907 161198
rect 419441 161195 419507 161198
rect 445661 161195 445727 161198
rect 284201 160712 286242 160714
rect 284201 160656 284206 160712
rect 284262 160656 286242 160712
rect 284201 160654 286242 160656
rect 473261 160714 473327 160717
rect 475150 160714 475210 161228
rect 500861 161200 500866 161256
rect 500922 161200 502044 161256
rect 500861 161198 502044 161200
rect 500861 161195 500927 161198
rect 473261 160712 475210 160714
rect 473261 160656 473266 160712
rect 473322 160656 475210 160712
rect 473261 160654 475210 160656
rect 68921 160651 68987 160654
rect 176561 160651 176627 160654
rect 284201 160651 284267 160654
rect 473261 160651 473327 160654
rect 64873 160578 64939 160581
rect 91093 160578 91159 160581
rect 118693 160578 118759 160581
rect 172513 160578 172579 160581
rect 200113 160578 200179 160581
rect 226333 160578 226399 160581
rect 280153 160578 280219 160581
rect 307753 160578 307819 160581
rect 335353 160578 335419 160581
rect 389173 160578 389239 160581
rect 415393 160578 415459 160581
rect 442993 160578 443059 160581
rect 496813 160578 496879 160581
rect 523033 160578 523099 160581
rect 550633 160578 550699 160581
rect 62836 160576 64939 160578
rect 35758 160170 35818 160548
rect 62836 160520 64878 160576
rect 64934 160520 64939 160576
rect 62836 160518 64939 160520
rect 89884 160576 91159 160578
rect 89884 160520 91098 160576
rect 91154 160520 91159 160576
rect 89884 160518 91159 160520
rect 116932 160576 118759 160578
rect 116932 160520 118698 160576
rect 118754 160520 118759 160576
rect 170844 160576 172579 160578
rect 116932 160518 118759 160520
rect 64873 160515 64939 160518
rect 91093 160515 91159 160518
rect 118693 160515 118759 160518
rect 37917 160170 37983 160173
rect 35758 160168 37983 160170
rect 35758 160112 37922 160168
rect 37978 160112 37983 160168
rect 35758 160110 37983 160112
rect 143766 160170 143826 160548
rect 170844 160520 172518 160576
rect 172574 160520 172579 160576
rect 170844 160518 172579 160520
rect 197892 160576 200179 160578
rect 197892 160520 200118 160576
rect 200174 160520 200179 160576
rect 197892 160518 200179 160520
rect 224940 160576 226399 160578
rect 224940 160520 226338 160576
rect 226394 160520 226399 160576
rect 278852 160576 280219 160578
rect 224940 160518 226399 160520
rect 172513 160515 172579 160518
rect 200113 160515 200179 160518
rect 226333 160515 226399 160518
rect 146293 160170 146359 160173
rect 143766 160168 146359 160170
rect 143766 160112 146298 160168
rect 146354 160112 146359 160168
rect 143766 160110 146359 160112
rect 251774 160170 251834 160548
rect 278852 160520 280158 160576
rect 280214 160520 280219 160576
rect 278852 160518 280219 160520
rect 305900 160576 307819 160578
rect 305900 160520 307758 160576
rect 307814 160520 307819 160576
rect 305900 160518 307819 160520
rect 332948 160576 335419 160578
rect 332948 160520 335358 160576
rect 335414 160520 335419 160576
rect 386860 160576 389239 160578
rect 332948 160518 335419 160520
rect 280153 160515 280219 160518
rect 307753 160515 307819 160518
rect 335353 160515 335419 160518
rect 253933 160170 253999 160173
rect 251774 160168 253999 160170
rect 251774 160112 253938 160168
rect 253994 160112 253999 160168
rect 251774 160110 253999 160112
rect 359782 160170 359842 160548
rect 386860 160520 389178 160576
rect 389234 160520 389239 160576
rect 386860 160518 389239 160520
rect 413908 160576 415459 160578
rect 413908 160520 415398 160576
rect 415454 160520 415459 160576
rect 413908 160518 415459 160520
rect 440956 160576 443059 160578
rect 440956 160520 442998 160576
rect 443054 160520 443059 160576
rect 494868 160576 496879 160578
rect 440956 160518 443059 160520
rect 389173 160515 389239 160518
rect 415393 160515 415459 160518
rect 442993 160515 443059 160518
rect 361573 160170 361639 160173
rect 359782 160168 361639 160170
rect 359782 160112 361578 160168
rect 361634 160112 361639 160168
rect 359782 160110 361639 160112
rect 467790 160170 467850 160548
rect 494868 160520 496818 160576
rect 496874 160520 496879 160576
rect 494868 160518 496879 160520
rect 521916 160576 523099 160578
rect 521916 160520 523038 160576
rect 523094 160520 523099 160576
rect 521916 160518 523099 160520
rect 548964 160576 550699 160578
rect 548964 160520 550638 160576
rect 550694 160520 550699 160576
rect 548964 160518 550699 160520
rect 496813 160515 496879 160518
rect 523033 160515 523099 160518
rect 550633 160515 550699 160518
rect 469213 160170 469279 160173
rect 467790 160168 469279 160170
rect 467790 160112 469218 160168
rect 469274 160112 469279 160168
rect 467790 160110 469279 160112
rect 37917 160107 37983 160110
rect 146293 160107 146359 160110
rect 253933 160107 253999 160110
rect 361573 160107 361639 160110
rect 469213 160107 469279 160110
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 526437 134330 526503 134333
rect 526437 134328 529092 134330
rect 526437 134272 526442 134328
rect 526498 134272 529092 134328
rect 526437 134270 529092 134272
rect 526437 134267 526503 134270
rect 13721 134194 13787 134197
rect 41321 134194 41387 134197
rect 95141 134194 95207 134197
rect 122741 134194 122807 134197
rect 148961 134194 149027 134197
rect 202781 134194 202847 134197
rect 230381 134194 230447 134197
rect 256601 134194 256667 134197
rect 311801 134194 311867 134197
rect 338021 134194 338087 134197
rect 365621 134194 365687 134197
rect 419441 134194 419507 134197
rect 445661 134194 445727 134197
rect 500861 134194 500927 134197
rect 13721 134192 16100 134194
rect 13721 134136 13726 134192
rect 13782 134136 16100 134192
rect 13721 134134 16100 134136
rect 41321 134192 43148 134194
rect 41321 134136 41326 134192
rect 41382 134136 43148 134192
rect 95141 134192 97060 134194
rect 41321 134134 43148 134136
rect 13721 134131 13787 134134
rect 41321 134131 41387 134134
rect 68921 133922 68987 133925
rect 70166 133922 70226 134164
rect 95141 134136 95146 134192
rect 95202 134136 97060 134192
rect 95141 134134 97060 134136
rect 122741 134192 124108 134194
rect 122741 134136 122746 134192
rect 122802 134136 124108 134192
rect 122741 134134 124108 134136
rect 148961 134192 151156 134194
rect 148961 134136 148966 134192
rect 149022 134136 151156 134192
rect 202781 134192 205068 134194
rect 148961 134134 151156 134136
rect 95141 134131 95207 134134
rect 122741 134131 122807 134134
rect 148961 134131 149027 134134
rect 68921 133920 70226 133922
rect 68921 133864 68926 133920
rect 68982 133864 70226 133920
rect 68921 133862 70226 133864
rect 176561 133922 176627 133925
rect 178174 133922 178234 134164
rect 202781 134136 202786 134192
rect 202842 134136 205068 134192
rect 202781 134134 205068 134136
rect 230381 134192 232116 134194
rect 230381 134136 230386 134192
rect 230442 134136 232116 134192
rect 230381 134134 232116 134136
rect 256601 134192 259164 134194
rect 256601 134136 256606 134192
rect 256662 134136 259164 134192
rect 311801 134192 313076 134194
rect 256601 134134 259164 134136
rect 202781 134131 202847 134134
rect 230381 134131 230447 134134
rect 256601 134131 256667 134134
rect 176561 133920 178234 133922
rect 176561 133864 176566 133920
rect 176622 133864 178234 133920
rect 176561 133862 178234 133864
rect 284201 133922 284267 133925
rect 286182 133922 286242 134164
rect 311801 134136 311806 134192
rect 311862 134136 313076 134192
rect 311801 134134 313076 134136
rect 338021 134192 340124 134194
rect 338021 134136 338026 134192
rect 338082 134136 340124 134192
rect 338021 134134 340124 134136
rect 365621 134192 367172 134194
rect 365621 134136 365626 134192
rect 365682 134136 367172 134192
rect 419441 134192 421084 134194
rect 365621 134134 367172 134136
rect 311801 134131 311867 134134
rect 338021 134131 338087 134134
rect 365621 134131 365687 134134
rect 284201 133920 286242 133922
rect 284201 133864 284206 133920
rect 284262 133864 286242 133920
rect 284201 133862 286242 133864
rect 391841 133922 391907 133925
rect 394006 133922 394066 134164
rect 419441 134136 419446 134192
rect 419502 134136 421084 134192
rect 419441 134134 421084 134136
rect 445661 134192 448132 134194
rect 445661 134136 445666 134192
rect 445722 134136 448132 134192
rect 500861 134192 502044 134194
rect 445661 134134 448132 134136
rect 419441 134131 419507 134134
rect 445661 134131 445727 134134
rect 391841 133920 394066 133922
rect 391841 133864 391846 133920
rect 391902 133864 394066 133920
rect 391841 133862 394066 133864
rect 473261 133922 473327 133925
rect 475150 133922 475210 134164
rect 500861 134136 500866 134192
rect 500922 134136 502044 134192
rect 500861 134134 502044 134136
rect 500861 134131 500927 134134
rect 473261 133920 475210 133922
rect 473261 133864 473266 133920
rect 473322 133864 475210 133920
rect 473261 133862 475210 133864
rect 68921 133859 68987 133862
rect 176561 133859 176627 133862
rect 284201 133859 284267 133862
rect 391841 133859 391907 133862
rect 473261 133859 473327 133862
rect 64873 133514 64939 133517
rect 91093 133514 91159 133517
rect 118693 133514 118759 133517
rect 172513 133514 172579 133517
rect 200113 133514 200179 133517
rect 226333 133514 226399 133517
rect 280153 133514 280219 133517
rect 307753 133514 307819 133517
rect 335353 133514 335419 133517
rect 389173 133514 389239 133517
rect 415393 133514 415459 133517
rect 442993 133514 443059 133517
rect 496813 133514 496879 133517
rect 523033 133514 523099 133517
rect 62836 133512 64939 133514
rect 35758 132970 35818 133484
rect 62836 133456 64878 133512
rect 64934 133456 64939 133512
rect 62836 133454 64939 133456
rect 89884 133512 91159 133514
rect 89884 133456 91098 133512
rect 91154 133456 91159 133512
rect 89884 133454 91159 133456
rect 116932 133512 118759 133514
rect 116932 133456 118698 133512
rect 118754 133456 118759 133512
rect 170844 133512 172579 133514
rect 116932 133454 118759 133456
rect 64873 133451 64939 133454
rect 91093 133451 91159 133454
rect 118693 133451 118759 133454
rect 37917 132970 37983 132973
rect 35758 132968 37983 132970
rect 35758 132912 37922 132968
rect 37978 132912 37983 132968
rect 35758 132910 37983 132912
rect 143766 132970 143826 133484
rect 170844 133456 172518 133512
rect 172574 133456 172579 133512
rect 170844 133454 172579 133456
rect 197892 133512 200179 133514
rect 197892 133456 200118 133512
rect 200174 133456 200179 133512
rect 197892 133454 200179 133456
rect 224940 133512 226399 133514
rect 224940 133456 226338 133512
rect 226394 133456 226399 133512
rect 278852 133512 280219 133514
rect 224940 133454 226399 133456
rect 172513 133451 172579 133454
rect 200113 133451 200179 133454
rect 226333 133451 226399 133454
rect 146293 132970 146359 132973
rect 143766 132968 146359 132970
rect 143766 132912 146298 132968
rect 146354 132912 146359 132968
rect 143766 132910 146359 132912
rect 251774 132970 251834 133484
rect 278852 133456 280158 133512
rect 280214 133456 280219 133512
rect 278852 133454 280219 133456
rect 305900 133512 307819 133514
rect 305900 133456 307758 133512
rect 307814 133456 307819 133512
rect 305900 133454 307819 133456
rect 332948 133512 335419 133514
rect 332948 133456 335358 133512
rect 335414 133456 335419 133512
rect 386860 133512 389239 133514
rect 332948 133454 335419 133456
rect 280153 133451 280219 133454
rect 307753 133451 307819 133454
rect 335353 133451 335419 133454
rect 253933 132970 253999 132973
rect 251774 132968 253999 132970
rect 251774 132912 253938 132968
rect 253994 132912 253999 132968
rect 251774 132910 253999 132912
rect 359782 132970 359842 133484
rect 386860 133456 389178 133512
rect 389234 133456 389239 133512
rect 386860 133454 389239 133456
rect 413908 133512 415459 133514
rect 413908 133456 415398 133512
rect 415454 133456 415459 133512
rect 413908 133454 415459 133456
rect 440956 133512 443059 133514
rect 440956 133456 442998 133512
rect 443054 133456 443059 133512
rect 494868 133512 496879 133514
rect 440956 133454 443059 133456
rect 389173 133451 389239 133454
rect 415393 133451 415459 133454
rect 442993 133451 443059 133454
rect 361573 132970 361639 132973
rect 359782 132968 361639 132970
rect 359782 132912 361578 132968
rect 361634 132912 361639 132968
rect 359782 132910 361639 132912
rect 467790 132970 467850 133484
rect 494868 133456 496818 133512
rect 496874 133456 496879 133512
rect 494868 133454 496879 133456
rect 521916 133512 523099 133514
rect 521916 133456 523038 133512
rect 523094 133456 523099 133512
rect 521916 133454 523099 133456
rect 496813 133451 496879 133454
rect 523033 133451 523099 133454
rect 469213 132970 469279 132973
rect 467790 132968 469279 132970
rect 467790 132912 469218 132968
rect 469274 132912 469279 132968
rect 467790 132910 469279 132912
rect 548934 132970 548994 133484
rect 550633 132970 550699 132973
rect 548934 132968 550699 132970
rect 548934 132912 550638 132968
rect 550694 132912 550699 132968
rect 548934 132910 550699 132912
rect 37917 132907 37983 132910
rect 146293 132907 146359 132910
rect 253933 132907 253999 132910
rect 361573 132907 361639 132910
rect 469213 132907 469279 132910
rect 550633 132907 550699 132910
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 526437 107402 526503 107405
rect 526437 107400 529092 107402
rect 526437 107344 526442 107400
rect 526498 107344 529092 107400
rect 526437 107342 529092 107344
rect 526437 107339 526503 107342
rect 13721 107266 13787 107269
rect 41321 107266 41387 107269
rect 95141 107266 95207 107269
rect 122741 107266 122807 107269
rect 148961 107266 149027 107269
rect 202781 107266 202847 107269
rect 230381 107266 230447 107269
rect 256601 107266 256667 107269
rect 311801 107266 311867 107269
rect 338021 107266 338087 107269
rect 365621 107266 365687 107269
rect 391841 107266 391907 107269
rect 419441 107266 419507 107269
rect 445661 107266 445727 107269
rect 500861 107266 500927 107269
rect 13721 107264 16100 107266
rect 13721 107208 13726 107264
rect 13782 107208 16100 107264
rect 13721 107206 16100 107208
rect 41321 107264 43148 107266
rect 41321 107208 41326 107264
rect 41382 107208 43148 107264
rect 95141 107264 97060 107266
rect 41321 107206 43148 107208
rect 13721 107203 13787 107206
rect 41321 107203 41387 107206
rect 68921 106722 68987 106725
rect 70166 106722 70226 107236
rect 95141 107208 95146 107264
rect 95202 107208 97060 107264
rect 95141 107206 97060 107208
rect 122741 107264 124108 107266
rect 122741 107208 122746 107264
rect 122802 107208 124108 107264
rect 122741 107206 124108 107208
rect 148961 107264 151156 107266
rect 148961 107208 148966 107264
rect 149022 107208 151156 107264
rect 202781 107264 205068 107266
rect 148961 107206 151156 107208
rect 95141 107203 95207 107206
rect 122741 107203 122807 107206
rect 148961 107203 149027 107206
rect 68921 106720 70226 106722
rect 68921 106664 68926 106720
rect 68982 106664 70226 106720
rect 68921 106662 70226 106664
rect 176561 106722 176627 106725
rect 178174 106722 178234 107236
rect 202781 107208 202786 107264
rect 202842 107208 205068 107264
rect 202781 107206 205068 107208
rect 230381 107264 232116 107266
rect 230381 107208 230386 107264
rect 230442 107208 232116 107264
rect 230381 107206 232116 107208
rect 256601 107264 259164 107266
rect 256601 107208 256606 107264
rect 256662 107208 259164 107264
rect 311801 107264 313076 107266
rect 256601 107206 259164 107208
rect 202781 107203 202847 107206
rect 230381 107203 230447 107206
rect 256601 107203 256667 107206
rect 176561 106720 178234 106722
rect 176561 106664 176566 106720
rect 176622 106664 178234 106720
rect 176561 106662 178234 106664
rect 284201 106722 284267 106725
rect 286182 106722 286242 107236
rect 311801 107208 311806 107264
rect 311862 107208 313076 107264
rect 311801 107206 313076 107208
rect 338021 107264 340124 107266
rect 338021 107208 338026 107264
rect 338082 107208 340124 107264
rect 338021 107206 340124 107208
rect 365621 107264 367172 107266
rect 365621 107208 365626 107264
rect 365682 107208 367172 107264
rect 365621 107206 367172 107208
rect 391841 107264 394036 107266
rect 391841 107208 391846 107264
rect 391902 107208 394036 107264
rect 391841 107206 394036 107208
rect 419441 107264 421084 107266
rect 419441 107208 419446 107264
rect 419502 107208 421084 107264
rect 419441 107206 421084 107208
rect 445661 107264 448132 107266
rect 445661 107208 445666 107264
rect 445722 107208 448132 107264
rect 500861 107264 502044 107266
rect 445661 107206 448132 107208
rect 311801 107203 311867 107206
rect 338021 107203 338087 107206
rect 365621 107203 365687 107206
rect 391841 107203 391907 107206
rect 419441 107203 419507 107206
rect 445661 107203 445727 107206
rect 284201 106720 286242 106722
rect 284201 106664 284206 106720
rect 284262 106664 286242 106720
rect 284201 106662 286242 106664
rect 473261 106722 473327 106725
rect 475150 106722 475210 107236
rect 500861 107208 500866 107264
rect 500922 107208 502044 107264
rect 500861 107206 502044 107208
rect 500861 107203 500927 107206
rect 473261 106720 475210 106722
rect 473261 106664 473266 106720
rect 473322 106664 475210 106720
rect 473261 106662 475210 106664
rect 68921 106659 68987 106662
rect 176561 106659 176627 106662
rect 284201 106659 284267 106662
rect 473261 106659 473327 106662
rect 37917 106586 37983 106589
rect 64873 106586 64939 106589
rect 91093 106586 91159 106589
rect 118693 106586 118759 106589
rect 172513 106586 172579 106589
rect 200113 106586 200179 106589
rect 226333 106586 226399 106589
rect 280153 106586 280219 106589
rect 307753 106586 307819 106589
rect 335353 106586 335419 106589
rect 389173 106586 389239 106589
rect 415393 106586 415459 106589
rect 442993 106586 443059 106589
rect 496813 106586 496879 106589
rect 523033 106586 523099 106589
rect 550633 106586 550699 106589
rect 35850 106584 37983 106586
rect 35574 106314 35634 106556
rect 35850 106528 37922 106584
rect 37978 106528 37983 106584
rect 35850 106526 37983 106528
rect 62836 106584 64939 106586
rect 62836 106528 64878 106584
rect 64934 106528 64939 106584
rect 62836 106526 64939 106528
rect 89884 106584 91159 106586
rect 89884 106528 91098 106584
rect 91154 106528 91159 106584
rect 89884 106526 91159 106528
rect 116932 106584 118759 106586
rect 116932 106528 118698 106584
rect 118754 106528 118759 106584
rect 170844 106584 172579 106586
rect 116932 106526 118759 106528
rect 35850 106314 35910 106526
rect 37917 106523 37983 106526
rect 64873 106523 64939 106526
rect 91093 106523 91159 106526
rect 118693 106523 118759 106526
rect 35574 106254 35910 106314
rect 143766 106314 143826 106556
rect 170844 106528 172518 106584
rect 172574 106528 172579 106584
rect 170844 106526 172579 106528
rect 197892 106584 200179 106586
rect 197892 106528 200118 106584
rect 200174 106528 200179 106584
rect 197892 106526 200179 106528
rect 224940 106584 226399 106586
rect 224940 106528 226338 106584
rect 226394 106528 226399 106584
rect 278852 106584 280219 106586
rect 224940 106526 226399 106528
rect 172513 106523 172579 106526
rect 200113 106523 200179 106526
rect 226333 106523 226399 106526
rect 146293 106314 146359 106317
rect 143766 106312 146359 106314
rect 143766 106256 146298 106312
rect 146354 106256 146359 106312
rect 143766 106254 146359 106256
rect 251774 106314 251834 106556
rect 278852 106528 280158 106584
rect 280214 106528 280219 106584
rect 278852 106526 280219 106528
rect 305900 106584 307819 106586
rect 305900 106528 307758 106584
rect 307814 106528 307819 106584
rect 305900 106526 307819 106528
rect 332948 106584 335419 106586
rect 332948 106528 335358 106584
rect 335414 106528 335419 106584
rect 386860 106584 389239 106586
rect 332948 106526 335419 106528
rect 280153 106523 280219 106526
rect 307753 106523 307819 106526
rect 335353 106523 335419 106526
rect 253933 106314 253999 106317
rect 251774 106312 253999 106314
rect 251774 106256 253938 106312
rect 253994 106256 253999 106312
rect 251774 106254 253999 106256
rect 359782 106314 359842 106556
rect 386860 106528 389178 106584
rect 389234 106528 389239 106584
rect 386860 106526 389239 106528
rect 413908 106584 415459 106586
rect 413908 106528 415398 106584
rect 415454 106528 415459 106584
rect 413908 106526 415459 106528
rect 440956 106584 443059 106586
rect 440956 106528 442998 106584
rect 443054 106528 443059 106584
rect 494868 106584 496879 106586
rect 440956 106526 443059 106528
rect 389173 106523 389239 106526
rect 415393 106523 415459 106526
rect 442993 106523 443059 106526
rect 361573 106314 361639 106317
rect 359782 106312 361639 106314
rect 359782 106256 361578 106312
rect 361634 106256 361639 106312
rect 359782 106254 361639 106256
rect 467790 106314 467850 106556
rect 494868 106528 496818 106584
rect 496874 106528 496879 106584
rect 494868 106526 496879 106528
rect 521916 106584 523099 106586
rect 521916 106528 523038 106584
rect 523094 106528 523099 106584
rect 521916 106526 523099 106528
rect 548964 106584 550699 106586
rect 548964 106528 550638 106584
rect 550694 106528 550699 106584
rect 548964 106526 550699 106528
rect 496813 106523 496879 106526
rect 523033 106523 523099 106526
rect 550633 106523 550699 106526
rect 469213 106314 469279 106317
rect 467790 106312 469279 106314
rect 467790 106256 469218 106312
rect 469274 106256 469279 106312
rect 467790 106254 469279 106256
rect 146293 106251 146359 106254
rect 253933 106251 253999 106254
rect 361573 106251 361639 106254
rect 469213 106251 469279 106254
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 68921 80882 68987 80885
rect 176561 80882 176627 80885
rect 284201 80882 284267 80885
rect 473261 80882 473327 80885
rect 68921 80880 70226 80882
rect 68921 80824 68926 80880
rect 68982 80824 70226 80880
rect 68921 80822 70226 80824
rect 68921 80819 68987 80822
rect 13721 80338 13787 80341
rect 41321 80338 41387 80341
rect 13721 80336 16100 80338
rect 13721 80280 13726 80336
rect 13782 80280 16100 80336
rect 13721 80278 16100 80280
rect 41321 80336 43148 80338
rect 41321 80280 41326 80336
rect 41382 80280 43148 80336
rect 70166 80308 70226 80822
rect 176561 80880 178234 80882
rect 176561 80824 176566 80880
rect 176622 80824 178234 80880
rect 176561 80822 178234 80824
rect 176561 80819 176627 80822
rect 95141 80338 95207 80341
rect 122741 80338 122807 80341
rect 148961 80338 149027 80341
rect 95141 80336 97060 80338
rect 41321 80278 43148 80280
rect 95141 80280 95146 80336
rect 95202 80280 97060 80336
rect 95141 80278 97060 80280
rect 122741 80336 124108 80338
rect 122741 80280 122746 80336
rect 122802 80280 124108 80336
rect 122741 80278 124108 80280
rect 148961 80336 151156 80338
rect 148961 80280 148966 80336
rect 149022 80280 151156 80336
rect 178174 80308 178234 80822
rect 284201 80880 286242 80882
rect 284201 80824 284206 80880
rect 284262 80824 286242 80880
rect 284201 80822 286242 80824
rect 284201 80819 284267 80822
rect 202781 80338 202847 80341
rect 230381 80338 230447 80341
rect 256601 80338 256667 80341
rect 202781 80336 205068 80338
rect 148961 80278 151156 80280
rect 202781 80280 202786 80336
rect 202842 80280 205068 80336
rect 202781 80278 205068 80280
rect 230381 80336 232116 80338
rect 230381 80280 230386 80336
rect 230442 80280 232116 80336
rect 230381 80278 232116 80280
rect 256601 80336 259164 80338
rect 256601 80280 256606 80336
rect 256662 80280 259164 80336
rect 286182 80308 286242 80822
rect 473261 80880 475210 80882
rect 473261 80824 473266 80880
rect 473322 80824 475210 80880
rect 473261 80822 475210 80824
rect 473261 80819 473327 80822
rect 311801 80338 311867 80341
rect 338021 80338 338087 80341
rect 365621 80338 365687 80341
rect 391841 80338 391907 80341
rect 419441 80338 419507 80341
rect 445661 80338 445727 80341
rect 311801 80336 313076 80338
rect 256601 80278 259164 80280
rect 311801 80280 311806 80336
rect 311862 80280 313076 80336
rect 311801 80278 313076 80280
rect 338021 80336 340124 80338
rect 338021 80280 338026 80336
rect 338082 80280 340124 80336
rect 338021 80278 340124 80280
rect 365621 80336 367172 80338
rect 365621 80280 365626 80336
rect 365682 80280 367172 80336
rect 365621 80278 367172 80280
rect 391841 80336 394036 80338
rect 391841 80280 391846 80336
rect 391902 80280 394036 80336
rect 391841 80278 394036 80280
rect 419441 80336 421084 80338
rect 419441 80280 419446 80336
rect 419502 80280 421084 80336
rect 419441 80278 421084 80280
rect 445661 80336 448132 80338
rect 445661 80280 445666 80336
rect 445722 80280 448132 80336
rect 475150 80308 475210 80822
rect 500861 80338 500927 80341
rect 526437 80338 526503 80341
rect 500861 80336 502044 80338
rect 445661 80278 448132 80280
rect 500861 80280 500866 80336
rect 500922 80280 502044 80336
rect 500861 80278 502044 80280
rect 526437 80336 529092 80338
rect 526437 80280 526442 80336
rect 526498 80280 529092 80336
rect 526437 80278 529092 80280
rect 13721 80275 13787 80278
rect 41321 80275 41387 80278
rect 95141 80275 95207 80278
rect 122741 80275 122807 80278
rect 148961 80275 149027 80278
rect 202781 80275 202847 80278
rect 230381 80275 230447 80278
rect 256601 80275 256667 80278
rect 311801 80275 311867 80278
rect 338021 80275 338087 80278
rect 365621 80275 365687 80278
rect 391841 80275 391907 80278
rect 419441 80275 419507 80278
rect 445661 80275 445727 80278
rect 500861 80275 500927 80278
rect 526437 80275 526503 80278
rect 146293 80066 146359 80069
rect 253933 80066 253999 80069
rect 361573 80066 361639 80069
rect 469213 80066 469279 80069
rect 143766 80064 146359 80066
rect 143766 80008 146298 80064
rect 146354 80008 146359 80064
rect 143766 80006 146359 80008
rect 64873 79658 64939 79661
rect 91093 79658 91159 79661
rect 118693 79658 118759 79661
rect 62836 79656 64939 79658
rect 62836 79600 64878 79656
rect 64934 79600 64939 79656
rect 62836 79598 64939 79600
rect 89884 79656 91159 79658
rect 89884 79600 91098 79656
rect 91154 79600 91159 79656
rect 89884 79598 91159 79600
rect 116932 79656 118759 79658
rect 116932 79600 118698 79656
rect 118754 79600 118759 79656
rect 143766 79628 143826 80006
rect 146293 80003 146359 80006
rect 251774 80064 253999 80066
rect 251774 80008 253938 80064
rect 253994 80008 253999 80064
rect 251774 80006 253999 80008
rect 172513 79658 172579 79661
rect 200113 79658 200179 79661
rect 226333 79658 226399 79661
rect 170844 79656 172579 79658
rect 116932 79598 118759 79600
rect 170844 79600 172518 79656
rect 172574 79600 172579 79656
rect 170844 79598 172579 79600
rect 197892 79656 200179 79658
rect 197892 79600 200118 79656
rect 200174 79600 200179 79656
rect 197892 79598 200179 79600
rect 224940 79656 226399 79658
rect 224940 79600 226338 79656
rect 226394 79600 226399 79656
rect 251774 79628 251834 80006
rect 253933 80003 253999 80006
rect 359782 80064 361639 80066
rect 359782 80008 361578 80064
rect 361634 80008 361639 80064
rect 359782 80006 361639 80008
rect 280153 79658 280219 79661
rect 307753 79658 307819 79661
rect 335353 79658 335419 79661
rect 278852 79656 280219 79658
rect 224940 79598 226399 79600
rect 278852 79600 280158 79656
rect 280214 79600 280219 79656
rect 278852 79598 280219 79600
rect 305900 79656 307819 79658
rect 305900 79600 307758 79656
rect 307814 79600 307819 79656
rect 305900 79598 307819 79600
rect 332948 79656 335419 79658
rect 332948 79600 335358 79656
rect 335414 79600 335419 79656
rect 359782 79628 359842 80006
rect 361573 80003 361639 80006
rect 467790 80064 469279 80066
rect 467790 80008 469218 80064
rect 469274 80008 469279 80064
rect 467790 80006 469279 80008
rect 389173 79658 389239 79661
rect 415393 79658 415459 79661
rect 442993 79658 443059 79661
rect 386860 79656 389239 79658
rect 332948 79598 335419 79600
rect 386860 79600 389178 79656
rect 389234 79600 389239 79656
rect 386860 79598 389239 79600
rect 413908 79656 415459 79658
rect 413908 79600 415398 79656
rect 415454 79600 415459 79656
rect 413908 79598 415459 79600
rect 440956 79656 443059 79658
rect 440956 79600 442998 79656
rect 443054 79600 443059 79656
rect 467790 79628 467850 80006
rect 469213 80003 469279 80006
rect 496813 79658 496879 79661
rect 523033 79658 523099 79661
rect 550633 79658 550699 79661
rect 494868 79656 496879 79658
rect 440956 79598 443059 79600
rect 494868 79600 496818 79656
rect 496874 79600 496879 79656
rect 494868 79598 496879 79600
rect 521916 79656 523099 79658
rect 521916 79600 523038 79656
rect 523094 79600 523099 79656
rect 521916 79598 523099 79600
rect 548964 79656 550699 79658
rect 548964 79600 550638 79656
rect 550694 79600 550699 79656
rect 548964 79598 550699 79600
rect 64873 79595 64939 79598
rect 91093 79595 91159 79598
rect 118693 79595 118759 79598
rect 172513 79595 172579 79598
rect 200113 79595 200179 79598
rect 226333 79595 226399 79598
rect 280153 79595 280219 79598
rect 307753 79595 307819 79598
rect 335353 79595 335419 79598
rect 389173 79595 389239 79598
rect 415393 79595 415459 79598
rect 442993 79595 443059 79598
rect 496813 79595 496879 79598
rect 523033 79595 523099 79598
rect 550633 79595 550699 79598
rect 35758 78978 35818 79492
rect 37917 78978 37983 78981
rect 35758 78976 37983 78978
rect 35758 78920 37922 78976
rect 37978 78920 37983 78976
rect 35758 78918 37983 78920
rect 37917 78915 37983 78918
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 68921 53818 68987 53821
rect 284201 53818 284267 53821
rect 473261 53818 473327 53821
rect 500861 53818 500927 53821
rect 68921 53816 70226 53818
rect 68921 53760 68926 53816
rect 68982 53760 70226 53816
rect 68921 53758 70226 53760
rect 68921 53755 68987 53758
rect 41321 53410 41387 53413
rect 41321 53408 43148 53410
rect 41321 53352 41326 53408
rect 41382 53352 43148 53408
rect 70166 53380 70226 53758
rect 284201 53816 286242 53818
rect 284201 53760 284206 53816
rect 284262 53760 286242 53816
rect 284201 53758 286242 53760
rect 284201 53755 284267 53758
rect 122741 53410 122807 53413
rect 148961 53410 149027 53413
rect 202781 53410 202847 53413
rect 230381 53410 230447 53413
rect 122741 53408 124108 53410
rect 41321 53350 43148 53352
rect 122741 53352 122746 53408
rect 122802 53352 124108 53408
rect 122741 53350 124108 53352
rect 148961 53408 151156 53410
rect 148961 53352 148966 53408
rect 149022 53352 151156 53408
rect 148961 53350 151156 53352
rect 202781 53408 205068 53410
rect 202781 53352 202786 53408
rect 202842 53352 205068 53408
rect 202781 53350 205068 53352
rect 230381 53408 232116 53410
rect 230381 53352 230386 53408
rect 230442 53352 232116 53408
rect 286182 53380 286242 53758
rect 473261 53816 475210 53818
rect 473261 53760 473266 53816
rect 473322 53760 475210 53816
rect 473261 53758 475210 53760
rect 473261 53755 473327 53758
rect 311801 53410 311867 53413
rect 365621 53410 365687 53413
rect 419441 53410 419507 53413
rect 311801 53408 313076 53410
rect 230381 53350 232116 53352
rect 311801 53352 311806 53408
rect 311862 53352 313076 53408
rect 311801 53350 313076 53352
rect 365621 53408 367172 53410
rect 365621 53352 365626 53408
rect 365682 53352 367172 53408
rect 365621 53350 367172 53352
rect 419441 53408 421084 53410
rect 419441 53352 419446 53408
rect 419502 53352 421084 53408
rect 475150 53380 475210 53758
rect 500861 53816 502074 53818
rect 500861 53760 500866 53816
rect 500922 53760 502074 53816
rect 500861 53758 502074 53760
rect 500861 53755 500927 53758
rect 502014 53380 502074 53758
rect 526437 53410 526503 53413
rect 526437 53408 529092 53410
rect 419441 53350 421084 53352
rect 526437 53352 526442 53408
rect 526498 53352 529092 53408
rect 526437 53350 529092 53352
rect 41321 53347 41387 53350
rect 122741 53347 122807 53350
rect 148961 53347 149027 53350
rect 202781 53347 202847 53350
rect 230381 53347 230447 53350
rect 311801 53347 311867 53350
rect 365621 53347 365687 53350
rect 419441 53347 419507 53350
rect 526437 53347 526503 53350
rect 13721 53274 13787 53277
rect 95141 53274 95207 53277
rect 253933 53274 253999 53277
rect 13721 53272 16100 53274
rect 13721 53216 13726 53272
rect 13782 53216 16100 53272
rect 13721 53214 16100 53216
rect 95141 53272 97060 53274
rect 95141 53216 95146 53272
rect 95202 53216 97060 53272
rect 251774 53272 253999 53274
rect 95141 53214 97060 53216
rect 13721 53211 13787 53214
rect 95141 53211 95207 53214
rect 37917 52866 37983 52869
rect 146293 52866 146359 52869
rect 35758 52864 37983 52866
rect 35758 52808 37922 52864
rect 37978 52808 37983 52864
rect 35758 52806 37983 52808
rect 35758 52700 35818 52806
rect 37917 52803 37983 52806
rect 143766 52864 146359 52866
rect 143766 52808 146298 52864
rect 146354 52808 146359 52864
rect 143766 52806 146359 52808
rect 91093 52730 91159 52733
rect 118693 52730 118759 52733
rect 89884 52728 91159 52730
rect 89884 52672 91098 52728
rect 91154 52672 91159 52728
rect 89884 52670 91159 52672
rect 116932 52728 118759 52730
rect 116932 52672 118698 52728
rect 118754 52672 118759 52728
rect 143766 52700 143826 52806
rect 146293 52803 146359 52806
rect 172513 52730 172579 52733
rect 170844 52728 172579 52730
rect 116932 52670 118759 52672
rect 170844 52672 172518 52728
rect 172574 52672 172579 52728
rect 170844 52670 172579 52672
rect 91093 52667 91159 52670
rect 118693 52667 118759 52670
rect 172513 52667 172579 52670
rect 176561 52730 176627 52733
rect 178174 52730 178234 53244
rect 251774 53216 253938 53272
rect 253994 53216 253999 53272
rect 251774 53214 253999 53216
rect 200113 52730 200179 52733
rect 176561 52728 178234 52730
rect 176561 52672 176566 52728
rect 176622 52672 178234 52728
rect 176561 52670 178234 52672
rect 197892 52728 200179 52730
rect 197892 52672 200118 52728
rect 200174 52672 200179 52728
rect 251774 52700 251834 53214
rect 253933 53211 253999 53214
rect 256601 53274 256667 53277
rect 338021 53274 338087 53277
rect 361573 53274 361639 53277
rect 256601 53272 259164 53274
rect 256601 53216 256606 53272
rect 256662 53216 259164 53272
rect 256601 53214 259164 53216
rect 338021 53272 340124 53274
rect 338021 53216 338026 53272
rect 338082 53216 340124 53272
rect 338021 53214 340124 53216
rect 359782 53272 361639 53274
rect 359782 53216 361578 53272
rect 361634 53216 361639 53272
rect 359782 53214 361639 53216
rect 256601 53211 256667 53214
rect 338021 53211 338087 53214
rect 280153 52730 280219 52733
rect 335353 52730 335419 52733
rect 278852 52728 280219 52730
rect 197892 52670 200179 52672
rect 278852 52672 280158 52728
rect 280214 52672 280219 52728
rect 278852 52670 280219 52672
rect 332948 52728 335419 52730
rect 332948 52672 335358 52728
rect 335414 52672 335419 52728
rect 359782 52700 359842 53214
rect 361573 53211 361639 53214
rect 391841 53274 391907 53277
rect 445661 53274 445727 53277
rect 469213 53274 469279 53277
rect 550633 53274 550699 53277
rect 391841 53272 394036 53274
rect 391841 53216 391846 53272
rect 391902 53216 394036 53272
rect 391841 53214 394036 53216
rect 445661 53272 448132 53274
rect 445661 53216 445666 53272
rect 445722 53216 448132 53272
rect 445661 53214 448132 53216
rect 467790 53272 469279 53274
rect 467790 53216 469218 53272
rect 469274 53216 469279 53272
rect 467790 53214 469279 53216
rect 391841 53211 391907 53214
rect 445661 53211 445727 53214
rect 415393 52730 415459 52733
rect 413908 52728 415459 52730
rect 332948 52670 335419 52672
rect 413908 52672 415398 52728
rect 415454 52672 415459 52728
rect 467790 52700 467850 53214
rect 469213 53211 469279 53214
rect 548934 53272 550699 53274
rect 548934 53216 550638 53272
rect 550694 53216 550699 53272
rect 548934 53214 550699 53216
rect 523033 52730 523099 52733
rect 521916 52728 523099 52730
rect 413908 52670 415459 52672
rect 521916 52672 523038 52728
rect 523094 52672 523099 52728
rect 548934 52700 548994 53214
rect 550633 53211 550699 53214
rect 521916 52670 523099 52672
rect 176561 52667 176627 52670
rect 200113 52667 200179 52670
rect 280153 52667 280219 52670
rect 335353 52667 335419 52670
rect 415393 52667 415459 52670
rect 523033 52667 523099 52670
rect 64873 52594 64939 52597
rect 226333 52594 226399 52597
rect 307753 52594 307819 52597
rect 389173 52594 389239 52597
rect 442993 52594 443059 52597
rect 496813 52594 496879 52597
rect 62836 52592 64939 52594
rect 62836 52536 64878 52592
rect 64934 52536 64939 52592
rect 62836 52534 64939 52536
rect 224940 52592 226399 52594
rect 224940 52536 226338 52592
rect 226394 52536 226399 52592
rect 224940 52534 226399 52536
rect 305900 52592 307819 52594
rect 305900 52536 307758 52592
rect 307814 52536 307819 52592
rect 305900 52534 307819 52536
rect 386860 52592 389239 52594
rect 386860 52536 389178 52592
rect 389234 52536 389239 52592
rect 386860 52534 389239 52536
rect 440956 52592 443059 52594
rect 440956 52536 442998 52592
rect 443054 52536 443059 52592
rect 440956 52534 443059 52536
rect 494868 52592 496879 52594
rect 494868 52536 496818 52592
rect 496874 52536 496879 52592
rect 494868 52534 496879 52536
rect 64873 52531 64939 52534
rect 226333 52531 226399 52534
rect 307753 52531 307819 52534
rect 389173 52531 389239 52534
rect 442993 52531 443059 52534
rect 496813 52531 496879 52534
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 68921 26890 68987 26893
rect 176561 26890 176627 26893
rect 284201 26890 284267 26893
rect 473261 26890 473327 26893
rect 68921 26888 70226 26890
rect 68921 26832 68926 26888
rect 68982 26832 70226 26888
rect 68921 26830 70226 26832
rect 68921 26827 68987 26830
rect 13721 26346 13787 26349
rect 41321 26346 41387 26349
rect 13721 26344 16100 26346
rect 13721 26288 13726 26344
rect 13782 26288 16100 26344
rect 13721 26286 16100 26288
rect 41321 26344 43148 26346
rect 41321 26288 41326 26344
rect 41382 26288 43148 26344
rect 70166 26316 70226 26830
rect 176561 26888 178234 26890
rect 176561 26832 176566 26888
rect 176622 26832 178234 26888
rect 176561 26830 178234 26832
rect 176561 26827 176627 26830
rect 95141 26346 95207 26349
rect 122741 26346 122807 26349
rect 148961 26346 149027 26349
rect 95141 26344 97060 26346
rect 41321 26286 43148 26288
rect 95141 26288 95146 26344
rect 95202 26288 97060 26344
rect 95141 26286 97060 26288
rect 122741 26344 124108 26346
rect 122741 26288 122746 26344
rect 122802 26288 124108 26344
rect 122741 26286 124108 26288
rect 148961 26344 151156 26346
rect 148961 26288 148966 26344
rect 149022 26288 151156 26344
rect 178174 26316 178234 26830
rect 284201 26888 286242 26890
rect 284201 26832 284206 26888
rect 284262 26832 286242 26888
rect 284201 26830 286242 26832
rect 284201 26827 284267 26830
rect 202781 26346 202847 26349
rect 230381 26346 230447 26349
rect 256601 26346 256667 26349
rect 202781 26344 205068 26346
rect 148961 26286 151156 26288
rect 202781 26288 202786 26344
rect 202842 26288 205068 26344
rect 202781 26286 205068 26288
rect 230381 26344 232116 26346
rect 230381 26288 230386 26344
rect 230442 26288 232116 26344
rect 230381 26286 232116 26288
rect 256601 26344 259164 26346
rect 256601 26288 256606 26344
rect 256662 26288 259164 26344
rect 286182 26316 286242 26830
rect 473261 26888 475210 26890
rect 473261 26832 473266 26888
rect 473322 26832 475210 26888
rect 473261 26830 475210 26832
rect 473261 26827 473327 26830
rect 311801 26346 311867 26349
rect 338021 26346 338087 26349
rect 365621 26346 365687 26349
rect 391841 26346 391907 26349
rect 419441 26346 419507 26349
rect 445661 26346 445727 26349
rect 311801 26344 313076 26346
rect 256601 26286 259164 26288
rect 311801 26288 311806 26344
rect 311862 26288 313076 26344
rect 311801 26286 313076 26288
rect 338021 26344 340124 26346
rect 338021 26288 338026 26344
rect 338082 26288 340124 26344
rect 338021 26286 340124 26288
rect 365621 26344 367070 26346
rect 365621 26288 365626 26344
rect 365682 26288 367070 26344
rect 365621 26286 367070 26288
rect 13721 26283 13787 26286
rect 41321 26283 41387 26286
rect 95141 26283 95207 26286
rect 122741 26283 122807 26286
rect 148961 26283 149027 26286
rect 202781 26283 202847 26286
rect 230381 26283 230447 26286
rect 256601 26283 256667 26286
rect 311801 26283 311867 26286
rect 338021 26283 338087 26286
rect 365621 26283 365687 26286
rect 38009 26210 38075 26213
rect 35758 26208 38075 26210
rect 35758 26152 38014 26208
rect 38070 26152 38075 26208
rect 35758 26150 38075 26152
rect 367010 26210 367070 26286
rect 391841 26344 394036 26346
rect 391841 26288 391846 26344
rect 391902 26288 394036 26344
rect 391841 26286 394036 26288
rect 419441 26344 421084 26346
rect 419441 26288 419446 26344
rect 419502 26288 421084 26344
rect 419441 26286 421084 26288
rect 445661 26344 448132 26346
rect 445661 26288 445666 26344
rect 445722 26288 448132 26344
rect 475150 26316 475210 26830
rect 500861 26346 500927 26349
rect 526437 26346 526503 26349
rect 500861 26344 502044 26346
rect 445661 26286 448132 26288
rect 500861 26288 500866 26344
rect 500922 26288 502044 26344
rect 500861 26286 502044 26288
rect 526437 26344 529092 26346
rect 526437 26288 526442 26344
rect 526498 26288 529092 26344
rect 526437 26286 529092 26288
rect 391841 26283 391907 26286
rect 419441 26283 419507 26286
rect 445661 26283 445727 26286
rect 500861 26283 500927 26286
rect 526437 26283 526503 26286
rect 367010 26150 367172 26210
rect 35758 25636 35818 26150
rect 38009 26147 38075 26150
rect 146293 25938 146359 25941
rect 253933 25938 253999 25941
rect 361573 25938 361639 25941
rect 469213 25938 469279 25941
rect 143766 25936 146359 25938
rect 143766 25880 146298 25936
rect 146354 25880 146359 25936
rect 143766 25878 146359 25880
rect 64873 25666 64939 25669
rect 91093 25666 91159 25669
rect 118693 25666 118759 25669
rect 62836 25664 64939 25666
rect 62836 25608 64878 25664
rect 64934 25608 64939 25664
rect 62836 25606 64939 25608
rect 89884 25664 91159 25666
rect 89884 25608 91098 25664
rect 91154 25608 91159 25664
rect 89884 25606 91159 25608
rect 116932 25664 118759 25666
rect 116932 25608 118698 25664
rect 118754 25608 118759 25664
rect 143766 25636 143826 25878
rect 146293 25875 146359 25878
rect 251774 25936 253999 25938
rect 251774 25880 253938 25936
rect 253994 25880 253999 25936
rect 251774 25878 253999 25880
rect 172513 25666 172579 25669
rect 200113 25666 200179 25669
rect 226333 25666 226399 25669
rect 170844 25664 172579 25666
rect 116932 25606 118759 25608
rect 170844 25608 172518 25664
rect 172574 25608 172579 25664
rect 170844 25606 172579 25608
rect 197892 25664 200179 25666
rect 197892 25608 200118 25664
rect 200174 25608 200179 25664
rect 197892 25606 200179 25608
rect 224940 25664 226399 25666
rect 224940 25608 226338 25664
rect 226394 25608 226399 25664
rect 251774 25636 251834 25878
rect 253933 25875 253999 25878
rect 359782 25936 361639 25938
rect 359782 25880 361578 25936
rect 361634 25880 361639 25936
rect 359782 25878 361639 25880
rect 280153 25666 280219 25669
rect 307753 25666 307819 25669
rect 335353 25666 335419 25669
rect 278852 25664 280219 25666
rect 224940 25606 226399 25608
rect 278852 25608 280158 25664
rect 280214 25608 280219 25664
rect 278852 25606 280219 25608
rect 305900 25664 307819 25666
rect 305900 25608 307758 25664
rect 307814 25608 307819 25664
rect 305900 25606 307819 25608
rect 332948 25664 335419 25666
rect 332948 25608 335358 25664
rect 335414 25608 335419 25664
rect 359782 25636 359842 25878
rect 361573 25875 361639 25878
rect 467790 25936 469279 25938
rect 467790 25880 469218 25936
rect 469274 25880 469279 25936
rect 467790 25878 469279 25880
rect 389173 25666 389239 25669
rect 415393 25666 415459 25669
rect 442993 25666 443059 25669
rect 386860 25664 389239 25666
rect 332948 25606 335419 25608
rect 386860 25608 389178 25664
rect 389234 25608 389239 25664
rect 386860 25606 389239 25608
rect 413908 25664 415459 25666
rect 413908 25608 415398 25664
rect 415454 25608 415459 25664
rect 413908 25606 415459 25608
rect 440956 25664 443059 25666
rect 440956 25608 442998 25664
rect 443054 25608 443059 25664
rect 467790 25636 467850 25878
rect 469213 25875 469279 25878
rect 496813 25666 496879 25669
rect 523033 25666 523099 25669
rect 550633 25666 550699 25669
rect 494868 25664 496879 25666
rect 440956 25606 443059 25608
rect 494868 25608 496818 25664
rect 496874 25608 496879 25664
rect 494868 25606 496879 25608
rect 521916 25664 523099 25666
rect 521916 25608 523038 25664
rect 523094 25608 523099 25664
rect 521916 25606 523099 25608
rect 548964 25664 550699 25666
rect 548964 25608 550638 25664
rect 550694 25608 550699 25664
rect 548964 25606 550699 25608
rect 64873 25603 64939 25606
rect 91093 25603 91159 25606
rect 118693 25603 118759 25606
rect 172513 25603 172579 25606
rect 200113 25603 200179 25606
rect 226333 25603 226399 25606
rect 280153 25603 280219 25606
rect 307753 25603 307819 25606
rect 335353 25603 335419 25606
rect 389173 25603 389239 25606
rect 415393 25603 415459 25606
rect 442993 25603 443059 25606
rect 496813 25603 496879 25606
rect 523033 25603 523099 25606
rect 550633 25603 550699 25606
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 583520 6476 584960 6716
<< metal4 >>
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 696454 -2346 705242
rect -2966 696218 -2934 696454
rect -2698 696218 -2614 696454
rect -2378 696218 -2346 696454
rect -2966 696134 -2346 696218
rect -2966 695898 -2934 696134
rect -2698 695898 -2614 696134
rect -2378 695898 -2346 696134
rect -2966 678454 -2346 695898
rect -2966 678218 -2934 678454
rect -2698 678218 -2614 678454
rect -2378 678218 -2346 678454
rect -2966 678134 -2346 678218
rect -2966 677898 -2934 678134
rect -2698 677898 -2614 678134
rect -2378 677898 -2346 678134
rect -2966 660454 -2346 677898
rect -2966 660218 -2934 660454
rect -2698 660218 -2614 660454
rect -2378 660218 -2346 660454
rect -2966 660134 -2346 660218
rect -2966 659898 -2934 660134
rect -2698 659898 -2614 660134
rect -2378 659898 -2346 660134
rect -2966 642454 -2346 659898
rect -2966 642218 -2934 642454
rect -2698 642218 -2614 642454
rect -2378 642218 -2346 642454
rect -2966 642134 -2346 642218
rect -2966 641898 -2934 642134
rect -2698 641898 -2614 642134
rect -2378 641898 -2346 642134
rect -2966 624454 -2346 641898
rect -2966 624218 -2934 624454
rect -2698 624218 -2614 624454
rect -2378 624218 -2346 624454
rect -2966 624134 -2346 624218
rect -2966 623898 -2934 624134
rect -2698 623898 -2614 624134
rect -2378 623898 -2346 624134
rect -2966 606454 -2346 623898
rect -2966 606218 -2934 606454
rect -2698 606218 -2614 606454
rect -2378 606218 -2346 606454
rect -2966 606134 -2346 606218
rect -2966 605898 -2934 606134
rect -2698 605898 -2614 606134
rect -2378 605898 -2346 606134
rect -2966 588454 -2346 605898
rect -2966 588218 -2934 588454
rect -2698 588218 -2614 588454
rect -2378 588218 -2346 588454
rect -2966 588134 -2346 588218
rect -2966 587898 -2934 588134
rect -2698 587898 -2614 588134
rect -2378 587898 -2346 588134
rect -2966 570454 -2346 587898
rect -2966 570218 -2934 570454
rect -2698 570218 -2614 570454
rect -2378 570218 -2346 570454
rect -2966 570134 -2346 570218
rect -2966 569898 -2934 570134
rect -2698 569898 -2614 570134
rect -2378 569898 -2346 570134
rect -2966 552454 -2346 569898
rect -2966 552218 -2934 552454
rect -2698 552218 -2614 552454
rect -2378 552218 -2346 552454
rect -2966 552134 -2346 552218
rect -2966 551898 -2934 552134
rect -2698 551898 -2614 552134
rect -2378 551898 -2346 552134
rect -2966 534454 -2346 551898
rect -2966 534218 -2934 534454
rect -2698 534218 -2614 534454
rect -2378 534218 -2346 534454
rect -2966 534134 -2346 534218
rect -2966 533898 -2934 534134
rect -2698 533898 -2614 534134
rect -2378 533898 -2346 534134
rect -2966 516454 -2346 533898
rect -2966 516218 -2934 516454
rect -2698 516218 -2614 516454
rect -2378 516218 -2346 516454
rect -2966 516134 -2346 516218
rect -2966 515898 -2934 516134
rect -2698 515898 -2614 516134
rect -2378 515898 -2346 516134
rect -2966 498454 -2346 515898
rect -2966 498218 -2934 498454
rect -2698 498218 -2614 498454
rect -2378 498218 -2346 498454
rect -2966 498134 -2346 498218
rect -2966 497898 -2934 498134
rect -2698 497898 -2614 498134
rect -2378 497898 -2346 498134
rect -2966 480454 -2346 497898
rect -2966 480218 -2934 480454
rect -2698 480218 -2614 480454
rect -2378 480218 -2346 480454
rect -2966 480134 -2346 480218
rect -2966 479898 -2934 480134
rect -2698 479898 -2614 480134
rect -2378 479898 -2346 480134
rect -2966 462454 -2346 479898
rect -2966 462218 -2934 462454
rect -2698 462218 -2614 462454
rect -2378 462218 -2346 462454
rect -2966 462134 -2346 462218
rect -2966 461898 -2934 462134
rect -2698 461898 -2614 462134
rect -2378 461898 -2346 462134
rect -2966 444454 -2346 461898
rect -2966 444218 -2934 444454
rect -2698 444218 -2614 444454
rect -2378 444218 -2346 444454
rect -2966 444134 -2346 444218
rect -2966 443898 -2934 444134
rect -2698 443898 -2614 444134
rect -2378 443898 -2346 444134
rect -2966 426454 -2346 443898
rect -2966 426218 -2934 426454
rect -2698 426218 -2614 426454
rect -2378 426218 -2346 426454
rect -2966 426134 -2346 426218
rect -2966 425898 -2934 426134
rect -2698 425898 -2614 426134
rect -2378 425898 -2346 426134
rect -2966 408454 -2346 425898
rect -2966 408218 -2934 408454
rect -2698 408218 -2614 408454
rect -2378 408218 -2346 408454
rect -2966 408134 -2346 408218
rect -2966 407898 -2934 408134
rect -2698 407898 -2614 408134
rect -2378 407898 -2346 408134
rect -2966 390454 -2346 407898
rect -2966 390218 -2934 390454
rect -2698 390218 -2614 390454
rect -2378 390218 -2346 390454
rect -2966 390134 -2346 390218
rect -2966 389898 -2934 390134
rect -2698 389898 -2614 390134
rect -2378 389898 -2346 390134
rect -2966 372454 -2346 389898
rect -2966 372218 -2934 372454
rect -2698 372218 -2614 372454
rect -2378 372218 -2346 372454
rect -2966 372134 -2346 372218
rect -2966 371898 -2934 372134
rect -2698 371898 -2614 372134
rect -2378 371898 -2346 372134
rect -2966 354454 -2346 371898
rect -2966 354218 -2934 354454
rect -2698 354218 -2614 354454
rect -2378 354218 -2346 354454
rect -2966 354134 -2346 354218
rect -2966 353898 -2934 354134
rect -2698 353898 -2614 354134
rect -2378 353898 -2346 354134
rect -2966 336454 -2346 353898
rect -2966 336218 -2934 336454
rect -2698 336218 -2614 336454
rect -2378 336218 -2346 336454
rect -2966 336134 -2346 336218
rect -2966 335898 -2934 336134
rect -2698 335898 -2614 336134
rect -2378 335898 -2346 336134
rect -2966 318454 -2346 335898
rect -2966 318218 -2934 318454
rect -2698 318218 -2614 318454
rect -2378 318218 -2346 318454
rect -2966 318134 -2346 318218
rect -2966 317898 -2934 318134
rect -2698 317898 -2614 318134
rect -2378 317898 -2346 318134
rect -2966 300454 -2346 317898
rect -2966 300218 -2934 300454
rect -2698 300218 -2614 300454
rect -2378 300218 -2346 300454
rect -2966 300134 -2346 300218
rect -2966 299898 -2934 300134
rect -2698 299898 -2614 300134
rect -2378 299898 -2346 300134
rect -2966 282454 -2346 299898
rect -2966 282218 -2934 282454
rect -2698 282218 -2614 282454
rect -2378 282218 -2346 282454
rect -2966 282134 -2346 282218
rect -2966 281898 -2934 282134
rect -2698 281898 -2614 282134
rect -2378 281898 -2346 282134
rect -2966 264454 -2346 281898
rect -2966 264218 -2934 264454
rect -2698 264218 -2614 264454
rect -2378 264218 -2346 264454
rect -2966 264134 -2346 264218
rect -2966 263898 -2934 264134
rect -2698 263898 -2614 264134
rect -2378 263898 -2346 264134
rect -2966 246454 -2346 263898
rect -2966 246218 -2934 246454
rect -2698 246218 -2614 246454
rect -2378 246218 -2346 246454
rect -2966 246134 -2346 246218
rect -2966 245898 -2934 246134
rect -2698 245898 -2614 246134
rect -2378 245898 -2346 246134
rect -2966 228454 -2346 245898
rect -2966 228218 -2934 228454
rect -2698 228218 -2614 228454
rect -2378 228218 -2346 228454
rect -2966 228134 -2346 228218
rect -2966 227898 -2934 228134
rect -2698 227898 -2614 228134
rect -2378 227898 -2346 228134
rect -2966 210454 -2346 227898
rect -2966 210218 -2934 210454
rect -2698 210218 -2614 210454
rect -2378 210218 -2346 210454
rect -2966 210134 -2346 210218
rect -2966 209898 -2934 210134
rect -2698 209898 -2614 210134
rect -2378 209898 -2346 210134
rect -2966 192454 -2346 209898
rect -2966 192218 -2934 192454
rect -2698 192218 -2614 192454
rect -2378 192218 -2346 192454
rect -2966 192134 -2346 192218
rect -2966 191898 -2934 192134
rect -2698 191898 -2614 192134
rect -2378 191898 -2346 192134
rect -2966 174454 -2346 191898
rect -2966 174218 -2934 174454
rect -2698 174218 -2614 174454
rect -2378 174218 -2346 174454
rect -2966 174134 -2346 174218
rect -2966 173898 -2934 174134
rect -2698 173898 -2614 174134
rect -2378 173898 -2346 174134
rect -2966 156454 -2346 173898
rect -2966 156218 -2934 156454
rect -2698 156218 -2614 156454
rect -2378 156218 -2346 156454
rect -2966 156134 -2346 156218
rect -2966 155898 -2934 156134
rect -2698 155898 -2614 156134
rect -2378 155898 -2346 156134
rect -2966 138454 -2346 155898
rect -2966 138218 -2934 138454
rect -2698 138218 -2614 138454
rect -2378 138218 -2346 138454
rect -2966 138134 -2346 138218
rect -2966 137898 -2934 138134
rect -2698 137898 -2614 138134
rect -2378 137898 -2346 138134
rect -2966 120454 -2346 137898
rect -2966 120218 -2934 120454
rect -2698 120218 -2614 120454
rect -2378 120218 -2346 120454
rect -2966 120134 -2346 120218
rect -2966 119898 -2934 120134
rect -2698 119898 -2614 120134
rect -2378 119898 -2346 120134
rect -2966 102454 -2346 119898
rect -2966 102218 -2934 102454
rect -2698 102218 -2614 102454
rect -2378 102218 -2346 102454
rect -2966 102134 -2346 102218
rect -2966 101898 -2934 102134
rect -2698 101898 -2614 102134
rect -2378 101898 -2346 102134
rect -2966 84454 -2346 101898
rect -2966 84218 -2934 84454
rect -2698 84218 -2614 84454
rect -2378 84218 -2346 84454
rect -2966 84134 -2346 84218
rect -2966 83898 -2934 84134
rect -2698 83898 -2614 84134
rect -2378 83898 -2346 84134
rect -2966 66454 -2346 83898
rect -2966 66218 -2934 66454
rect -2698 66218 -2614 66454
rect -2378 66218 -2346 66454
rect -2966 66134 -2346 66218
rect -2966 65898 -2934 66134
rect -2698 65898 -2614 66134
rect -2378 65898 -2346 66134
rect -2966 48454 -2346 65898
rect -2966 48218 -2934 48454
rect -2698 48218 -2614 48454
rect -2378 48218 -2346 48454
rect -2966 48134 -2346 48218
rect -2966 47898 -2934 48134
rect -2698 47898 -2614 48134
rect -2378 47898 -2346 48134
rect -2966 30454 -2346 47898
rect -2966 30218 -2934 30454
rect -2698 30218 -2614 30454
rect -2378 30218 -2346 30454
rect -2966 30134 -2346 30218
rect -2966 29898 -2934 30134
rect -2698 29898 -2614 30134
rect -2378 29898 -2346 30134
rect -2966 12454 -2346 29898
rect -2966 12218 -2934 12454
rect -2698 12218 -2614 12454
rect -2378 12218 -2346 12454
rect -2966 12134 -2346 12218
rect -2966 11898 -2934 12134
rect -2698 11898 -2614 12134
rect -2378 11898 -2346 12134
rect -2966 -1306 -2346 11898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 669454 -1386 686898
rect -2006 669218 -1974 669454
rect -1738 669218 -1654 669454
rect -1418 669218 -1386 669454
rect -2006 669134 -1386 669218
rect -2006 668898 -1974 669134
rect -1738 668898 -1654 669134
rect -1418 668898 -1386 669134
rect -2006 651454 -1386 668898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 633454 -1386 650898
rect -2006 633218 -1974 633454
rect -1738 633218 -1654 633454
rect -1418 633218 -1386 633454
rect -2006 633134 -1386 633218
rect -2006 632898 -1974 633134
rect -1738 632898 -1654 633134
rect -1418 632898 -1386 633134
rect -2006 615454 -1386 632898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 597454 -1386 614898
rect -2006 597218 -1974 597454
rect -1738 597218 -1654 597454
rect -1418 597218 -1386 597454
rect -2006 597134 -1386 597218
rect -2006 596898 -1974 597134
rect -1738 596898 -1654 597134
rect -1418 596898 -1386 597134
rect -2006 579454 -1386 596898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 561454 -1386 578898
rect -2006 561218 -1974 561454
rect -1738 561218 -1654 561454
rect -1418 561218 -1386 561454
rect -2006 561134 -1386 561218
rect -2006 560898 -1974 561134
rect -1738 560898 -1654 561134
rect -1418 560898 -1386 561134
rect -2006 543454 -1386 560898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 525454 -1386 542898
rect -2006 525218 -1974 525454
rect -1738 525218 -1654 525454
rect -1418 525218 -1386 525454
rect -2006 525134 -1386 525218
rect -2006 524898 -1974 525134
rect -1738 524898 -1654 525134
rect -1418 524898 -1386 525134
rect -2006 507454 -1386 524898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 489454 -1386 506898
rect -2006 489218 -1974 489454
rect -1738 489218 -1654 489454
rect -1418 489218 -1386 489454
rect -2006 489134 -1386 489218
rect -2006 488898 -1974 489134
rect -1738 488898 -1654 489134
rect -1418 488898 -1386 489134
rect -2006 471454 -1386 488898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 453454 -1386 470898
rect -2006 453218 -1974 453454
rect -1738 453218 -1654 453454
rect -1418 453218 -1386 453454
rect -2006 453134 -1386 453218
rect -2006 452898 -1974 453134
rect -1738 452898 -1654 453134
rect -1418 452898 -1386 453134
rect -2006 435454 -1386 452898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 417454 -1386 434898
rect -2006 417218 -1974 417454
rect -1738 417218 -1654 417454
rect -1418 417218 -1386 417454
rect -2006 417134 -1386 417218
rect -2006 416898 -1974 417134
rect -1738 416898 -1654 417134
rect -1418 416898 -1386 417134
rect -2006 399454 -1386 416898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 381454 -1386 398898
rect -2006 381218 -1974 381454
rect -1738 381218 -1654 381454
rect -1418 381218 -1386 381454
rect -2006 381134 -1386 381218
rect -2006 380898 -1974 381134
rect -1738 380898 -1654 381134
rect -1418 380898 -1386 381134
rect -2006 363454 -1386 380898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 345454 -1386 362898
rect -2006 345218 -1974 345454
rect -1738 345218 -1654 345454
rect -1418 345218 -1386 345454
rect -2006 345134 -1386 345218
rect -2006 344898 -1974 345134
rect -1738 344898 -1654 345134
rect -1418 344898 -1386 345134
rect -2006 327454 -1386 344898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 309454 -1386 326898
rect -2006 309218 -1974 309454
rect -1738 309218 -1654 309454
rect -1418 309218 -1386 309454
rect -2006 309134 -1386 309218
rect -2006 308898 -1974 309134
rect -1738 308898 -1654 309134
rect -1418 308898 -1386 309134
rect -2006 291454 -1386 308898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 273454 -1386 290898
rect -2006 273218 -1974 273454
rect -1738 273218 -1654 273454
rect -1418 273218 -1386 273454
rect -2006 273134 -1386 273218
rect -2006 272898 -1974 273134
rect -1738 272898 -1654 273134
rect -1418 272898 -1386 273134
rect -2006 255454 -1386 272898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 237454 -1386 254898
rect -2006 237218 -1974 237454
rect -1738 237218 -1654 237454
rect -1418 237218 -1386 237454
rect -2006 237134 -1386 237218
rect -2006 236898 -1974 237134
rect -1738 236898 -1654 237134
rect -1418 236898 -1386 237134
rect -2006 219454 -1386 236898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 201454 -1386 218898
rect -2006 201218 -1974 201454
rect -1738 201218 -1654 201454
rect -1418 201218 -1386 201454
rect -2006 201134 -1386 201218
rect -2006 200898 -1974 201134
rect -1738 200898 -1654 201134
rect -1418 200898 -1386 201134
rect -2006 183454 -1386 200898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 165454 -1386 182898
rect -2006 165218 -1974 165454
rect -1738 165218 -1654 165454
rect -1418 165218 -1386 165454
rect -2006 165134 -1386 165218
rect -2006 164898 -1974 165134
rect -1738 164898 -1654 165134
rect -1418 164898 -1386 165134
rect -2006 147454 -1386 164898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 129454 -1386 146898
rect -2006 129218 -1974 129454
rect -1738 129218 -1654 129454
rect -1418 129218 -1386 129454
rect -2006 129134 -1386 129218
rect -2006 128898 -1974 129134
rect -1738 128898 -1654 129134
rect -1418 128898 -1386 129134
rect -2006 111454 -1386 128898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 93454 -1386 110898
rect -2006 93218 -1974 93454
rect -1738 93218 -1654 93454
rect -1418 93218 -1386 93454
rect -2006 93134 -1386 93218
rect -2006 92898 -1974 93134
rect -1738 92898 -1654 93134
rect -1418 92898 -1386 93134
rect -2006 75454 -1386 92898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 57454 -1386 74898
rect -2006 57218 -1974 57454
rect -1738 57218 -1654 57454
rect -1418 57218 -1386 57454
rect -2006 57134 -1386 57218
rect -2006 56898 -1974 57134
rect -1738 56898 -1654 57134
rect -1418 56898 -1386 57134
rect -2006 39454 -1386 56898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 21454 -1386 38898
rect -2006 21218 -1974 21454
rect -1738 21218 -1654 21454
rect -1418 21218 -1386 21454
rect -2006 21134 -1386 21218
rect -2006 20898 -1974 21134
rect -1738 20898 -1654 21134
rect -1418 20898 -1386 21134
rect -2006 3454 -1386 20898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 669454 2414 686898
rect 1794 669218 1826 669454
rect 2062 669218 2146 669454
rect 2382 669218 2414 669454
rect 1794 669134 2414 669218
rect 1794 668898 1826 669134
rect 2062 668898 2146 669134
rect 2382 668898 2414 669134
rect 1794 651454 2414 668898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 633454 2414 650898
rect 1794 633218 1826 633454
rect 2062 633218 2146 633454
rect 2382 633218 2414 633454
rect 1794 633134 2414 633218
rect 1794 632898 1826 633134
rect 2062 632898 2146 633134
rect 2382 632898 2414 633134
rect 1794 615454 2414 632898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 597454 2414 614898
rect 1794 597218 1826 597454
rect 2062 597218 2146 597454
rect 2382 597218 2414 597454
rect 1794 597134 2414 597218
rect 1794 596898 1826 597134
rect 2062 596898 2146 597134
rect 2382 596898 2414 597134
rect 1794 579454 2414 596898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 561454 2414 578898
rect 1794 561218 1826 561454
rect 2062 561218 2146 561454
rect 2382 561218 2414 561454
rect 1794 561134 2414 561218
rect 1794 560898 1826 561134
rect 2062 560898 2146 561134
rect 2382 560898 2414 561134
rect 1794 543454 2414 560898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 525454 2414 542898
rect 1794 525218 1826 525454
rect 2062 525218 2146 525454
rect 2382 525218 2414 525454
rect 1794 525134 2414 525218
rect 1794 524898 1826 525134
rect 2062 524898 2146 525134
rect 2382 524898 2414 525134
rect 1794 507454 2414 524898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 489454 2414 506898
rect 1794 489218 1826 489454
rect 2062 489218 2146 489454
rect 2382 489218 2414 489454
rect 1794 489134 2414 489218
rect 1794 488898 1826 489134
rect 2062 488898 2146 489134
rect 2382 488898 2414 489134
rect 1794 471454 2414 488898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 453454 2414 470898
rect 1794 453218 1826 453454
rect 2062 453218 2146 453454
rect 2382 453218 2414 453454
rect 1794 453134 2414 453218
rect 1794 452898 1826 453134
rect 2062 452898 2146 453134
rect 2382 452898 2414 453134
rect 1794 435454 2414 452898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 417454 2414 434898
rect 1794 417218 1826 417454
rect 2062 417218 2146 417454
rect 2382 417218 2414 417454
rect 1794 417134 2414 417218
rect 1794 416898 1826 417134
rect 2062 416898 2146 417134
rect 2382 416898 2414 417134
rect 1794 399454 2414 416898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 381454 2414 398898
rect 1794 381218 1826 381454
rect 2062 381218 2146 381454
rect 2382 381218 2414 381454
rect 1794 381134 2414 381218
rect 1794 380898 1826 381134
rect 2062 380898 2146 381134
rect 2382 380898 2414 381134
rect 1794 363454 2414 380898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 345454 2414 362898
rect 1794 345218 1826 345454
rect 2062 345218 2146 345454
rect 2382 345218 2414 345454
rect 1794 345134 2414 345218
rect 1794 344898 1826 345134
rect 2062 344898 2146 345134
rect 2382 344898 2414 345134
rect 1794 327454 2414 344898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 309454 2414 326898
rect 1794 309218 1826 309454
rect 2062 309218 2146 309454
rect 2382 309218 2414 309454
rect 1794 309134 2414 309218
rect 1794 308898 1826 309134
rect 2062 308898 2146 309134
rect 2382 308898 2414 309134
rect 1794 291454 2414 308898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 273454 2414 290898
rect 1794 273218 1826 273454
rect 2062 273218 2146 273454
rect 2382 273218 2414 273454
rect 1794 273134 2414 273218
rect 1794 272898 1826 273134
rect 2062 272898 2146 273134
rect 2382 272898 2414 273134
rect 1794 255454 2414 272898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 237454 2414 254898
rect 1794 237218 1826 237454
rect 2062 237218 2146 237454
rect 2382 237218 2414 237454
rect 1794 237134 2414 237218
rect 1794 236898 1826 237134
rect 2062 236898 2146 237134
rect 2382 236898 2414 237134
rect 1794 219454 2414 236898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 201454 2414 218898
rect 1794 201218 1826 201454
rect 2062 201218 2146 201454
rect 2382 201218 2414 201454
rect 1794 201134 2414 201218
rect 1794 200898 1826 201134
rect 2062 200898 2146 201134
rect 2382 200898 2414 201134
rect 1794 183454 2414 200898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 165454 2414 182898
rect 1794 165218 1826 165454
rect 2062 165218 2146 165454
rect 2382 165218 2414 165454
rect 1794 165134 2414 165218
rect 1794 164898 1826 165134
rect 2062 164898 2146 165134
rect 2382 164898 2414 165134
rect 1794 147454 2414 164898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 129454 2414 146898
rect 1794 129218 1826 129454
rect 2062 129218 2146 129454
rect 2382 129218 2414 129454
rect 1794 129134 2414 129218
rect 1794 128898 1826 129134
rect 2062 128898 2146 129134
rect 2382 128898 2414 129134
rect 1794 111454 2414 128898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 93454 2414 110898
rect 1794 93218 1826 93454
rect 2062 93218 2146 93454
rect 2382 93218 2414 93454
rect 1794 93134 2414 93218
rect 1794 92898 1826 93134
rect 2062 92898 2146 93134
rect 2382 92898 2414 93134
rect 1794 75454 2414 92898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 57454 2414 74898
rect 1794 57218 1826 57454
rect 2062 57218 2146 57454
rect 2382 57218 2414 57454
rect 1794 57134 2414 57218
rect 1794 56898 1826 57134
rect 2062 56898 2146 57134
rect 2382 56898 2414 57134
rect 1794 39454 2414 56898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 21454 2414 38898
rect 1794 21218 1826 21454
rect 2062 21218 2146 21454
rect 2382 21218 2414 21454
rect 1794 21134 2414 21218
rect 1794 20898 1826 21134
rect 2062 20898 2146 21134
rect 2382 20898 2414 21134
rect 1794 3454 2414 20898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 10794 705798 11414 705830
rect 10794 705562 10826 705798
rect 11062 705562 11146 705798
rect 11382 705562 11414 705798
rect 10794 705478 11414 705562
rect 10794 705242 10826 705478
rect 11062 705242 11146 705478
rect 11382 705242 11414 705478
rect 10794 696454 11414 705242
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 678454 11414 695898
rect 19794 704838 20414 705830
rect 19794 704602 19826 704838
rect 20062 704602 20146 704838
rect 20382 704602 20414 704838
rect 19794 704518 20414 704602
rect 19794 704282 19826 704518
rect 20062 704282 20146 704518
rect 20382 704282 20414 704518
rect 19794 687454 20414 704282
rect 19794 687218 19826 687454
rect 20062 687218 20146 687454
rect 20382 687218 20414 687454
rect 19794 687134 20414 687218
rect 19794 686898 19826 687134
rect 20062 686898 20146 687134
rect 20382 686898 20414 687134
rect 19794 686000 20414 686898
rect 28794 705798 29414 705830
rect 28794 705562 28826 705798
rect 29062 705562 29146 705798
rect 29382 705562 29414 705798
rect 28794 705478 29414 705562
rect 28794 705242 28826 705478
rect 29062 705242 29146 705478
rect 29382 705242 29414 705478
rect 28794 696454 29414 705242
rect 28794 696218 28826 696454
rect 29062 696218 29146 696454
rect 29382 696218 29414 696454
rect 28794 696134 29414 696218
rect 28794 695898 28826 696134
rect 29062 695898 29146 696134
rect 29382 695898 29414 696134
rect 28794 686000 29414 695898
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 686000 38414 686898
rect 46794 705798 47414 705830
rect 46794 705562 46826 705798
rect 47062 705562 47146 705798
rect 47382 705562 47414 705798
rect 46794 705478 47414 705562
rect 46794 705242 46826 705478
rect 47062 705242 47146 705478
rect 47382 705242 47414 705478
rect 46794 696454 47414 705242
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 686000 47414 695898
rect 55794 704838 56414 705830
rect 55794 704602 55826 704838
rect 56062 704602 56146 704838
rect 56382 704602 56414 704838
rect 55794 704518 56414 704602
rect 55794 704282 55826 704518
rect 56062 704282 56146 704518
rect 56382 704282 56414 704518
rect 55794 687454 56414 704282
rect 55794 687218 55826 687454
rect 56062 687218 56146 687454
rect 56382 687218 56414 687454
rect 55794 687134 56414 687218
rect 55794 686898 55826 687134
rect 56062 686898 56146 687134
rect 56382 686898 56414 687134
rect 55794 686000 56414 686898
rect 64794 705798 65414 705830
rect 64794 705562 64826 705798
rect 65062 705562 65146 705798
rect 65382 705562 65414 705798
rect 64794 705478 65414 705562
rect 64794 705242 64826 705478
rect 65062 705242 65146 705478
rect 65382 705242 65414 705478
rect 64794 696454 65414 705242
rect 64794 696218 64826 696454
rect 65062 696218 65146 696454
rect 65382 696218 65414 696454
rect 64794 696134 65414 696218
rect 64794 695898 64826 696134
rect 65062 695898 65146 696134
rect 65382 695898 65414 696134
rect 64794 686000 65414 695898
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 686000 74414 686898
rect 82794 705798 83414 705830
rect 82794 705562 82826 705798
rect 83062 705562 83146 705798
rect 83382 705562 83414 705798
rect 82794 705478 83414 705562
rect 82794 705242 82826 705478
rect 83062 705242 83146 705478
rect 83382 705242 83414 705478
rect 82794 696454 83414 705242
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 686000 83414 695898
rect 91794 704838 92414 705830
rect 91794 704602 91826 704838
rect 92062 704602 92146 704838
rect 92382 704602 92414 704838
rect 91794 704518 92414 704602
rect 91794 704282 91826 704518
rect 92062 704282 92146 704518
rect 92382 704282 92414 704518
rect 91794 687454 92414 704282
rect 91794 687218 91826 687454
rect 92062 687218 92146 687454
rect 92382 687218 92414 687454
rect 91794 687134 92414 687218
rect 91794 686898 91826 687134
rect 92062 686898 92146 687134
rect 92382 686898 92414 687134
rect 91794 686000 92414 686898
rect 100794 705798 101414 705830
rect 100794 705562 100826 705798
rect 101062 705562 101146 705798
rect 101382 705562 101414 705798
rect 100794 705478 101414 705562
rect 100794 705242 100826 705478
rect 101062 705242 101146 705478
rect 101382 705242 101414 705478
rect 100794 696454 101414 705242
rect 100794 696218 100826 696454
rect 101062 696218 101146 696454
rect 101382 696218 101414 696454
rect 100794 696134 101414 696218
rect 100794 695898 100826 696134
rect 101062 695898 101146 696134
rect 101382 695898 101414 696134
rect 100794 686000 101414 695898
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 686000 110414 686898
rect 118794 705798 119414 705830
rect 118794 705562 118826 705798
rect 119062 705562 119146 705798
rect 119382 705562 119414 705798
rect 118794 705478 119414 705562
rect 118794 705242 118826 705478
rect 119062 705242 119146 705478
rect 119382 705242 119414 705478
rect 118794 696454 119414 705242
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 686000 119414 695898
rect 127794 704838 128414 705830
rect 127794 704602 127826 704838
rect 128062 704602 128146 704838
rect 128382 704602 128414 704838
rect 127794 704518 128414 704602
rect 127794 704282 127826 704518
rect 128062 704282 128146 704518
rect 128382 704282 128414 704518
rect 127794 687454 128414 704282
rect 127794 687218 127826 687454
rect 128062 687218 128146 687454
rect 128382 687218 128414 687454
rect 127794 687134 128414 687218
rect 127794 686898 127826 687134
rect 128062 686898 128146 687134
rect 128382 686898 128414 687134
rect 127794 686000 128414 686898
rect 136794 705798 137414 705830
rect 136794 705562 136826 705798
rect 137062 705562 137146 705798
rect 137382 705562 137414 705798
rect 136794 705478 137414 705562
rect 136794 705242 136826 705478
rect 137062 705242 137146 705478
rect 137382 705242 137414 705478
rect 136794 696454 137414 705242
rect 136794 696218 136826 696454
rect 137062 696218 137146 696454
rect 137382 696218 137414 696454
rect 136794 696134 137414 696218
rect 136794 695898 136826 696134
rect 137062 695898 137146 696134
rect 137382 695898 137414 696134
rect 136794 686000 137414 695898
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 686000 146414 686898
rect 154794 705798 155414 705830
rect 154794 705562 154826 705798
rect 155062 705562 155146 705798
rect 155382 705562 155414 705798
rect 154794 705478 155414 705562
rect 154794 705242 154826 705478
rect 155062 705242 155146 705478
rect 155382 705242 155414 705478
rect 154794 696454 155414 705242
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 686000 155414 695898
rect 163794 704838 164414 705830
rect 163794 704602 163826 704838
rect 164062 704602 164146 704838
rect 164382 704602 164414 704838
rect 163794 704518 164414 704602
rect 163794 704282 163826 704518
rect 164062 704282 164146 704518
rect 164382 704282 164414 704518
rect 163794 687454 164414 704282
rect 163794 687218 163826 687454
rect 164062 687218 164146 687454
rect 164382 687218 164414 687454
rect 163794 687134 164414 687218
rect 163794 686898 163826 687134
rect 164062 686898 164146 687134
rect 164382 686898 164414 687134
rect 163794 686000 164414 686898
rect 172794 705798 173414 705830
rect 172794 705562 172826 705798
rect 173062 705562 173146 705798
rect 173382 705562 173414 705798
rect 172794 705478 173414 705562
rect 172794 705242 172826 705478
rect 173062 705242 173146 705478
rect 173382 705242 173414 705478
rect 172794 696454 173414 705242
rect 172794 696218 172826 696454
rect 173062 696218 173146 696454
rect 173382 696218 173414 696454
rect 172794 696134 173414 696218
rect 172794 695898 172826 696134
rect 173062 695898 173146 696134
rect 173382 695898 173414 696134
rect 172794 686000 173414 695898
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 686000 182414 686898
rect 190794 705798 191414 705830
rect 190794 705562 190826 705798
rect 191062 705562 191146 705798
rect 191382 705562 191414 705798
rect 190794 705478 191414 705562
rect 190794 705242 190826 705478
rect 191062 705242 191146 705478
rect 191382 705242 191414 705478
rect 190794 696454 191414 705242
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 686000 191414 695898
rect 199794 704838 200414 705830
rect 199794 704602 199826 704838
rect 200062 704602 200146 704838
rect 200382 704602 200414 704838
rect 199794 704518 200414 704602
rect 199794 704282 199826 704518
rect 200062 704282 200146 704518
rect 200382 704282 200414 704518
rect 199794 687454 200414 704282
rect 199794 687218 199826 687454
rect 200062 687218 200146 687454
rect 200382 687218 200414 687454
rect 199794 687134 200414 687218
rect 199794 686898 199826 687134
rect 200062 686898 200146 687134
rect 200382 686898 200414 687134
rect 199794 686000 200414 686898
rect 208794 705798 209414 705830
rect 208794 705562 208826 705798
rect 209062 705562 209146 705798
rect 209382 705562 209414 705798
rect 208794 705478 209414 705562
rect 208794 705242 208826 705478
rect 209062 705242 209146 705478
rect 209382 705242 209414 705478
rect 208794 696454 209414 705242
rect 208794 696218 208826 696454
rect 209062 696218 209146 696454
rect 209382 696218 209414 696454
rect 208794 696134 209414 696218
rect 208794 695898 208826 696134
rect 209062 695898 209146 696134
rect 209382 695898 209414 696134
rect 208794 686000 209414 695898
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 686000 218414 686898
rect 226794 705798 227414 705830
rect 226794 705562 226826 705798
rect 227062 705562 227146 705798
rect 227382 705562 227414 705798
rect 226794 705478 227414 705562
rect 226794 705242 226826 705478
rect 227062 705242 227146 705478
rect 227382 705242 227414 705478
rect 226794 696454 227414 705242
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 686000 227414 695898
rect 235794 704838 236414 705830
rect 235794 704602 235826 704838
rect 236062 704602 236146 704838
rect 236382 704602 236414 704838
rect 235794 704518 236414 704602
rect 235794 704282 235826 704518
rect 236062 704282 236146 704518
rect 236382 704282 236414 704518
rect 235794 687454 236414 704282
rect 235794 687218 235826 687454
rect 236062 687218 236146 687454
rect 236382 687218 236414 687454
rect 235794 687134 236414 687218
rect 235794 686898 235826 687134
rect 236062 686898 236146 687134
rect 236382 686898 236414 687134
rect 235794 686000 236414 686898
rect 244794 705798 245414 705830
rect 244794 705562 244826 705798
rect 245062 705562 245146 705798
rect 245382 705562 245414 705798
rect 244794 705478 245414 705562
rect 244794 705242 244826 705478
rect 245062 705242 245146 705478
rect 245382 705242 245414 705478
rect 244794 696454 245414 705242
rect 244794 696218 244826 696454
rect 245062 696218 245146 696454
rect 245382 696218 245414 696454
rect 244794 696134 245414 696218
rect 244794 695898 244826 696134
rect 245062 695898 245146 696134
rect 245382 695898 245414 696134
rect 244794 686000 245414 695898
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 686000 254414 686898
rect 262794 705798 263414 705830
rect 262794 705562 262826 705798
rect 263062 705562 263146 705798
rect 263382 705562 263414 705798
rect 262794 705478 263414 705562
rect 262794 705242 262826 705478
rect 263062 705242 263146 705478
rect 263382 705242 263414 705478
rect 262794 696454 263414 705242
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 686000 263414 695898
rect 271794 704838 272414 705830
rect 271794 704602 271826 704838
rect 272062 704602 272146 704838
rect 272382 704602 272414 704838
rect 271794 704518 272414 704602
rect 271794 704282 271826 704518
rect 272062 704282 272146 704518
rect 272382 704282 272414 704518
rect 271794 687454 272414 704282
rect 271794 687218 271826 687454
rect 272062 687218 272146 687454
rect 272382 687218 272414 687454
rect 271794 687134 272414 687218
rect 271794 686898 271826 687134
rect 272062 686898 272146 687134
rect 272382 686898 272414 687134
rect 271794 686000 272414 686898
rect 280794 705798 281414 705830
rect 280794 705562 280826 705798
rect 281062 705562 281146 705798
rect 281382 705562 281414 705798
rect 280794 705478 281414 705562
rect 280794 705242 280826 705478
rect 281062 705242 281146 705478
rect 281382 705242 281414 705478
rect 280794 696454 281414 705242
rect 280794 696218 280826 696454
rect 281062 696218 281146 696454
rect 281382 696218 281414 696454
rect 280794 696134 281414 696218
rect 280794 695898 280826 696134
rect 281062 695898 281146 696134
rect 281382 695898 281414 696134
rect 280794 686000 281414 695898
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 686000 290414 686898
rect 298794 705798 299414 705830
rect 298794 705562 298826 705798
rect 299062 705562 299146 705798
rect 299382 705562 299414 705798
rect 298794 705478 299414 705562
rect 298794 705242 298826 705478
rect 299062 705242 299146 705478
rect 299382 705242 299414 705478
rect 298794 696454 299414 705242
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 686000 299414 695898
rect 307794 704838 308414 705830
rect 307794 704602 307826 704838
rect 308062 704602 308146 704838
rect 308382 704602 308414 704838
rect 307794 704518 308414 704602
rect 307794 704282 307826 704518
rect 308062 704282 308146 704518
rect 308382 704282 308414 704518
rect 307794 687454 308414 704282
rect 307794 687218 307826 687454
rect 308062 687218 308146 687454
rect 308382 687218 308414 687454
rect 307794 687134 308414 687218
rect 307794 686898 307826 687134
rect 308062 686898 308146 687134
rect 308382 686898 308414 687134
rect 307794 686000 308414 686898
rect 316794 705798 317414 705830
rect 316794 705562 316826 705798
rect 317062 705562 317146 705798
rect 317382 705562 317414 705798
rect 316794 705478 317414 705562
rect 316794 705242 316826 705478
rect 317062 705242 317146 705478
rect 317382 705242 317414 705478
rect 316794 696454 317414 705242
rect 316794 696218 316826 696454
rect 317062 696218 317146 696454
rect 317382 696218 317414 696454
rect 316794 696134 317414 696218
rect 316794 695898 316826 696134
rect 317062 695898 317146 696134
rect 317382 695898 317414 696134
rect 316794 686000 317414 695898
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 686000 326414 686898
rect 334794 705798 335414 705830
rect 334794 705562 334826 705798
rect 335062 705562 335146 705798
rect 335382 705562 335414 705798
rect 334794 705478 335414 705562
rect 334794 705242 334826 705478
rect 335062 705242 335146 705478
rect 335382 705242 335414 705478
rect 334794 696454 335414 705242
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 686000 335414 695898
rect 343794 704838 344414 705830
rect 343794 704602 343826 704838
rect 344062 704602 344146 704838
rect 344382 704602 344414 704838
rect 343794 704518 344414 704602
rect 343794 704282 343826 704518
rect 344062 704282 344146 704518
rect 344382 704282 344414 704518
rect 343794 687454 344414 704282
rect 343794 687218 343826 687454
rect 344062 687218 344146 687454
rect 344382 687218 344414 687454
rect 343794 687134 344414 687218
rect 343794 686898 343826 687134
rect 344062 686898 344146 687134
rect 344382 686898 344414 687134
rect 343794 686000 344414 686898
rect 352794 705798 353414 705830
rect 352794 705562 352826 705798
rect 353062 705562 353146 705798
rect 353382 705562 353414 705798
rect 352794 705478 353414 705562
rect 352794 705242 352826 705478
rect 353062 705242 353146 705478
rect 353382 705242 353414 705478
rect 352794 696454 353414 705242
rect 352794 696218 352826 696454
rect 353062 696218 353146 696454
rect 353382 696218 353414 696454
rect 352794 696134 353414 696218
rect 352794 695898 352826 696134
rect 353062 695898 353146 696134
rect 353382 695898 353414 696134
rect 352794 686000 353414 695898
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 686000 362414 686898
rect 370794 705798 371414 705830
rect 370794 705562 370826 705798
rect 371062 705562 371146 705798
rect 371382 705562 371414 705798
rect 370794 705478 371414 705562
rect 370794 705242 370826 705478
rect 371062 705242 371146 705478
rect 371382 705242 371414 705478
rect 370794 696454 371414 705242
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 686000 371414 695898
rect 379794 704838 380414 705830
rect 379794 704602 379826 704838
rect 380062 704602 380146 704838
rect 380382 704602 380414 704838
rect 379794 704518 380414 704602
rect 379794 704282 379826 704518
rect 380062 704282 380146 704518
rect 380382 704282 380414 704518
rect 379794 687454 380414 704282
rect 379794 687218 379826 687454
rect 380062 687218 380146 687454
rect 380382 687218 380414 687454
rect 379794 687134 380414 687218
rect 379794 686898 379826 687134
rect 380062 686898 380146 687134
rect 380382 686898 380414 687134
rect 379794 686000 380414 686898
rect 388794 705798 389414 705830
rect 388794 705562 388826 705798
rect 389062 705562 389146 705798
rect 389382 705562 389414 705798
rect 388794 705478 389414 705562
rect 388794 705242 388826 705478
rect 389062 705242 389146 705478
rect 389382 705242 389414 705478
rect 388794 696454 389414 705242
rect 388794 696218 388826 696454
rect 389062 696218 389146 696454
rect 389382 696218 389414 696454
rect 388794 696134 389414 696218
rect 388794 695898 388826 696134
rect 389062 695898 389146 696134
rect 389382 695898 389414 696134
rect 388794 686000 389414 695898
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 686000 398414 686898
rect 406794 705798 407414 705830
rect 406794 705562 406826 705798
rect 407062 705562 407146 705798
rect 407382 705562 407414 705798
rect 406794 705478 407414 705562
rect 406794 705242 406826 705478
rect 407062 705242 407146 705478
rect 407382 705242 407414 705478
rect 406794 696454 407414 705242
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 686000 407414 695898
rect 415794 704838 416414 705830
rect 415794 704602 415826 704838
rect 416062 704602 416146 704838
rect 416382 704602 416414 704838
rect 415794 704518 416414 704602
rect 415794 704282 415826 704518
rect 416062 704282 416146 704518
rect 416382 704282 416414 704518
rect 415794 687454 416414 704282
rect 415794 687218 415826 687454
rect 416062 687218 416146 687454
rect 416382 687218 416414 687454
rect 415794 687134 416414 687218
rect 415794 686898 415826 687134
rect 416062 686898 416146 687134
rect 416382 686898 416414 687134
rect 415794 686000 416414 686898
rect 424794 705798 425414 705830
rect 424794 705562 424826 705798
rect 425062 705562 425146 705798
rect 425382 705562 425414 705798
rect 424794 705478 425414 705562
rect 424794 705242 424826 705478
rect 425062 705242 425146 705478
rect 425382 705242 425414 705478
rect 424794 696454 425414 705242
rect 424794 696218 424826 696454
rect 425062 696218 425146 696454
rect 425382 696218 425414 696454
rect 424794 696134 425414 696218
rect 424794 695898 424826 696134
rect 425062 695898 425146 696134
rect 425382 695898 425414 696134
rect 424794 686000 425414 695898
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 686000 434414 686898
rect 442794 705798 443414 705830
rect 442794 705562 442826 705798
rect 443062 705562 443146 705798
rect 443382 705562 443414 705798
rect 442794 705478 443414 705562
rect 442794 705242 442826 705478
rect 443062 705242 443146 705478
rect 443382 705242 443414 705478
rect 442794 696454 443414 705242
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 686000 443414 695898
rect 451794 704838 452414 705830
rect 451794 704602 451826 704838
rect 452062 704602 452146 704838
rect 452382 704602 452414 704838
rect 451794 704518 452414 704602
rect 451794 704282 451826 704518
rect 452062 704282 452146 704518
rect 452382 704282 452414 704518
rect 451794 687454 452414 704282
rect 451794 687218 451826 687454
rect 452062 687218 452146 687454
rect 452382 687218 452414 687454
rect 451794 687134 452414 687218
rect 451794 686898 451826 687134
rect 452062 686898 452146 687134
rect 452382 686898 452414 687134
rect 451794 686000 452414 686898
rect 460794 705798 461414 705830
rect 460794 705562 460826 705798
rect 461062 705562 461146 705798
rect 461382 705562 461414 705798
rect 460794 705478 461414 705562
rect 460794 705242 460826 705478
rect 461062 705242 461146 705478
rect 461382 705242 461414 705478
rect 460794 696454 461414 705242
rect 460794 696218 460826 696454
rect 461062 696218 461146 696454
rect 461382 696218 461414 696454
rect 460794 696134 461414 696218
rect 460794 695898 460826 696134
rect 461062 695898 461146 696134
rect 461382 695898 461414 696134
rect 460794 686000 461414 695898
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 686000 470414 686898
rect 478794 705798 479414 705830
rect 478794 705562 478826 705798
rect 479062 705562 479146 705798
rect 479382 705562 479414 705798
rect 478794 705478 479414 705562
rect 478794 705242 478826 705478
rect 479062 705242 479146 705478
rect 479382 705242 479414 705478
rect 478794 696454 479414 705242
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 686000 479414 695898
rect 487794 704838 488414 705830
rect 487794 704602 487826 704838
rect 488062 704602 488146 704838
rect 488382 704602 488414 704838
rect 487794 704518 488414 704602
rect 487794 704282 487826 704518
rect 488062 704282 488146 704518
rect 488382 704282 488414 704518
rect 487794 687454 488414 704282
rect 487794 687218 487826 687454
rect 488062 687218 488146 687454
rect 488382 687218 488414 687454
rect 487794 687134 488414 687218
rect 487794 686898 487826 687134
rect 488062 686898 488146 687134
rect 488382 686898 488414 687134
rect 487794 686000 488414 686898
rect 496794 705798 497414 705830
rect 496794 705562 496826 705798
rect 497062 705562 497146 705798
rect 497382 705562 497414 705798
rect 496794 705478 497414 705562
rect 496794 705242 496826 705478
rect 497062 705242 497146 705478
rect 497382 705242 497414 705478
rect 496794 696454 497414 705242
rect 496794 696218 496826 696454
rect 497062 696218 497146 696454
rect 497382 696218 497414 696454
rect 496794 696134 497414 696218
rect 496794 695898 496826 696134
rect 497062 695898 497146 696134
rect 497382 695898 497414 696134
rect 496794 686000 497414 695898
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 686000 506414 686898
rect 514794 705798 515414 705830
rect 514794 705562 514826 705798
rect 515062 705562 515146 705798
rect 515382 705562 515414 705798
rect 514794 705478 515414 705562
rect 514794 705242 514826 705478
rect 515062 705242 515146 705478
rect 515382 705242 515414 705478
rect 514794 696454 515414 705242
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 686000 515414 695898
rect 523794 704838 524414 705830
rect 523794 704602 523826 704838
rect 524062 704602 524146 704838
rect 524382 704602 524414 704838
rect 523794 704518 524414 704602
rect 523794 704282 523826 704518
rect 524062 704282 524146 704518
rect 524382 704282 524414 704518
rect 523794 687454 524414 704282
rect 523794 687218 523826 687454
rect 524062 687218 524146 687454
rect 524382 687218 524414 687454
rect 523794 687134 524414 687218
rect 523794 686898 523826 687134
rect 524062 686898 524146 687134
rect 524382 686898 524414 687134
rect 523794 686000 524414 686898
rect 532794 705798 533414 705830
rect 532794 705562 532826 705798
rect 533062 705562 533146 705798
rect 533382 705562 533414 705798
rect 532794 705478 533414 705562
rect 532794 705242 532826 705478
rect 533062 705242 533146 705478
rect 533382 705242 533414 705478
rect 532794 696454 533414 705242
rect 532794 696218 532826 696454
rect 533062 696218 533146 696454
rect 533382 696218 533414 696454
rect 532794 696134 533414 696218
rect 532794 695898 532826 696134
rect 533062 695898 533146 696134
rect 533382 695898 533414 696134
rect 532794 686000 533414 695898
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 686000 542414 686898
rect 550794 705798 551414 705830
rect 550794 705562 550826 705798
rect 551062 705562 551146 705798
rect 551382 705562 551414 705798
rect 550794 705478 551414 705562
rect 550794 705242 550826 705478
rect 551062 705242 551146 705478
rect 551382 705242 551414 705478
rect 550794 696454 551414 705242
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 686000 551414 695898
rect 559794 704838 560414 705830
rect 559794 704602 559826 704838
rect 560062 704602 560146 704838
rect 560382 704602 560414 704838
rect 559794 704518 560414 704602
rect 559794 704282 559826 704518
rect 560062 704282 560146 704518
rect 560382 704282 560414 704518
rect 559794 687454 560414 704282
rect 559794 687218 559826 687454
rect 560062 687218 560146 687454
rect 560382 687218 560414 687454
rect 559794 687134 560414 687218
rect 559794 686898 559826 687134
rect 560062 686898 560146 687134
rect 560382 686898 560414 687134
rect 10794 678218 10826 678454
rect 11062 678218 11146 678454
rect 11382 678218 11414 678454
rect 10794 678134 11414 678218
rect 10794 677898 10826 678134
rect 11062 677898 11146 678134
rect 11382 677898 11414 678134
rect 10794 660454 11414 677898
rect 22874 678454 23194 678486
rect 22874 678218 22916 678454
rect 23152 678218 23194 678454
rect 22874 678134 23194 678218
rect 22874 677898 22916 678134
rect 23152 677898 23194 678134
rect 22874 677866 23194 677898
rect 28805 678454 29125 678486
rect 28805 678218 28847 678454
rect 29083 678218 29125 678454
rect 28805 678134 29125 678218
rect 28805 677898 28847 678134
rect 29083 677898 29125 678134
rect 28805 677866 29125 677898
rect 49874 678454 50194 678486
rect 49874 678218 49916 678454
rect 50152 678218 50194 678454
rect 49874 678134 50194 678218
rect 49874 677898 49916 678134
rect 50152 677898 50194 678134
rect 49874 677866 50194 677898
rect 55805 678454 56125 678486
rect 55805 678218 55847 678454
rect 56083 678218 56125 678454
rect 55805 678134 56125 678218
rect 55805 677898 55847 678134
rect 56083 677898 56125 678134
rect 55805 677866 56125 677898
rect 76874 678454 77194 678486
rect 76874 678218 76916 678454
rect 77152 678218 77194 678454
rect 76874 678134 77194 678218
rect 76874 677898 76916 678134
rect 77152 677898 77194 678134
rect 76874 677866 77194 677898
rect 82805 678454 83125 678486
rect 82805 678218 82847 678454
rect 83083 678218 83125 678454
rect 82805 678134 83125 678218
rect 82805 677898 82847 678134
rect 83083 677898 83125 678134
rect 82805 677866 83125 677898
rect 103874 678454 104194 678486
rect 103874 678218 103916 678454
rect 104152 678218 104194 678454
rect 103874 678134 104194 678218
rect 103874 677898 103916 678134
rect 104152 677898 104194 678134
rect 103874 677866 104194 677898
rect 109805 678454 110125 678486
rect 109805 678218 109847 678454
rect 110083 678218 110125 678454
rect 109805 678134 110125 678218
rect 109805 677898 109847 678134
rect 110083 677898 110125 678134
rect 109805 677866 110125 677898
rect 130874 678454 131194 678486
rect 130874 678218 130916 678454
rect 131152 678218 131194 678454
rect 130874 678134 131194 678218
rect 130874 677898 130916 678134
rect 131152 677898 131194 678134
rect 130874 677866 131194 677898
rect 136805 678454 137125 678486
rect 136805 678218 136847 678454
rect 137083 678218 137125 678454
rect 136805 678134 137125 678218
rect 136805 677898 136847 678134
rect 137083 677898 137125 678134
rect 136805 677866 137125 677898
rect 157874 678454 158194 678486
rect 157874 678218 157916 678454
rect 158152 678218 158194 678454
rect 157874 678134 158194 678218
rect 157874 677898 157916 678134
rect 158152 677898 158194 678134
rect 157874 677866 158194 677898
rect 163805 678454 164125 678486
rect 163805 678218 163847 678454
rect 164083 678218 164125 678454
rect 163805 678134 164125 678218
rect 163805 677898 163847 678134
rect 164083 677898 164125 678134
rect 163805 677866 164125 677898
rect 184874 678454 185194 678486
rect 184874 678218 184916 678454
rect 185152 678218 185194 678454
rect 184874 678134 185194 678218
rect 184874 677898 184916 678134
rect 185152 677898 185194 678134
rect 184874 677866 185194 677898
rect 190805 678454 191125 678486
rect 190805 678218 190847 678454
rect 191083 678218 191125 678454
rect 190805 678134 191125 678218
rect 190805 677898 190847 678134
rect 191083 677898 191125 678134
rect 190805 677866 191125 677898
rect 211874 678454 212194 678486
rect 211874 678218 211916 678454
rect 212152 678218 212194 678454
rect 211874 678134 212194 678218
rect 211874 677898 211916 678134
rect 212152 677898 212194 678134
rect 211874 677866 212194 677898
rect 217805 678454 218125 678486
rect 217805 678218 217847 678454
rect 218083 678218 218125 678454
rect 217805 678134 218125 678218
rect 217805 677898 217847 678134
rect 218083 677898 218125 678134
rect 217805 677866 218125 677898
rect 238874 678454 239194 678486
rect 238874 678218 238916 678454
rect 239152 678218 239194 678454
rect 238874 678134 239194 678218
rect 238874 677898 238916 678134
rect 239152 677898 239194 678134
rect 238874 677866 239194 677898
rect 244805 678454 245125 678486
rect 244805 678218 244847 678454
rect 245083 678218 245125 678454
rect 244805 678134 245125 678218
rect 244805 677898 244847 678134
rect 245083 677898 245125 678134
rect 244805 677866 245125 677898
rect 265874 678454 266194 678486
rect 265874 678218 265916 678454
rect 266152 678218 266194 678454
rect 265874 678134 266194 678218
rect 265874 677898 265916 678134
rect 266152 677898 266194 678134
rect 265874 677866 266194 677898
rect 271805 678454 272125 678486
rect 271805 678218 271847 678454
rect 272083 678218 272125 678454
rect 271805 678134 272125 678218
rect 271805 677898 271847 678134
rect 272083 677898 272125 678134
rect 271805 677866 272125 677898
rect 292874 678454 293194 678486
rect 292874 678218 292916 678454
rect 293152 678218 293194 678454
rect 292874 678134 293194 678218
rect 292874 677898 292916 678134
rect 293152 677898 293194 678134
rect 292874 677866 293194 677898
rect 298805 678454 299125 678486
rect 298805 678218 298847 678454
rect 299083 678218 299125 678454
rect 298805 678134 299125 678218
rect 298805 677898 298847 678134
rect 299083 677898 299125 678134
rect 298805 677866 299125 677898
rect 319874 678454 320194 678486
rect 319874 678218 319916 678454
rect 320152 678218 320194 678454
rect 319874 678134 320194 678218
rect 319874 677898 319916 678134
rect 320152 677898 320194 678134
rect 319874 677866 320194 677898
rect 325805 678454 326125 678486
rect 325805 678218 325847 678454
rect 326083 678218 326125 678454
rect 325805 678134 326125 678218
rect 325805 677898 325847 678134
rect 326083 677898 326125 678134
rect 325805 677866 326125 677898
rect 346874 678454 347194 678486
rect 346874 678218 346916 678454
rect 347152 678218 347194 678454
rect 346874 678134 347194 678218
rect 346874 677898 346916 678134
rect 347152 677898 347194 678134
rect 346874 677866 347194 677898
rect 352805 678454 353125 678486
rect 352805 678218 352847 678454
rect 353083 678218 353125 678454
rect 352805 678134 353125 678218
rect 352805 677898 352847 678134
rect 353083 677898 353125 678134
rect 352805 677866 353125 677898
rect 373874 678454 374194 678486
rect 373874 678218 373916 678454
rect 374152 678218 374194 678454
rect 373874 678134 374194 678218
rect 373874 677898 373916 678134
rect 374152 677898 374194 678134
rect 373874 677866 374194 677898
rect 379805 678454 380125 678486
rect 379805 678218 379847 678454
rect 380083 678218 380125 678454
rect 379805 678134 380125 678218
rect 379805 677898 379847 678134
rect 380083 677898 380125 678134
rect 379805 677866 380125 677898
rect 400874 678454 401194 678486
rect 400874 678218 400916 678454
rect 401152 678218 401194 678454
rect 400874 678134 401194 678218
rect 400874 677898 400916 678134
rect 401152 677898 401194 678134
rect 400874 677866 401194 677898
rect 406805 678454 407125 678486
rect 406805 678218 406847 678454
rect 407083 678218 407125 678454
rect 406805 678134 407125 678218
rect 406805 677898 406847 678134
rect 407083 677898 407125 678134
rect 406805 677866 407125 677898
rect 427874 678454 428194 678486
rect 427874 678218 427916 678454
rect 428152 678218 428194 678454
rect 427874 678134 428194 678218
rect 427874 677898 427916 678134
rect 428152 677898 428194 678134
rect 427874 677866 428194 677898
rect 433805 678454 434125 678486
rect 433805 678218 433847 678454
rect 434083 678218 434125 678454
rect 433805 678134 434125 678218
rect 433805 677898 433847 678134
rect 434083 677898 434125 678134
rect 433805 677866 434125 677898
rect 454874 678454 455194 678486
rect 454874 678218 454916 678454
rect 455152 678218 455194 678454
rect 454874 678134 455194 678218
rect 454874 677898 454916 678134
rect 455152 677898 455194 678134
rect 454874 677866 455194 677898
rect 460805 678454 461125 678486
rect 460805 678218 460847 678454
rect 461083 678218 461125 678454
rect 460805 678134 461125 678218
rect 460805 677898 460847 678134
rect 461083 677898 461125 678134
rect 460805 677866 461125 677898
rect 481874 678454 482194 678486
rect 481874 678218 481916 678454
rect 482152 678218 482194 678454
rect 481874 678134 482194 678218
rect 481874 677898 481916 678134
rect 482152 677898 482194 678134
rect 481874 677866 482194 677898
rect 487805 678454 488125 678486
rect 487805 678218 487847 678454
rect 488083 678218 488125 678454
rect 487805 678134 488125 678218
rect 487805 677898 487847 678134
rect 488083 677898 488125 678134
rect 487805 677866 488125 677898
rect 508874 678454 509194 678486
rect 508874 678218 508916 678454
rect 509152 678218 509194 678454
rect 508874 678134 509194 678218
rect 508874 677898 508916 678134
rect 509152 677898 509194 678134
rect 508874 677866 509194 677898
rect 514805 678454 515125 678486
rect 514805 678218 514847 678454
rect 515083 678218 515125 678454
rect 514805 678134 515125 678218
rect 514805 677898 514847 678134
rect 515083 677898 515125 678134
rect 514805 677866 515125 677898
rect 535874 678454 536194 678486
rect 535874 678218 535916 678454
rect 536152 678218 536194 678454
rect 535874 678134 536194 678218
rect 535874 677898 535916 678134
rect 536152 677898 536194 678134
rect 535874 677866 536194 677898
rect 541805 678454 542125 678486
rect 541805 678218 541847 678454
rect 542083 678218 542125 678454
rect 541805 678134 542125 678218
rect 541805 677898 541847 678134
rect 542083 677898 542125 678134
rect 541805 677866 542125 677898
rect 19910 669454 20230 669486
rect 19910 669218 19952 669454
rect 20188 669218 20230 669454
rect 19910 669134 20230 669218
rect 19910 668898 19952 669134
rect 20188 668898 20230 669134
rect 19910 668866 20230 668898
rect 25840 669454 26160 669486
rect 25840 669218 25882 669454
rect 26118 669218 26160 669454
rect 25840 669134 26160 669218
rect 25840 668898 25882 669134
rect 26118 668898 26160 669134
rect 25840 668866 26160 668898
rect 31771 669454 32091 669486
rect 31771 669218 31813 669454
rect 32049 669218 32091 669454
rect 31771 669134 32091 669218
rect 31771 668898 31813 669134
rect 32049 668898 32091 669134
rect 31771 668866 32091 668898
rect 46910 669454 47230 669486
rect 46910 669218 46952 669454
rect 47188 669218 47230 669454
rect 46910 669134 47230 669218
rect 46910 668898 46952 669134
rect 47188 668898 47230 669134
rect 46910 668866 47230 668898
rect 52840 669454 53160 669486
rect 52840 669218 52882 669454
rect 53118 669218 53160 669454
rect 52840 669134 53160 669218
rect 52840 668898 52882 669134
rect 53118 668898 53160 669134
rect 52840 668866 53160 668898
rect 58771 669454 59091 669486
rect 58771 669218 58813 669454
rect 59049 669218 59091 669454
rect 58771 669134 59091 669218
rect 58771 668898 58813 669134
rect 59049 668898 59091 669134
rect 58771 668866 59091 668898
rect 73910 669454 74230 669486
rect 73910 669218 73952 669454
rect 74188 669218 74230 669454
rect 73910 669134 74230 669218
rect 73910 668898 73952 669134
rect 74188 668898 74230 669134
rect 73910 668866 74230 668898
rect 79840 669454 80160 669486
rect 79840 669218 79882 669454
rect 80118 669218 80160 669454
rect 79840 669134 80160 669218
rect 79840 668898 79882 669134
rect 80118 668898 80160 669134
rect 79840 668866 80160 668898
rect 85771 669454 86091 669486
rect 85771 669218 85813 669454
rect 86049 669218 86091 669454
rect 85771 669134 86091 669218
rect 85771 668898 85813 669134
rect 86049 668898 86091 669134
rect 85771 668866 86091 668898
rect 100910 669454 101230 669486
rect 100910 669218 100952 669454
rect 101188 669218 101230 669454
rect 100910 669134 101230 669218
rect 100910 668898 100952 669134
rect 101188 668898 101230 669134
rect 100910 668866 101230 668898
rect 106840 669454 107160 669486
rect 106840 669218 106882 669454
rect 107118 669218 107160 669454
rect 106840 669134 107160 669218
rect 106840 668898 106882 669134
rect 107118 668898 107160 669134
rect 106840 668866 107160 668898
rect 112771 669454 113091 669486
rect 112771 669218 112813 669454
rect 113049 669218 113091 669454
rect 112771 669134 113091 669218
rect 112771 668898 112813 669134
rect 113049 668898 113091 669134
rect 112771 668866 113091 668898
rect 127910 669454 128230 669486
rect 127910 669218 127952 669454
rect 128188 669218 128230 669454
rect 127910 669134 128230 669218
rect 127910 668898 127952 669134
rect 128188 668898 128230 669134
rect 127910 668866 128230 668898
rect 133840 669454 134160 669486
rect 133840 669218 133882 669454
rect 134118 669218 134160 669454
rect 133840 669134 134160 669218
rect 133840 668898 133882 669134
rect 134118 668898 134160 669134
rect 133840 668866 134160 668898
rect 139771 669454 140091 669486
rect 139771 669218 139813 669454
rect 140049 669218 140091 669454
rect 139771 669134 140091 669218
rect 139771 668898 139813 669134
rect 140049 668898 140091 669134
rect 139771 668866 140091 668898
rect 154910 669454 155230 669486
rect 154910 669218 154952 669454
rect 155188 669218 155230 669454
rect 154910 669134 155230 669218
rect 154910 668898 154952 669134
rect 155188 668898 155230 669134
rect 154910 668866 155230 668898
rect 160840 669454 161160 669486
rect 160840 669218 160882 669454
rect 161118 669218 161160 669454
rect 160840 669134 161160 669218
rect 160840 668898 160882 669134
rect 161118 668898 161160 669134
rect 160840 668866 161160 668898
rect 166771 669454 167091 669486
rect 166771 669218 166813 669454
rect 167049 669218 167091 669454
rect 166771 669134 167091 669218
rect 166771 668898 166813 669134
rect 167049 668898 167091 669134
rect 166771 668866 167091 668898
rect 181910 669454 182230 669486
rect 181910 669218 181952 669454
rect 182188 669218 182230 669454
rect 181910 669134 182230 669218
rect 181910 668898 181952 669134
rect 182188 668898 182230 669134
rect 181910 668866 182230 668898
rect 187840 669454 188160 669486
rect 187840 669218 187882 669454
rect 188118 669218 188160 669454
rect 187840 669134 188160 669218
rect 187840 668898 187882 669134
rect 188118 668898 188160 669134
rect 187840 668866 188160 668898
rect 193771 669454 194091 669486
rect 193771 669218 193813 669454
rect 194049 669218 194091 669454
rect 193771 669134 194091 669218
rect 193771 668898 193813 669134
rect 194049 668898 194091 669134
rect 193771 668866 194091 668898
rect 208910 669454 209230 669486
rect 208910 669218 208952 669454
rect 209188 669218 209230 669454
rect 208910 669134 209230 669218
rect 208910 668898 208952 669134
rect 209188 668898 209230 669134
rect 208910 668866 209230 668898
rect 214840 669454 215160 669486
rect 214840 669218 214882 669454
rect 215118 669218 215160 669454
rect 214840 669134 215160 669218
rect 214840 668898 214882 669134
rect 215118 668898 215160 669134
rect 214840 668866 215160 668898
rect 220771 669454 221091 669486
rect 220771 669218 220813 669454
rect 221049 669218 221091 669454
rect 220771 669134 221091 669218
rect 220771 668898 220813 669134
rect 221049 668898 221091 669134
rect 220771 668866 221091 668898
rect 235910 669454 236230 669486
rect 235910 669218 235952 669454
rect 236188 669218 236230 669454
rect 235910 669134 236230 669218
rect 235910 668898 235952 669134
rect 236188 668898 236230 669134
rect 235910 668866 236230 668898
rect 241840 669454 242160 669486
rect 241840 669218 241882 669454
rect 242118 669218 242160 669454
rect 241840 669134 242160 669218
rect 241840 668898 241882 669134
rect 242118 668898 242160 669134
rect 241840 668866 242160 668898
rect 247771 669454 248091 669486
rect 247771 669218 247813 669454
rect 248049 669218 248091 669454
rect 247771 669134 248091 669218
rect 247771 668898 247813 669134
rect 248049 668898 248091 669134
rect 247771 668866 248091 668898
rect 262910 669454 263230 669486
rect 262910 669218 262952 669454
rect 263188 669218 263230 669454
rect 262910 669134 263230 669218
rect 262910 668898 262952 669134
rect 263188 668898 263230 669134
rect 262910 668866 263230 668898
rect 268840 669454 269160 669486
rect 268840 669218 268882 669454
rect 269118 669218 269160 669454
rect 268840 669134 269160 669218
rect 268840 668898 268882 669134
rect 269118 668898 269160 669134
rect 268840 668866 269160 668898
rect 274771 669454 275091 669486
rect 274771 669218 274813 669454
rect 275049 669218 275091 669454
rect 274771 669134 275091 669218
rect 274771 668898 274813 669134
rect 275049 668898 275091 669134
rect 274771 668866 275091 668898
rect 289910 669454 290230 669486
rect 289910 669218 289952 669454
rect 290188 669218 290230 669454
rect 289910 669134 290230 669218
rect 289910 668898 289952 669134
rect 290188 668898 290230 669134
rect 289910 668866 290230 668898
rect 295840 669454 296160 669486
rect 295840 669218 295882 669454
rect 296118 669218 296160 669454
rect 295840 669134 296160 669218
rect 295840 668898 295882 669134
rect 296118 668898 296160 669134
rect 295840 668866 296160 668898
rect 301771 669454 302091 669486
rect 301771 669218 301813 669454
rect 302049 669218 302091 669454
rect 301771 669134 302091 669218
rect 301771 668898 301813 669134
rect 302049 668898 302091 669134
rect 301771 668866 302091 668898
rect 316910 669454 317230 669486
rect 316910 669218 316952 669454
rect 317188 669218 317230 669454
rect 316910 669134 317230 669218
rect 316910 668898 316952 669134
rect 317188 668898 317230 669134
rect 316910 668866 317230 668898
rect 322840 669454 323160 669486
rect 322840 669218 322882 669454
rect 323118 669218 323160 669454
rect 322840 669134 323160 669218
rect 322840 668898 322882 669134
rect 323118 668898 323160 669134
rect 322840 668866 323160 668898
rect 328771 669454 329091 669486
rect 328771 669218 328813 669454
rect 329049 669218 329091 669454
rect 328771 669134 329091 669218
rect 328771 668898 328813 669134
rect 329049 668898 329091 669134
rect 328771 668866 329091 668898
rect 343910 669454 344230 669486
rect 343910 669218 343952 669454
rect 344188 669218 344230 669454
rect 343910 669134 344230 669218
rect 343910 668898 343952 669134
rect 344188 668898 344230 669134
rect 343910 668866 344230 668898
rect 349840 669454 350160 669486
rect 349840 669218 349882 669454
rect 350118 669218 350160 669454
rect 349840 669134 350160 669218
rect 349840 668898 349882 669134
rect 350118 668898 350160 669134
rect 349840 668866 350160 668898
rect 355771 669454 356091 669486
rect 355771 669218 355813 669454
rect 356049 669218 356091 669454
rect 355771 669134 356091 669218
rect 355771 668898 355813 669134
rect 356049 668898 356091 669134
rect 355771 668866 356091 668898
rect 370910 669454 371230 669486
rect 370910 669218 370952 669454
rect 371188 669218 371230 669454
rect 370910 669134 371230 669218
rect 370910 668898 370952 669134
rect 371188 668898 371230 669134
rect 370910 668866 371230 668898
rect 376840 669454 377160 669486
rect 376840 669218 376882 669454
rect 377118 669218 377160 669454
rect 376840 669134 377160 669218
rect 376840 668898 376882 669134
rect 377118 668898 377160 669134
rect 376840 668866 377160 668898
rect 382771 669454 383091 669486
rect 382771 669218 382813 669454
rect 383049 669218 383091 669454
rect 382771 669134 383091 669218
rect 382771 668898 382813 669134
rect 383049 668898 383091 669134
rect 382771 668866 383091 668898
rect 397910 669454 398230 669486
rect 397910 669218 397952 669454
rect 398188 669218 398230 669454
rect 397910 669134 398230 669218
rect 397910 668898 397952 669134
rect 398188 668898 398230 669134
rect 397910 668866 398230 668898
rect 403840 669454 404160 669486
rect 403840 669218 403882 669454
rect 404118 669218 404160 669454
rect 403840 669134 404160 669218
rect 403840 668898 403882 669134
rect 404118 668898 404160 669134
rect 403840 668866 404160 668898
rect 409771 669454 410091 669486
rect 409771 669218 409813 669454
rect 410049 669218 410091 669454
rect 409771 669134 410091 669218
rect 409771 668898 409813 669134
rect 410049 668898 410091 669134
rect 409771 668866 410091 668898
rect 424910 669454 425230 669486
rect 424910 669218 424952 669454
rect 425188 669218 425230 669454
rect 424910 669134 425230 669218
rect 424910 668898 424952 669134
rect 425188 668898 425230 669134
rect 424910 668866 425230 668898
rect 430840 669454 431160 669486
rect 430840 669218 430882 669454
rect 431118 669218 431160 669454
rect 430840 669134 431160 669218
rect 430840 668898 430882 669134
rect 431118 668898 431160 669134
rect 430840 668866 431160 668898
rect 436771 669454 437091 669486
rect 436771 669218 436813 669454
rect 437049 669218 437091 669454
rect 436771 669134 437091 669218
rect 436771 668898 436813 669134
rect 437049 668898 437091 669134
rect 436771 668866 437091 668898
rect 451910 669454 452230 669486
rect 451910 669218 451952 669454
rect 452188 669218 452230 669454
rect 451910 669134 452230 669218
rect 451910 668898 451952 669134
rect 452188 668898 452230 669134
rect 451910 668866 452230 668898
rect 457840 669454 458160 669486
rect 457840 669218 457882 669454
rect 458118 669218 458160 669454
rect 457840 669134 458160 669218
rect 457840 668898 457882 669134
rect 458118 668898 458160 669134
rect 457840 668866 458160 668898
rect 463771 669454 464091 669486
rect 463771 669218 463813 669454
rect 464049 669218 464091 669454
rect 463771 669134 464091 669218
rect 463771 668898 463813 669134
rect 464049 668898 464091 669134
rect 463771 668866 464091 668898
rect 478910 669454 479230 669486
rect 478910 669218 478952 669454
rect 479188 669218 479230 669454
rect 478910 669134 479230 669218
rect 478910 668898 478952 669134
rect 479188 668898 479230 669134
rect 478910 668866 479230 668898
rect 484840 669454 485160 669486
rect 484840 669218 484882 669454
rect 485118 669218 485160 669454
rect 484840 669134 485160 669218
rect 484840 668898 484882 669134
rect 485118 668898 485160 669134
rect 484840 668866 485160 668898
rect 490771 669454 491091 669486
rect 490771 669218 490813 669454
rect 491049 669218 491091 669454
rect 490771 669134 491091 669218
rect 490771 668898 490813 669134
rect 491049 668898 491091 669134
rect 490771 668866 491091 668898
rect 505910 669454 506230 669486
rect 505910 669218 505952 669454
rect 506188 669218 506230 669454
rect 505910 669134 506230 669218
rect 505910 668898 505952 669134
rect 506188 668898 506230 669134
rect 505910 668866 506230 668898
rect 511840 669454 512160 669486
rect 511840 669218 511882 669454
rect 512118 669218 512160 669454
rect 511840 669134 512160 669218
rect 511840 668898 511882 669134
rect 512118 668898 512160 669134
rect 511840 668866 512160 668898
rect 517771 669454 518091 669486
rect 517771 669218 517813 669454
rect 518049 669218 518091 669454
rect 517771 669134 518091 669218
rect 517771 668898 517813 669134
rect 518049 668898 518091 669134
rect 517771 668866 518091 668898
rect 532910 669454 533230 669486
rect 532910 669218 532952 669454
rect 533188 669218 533230 669454
rect 532910 669134 533230 669218
rect 532910 668898 532952 669134
rect 533188 668898 533230 669134
rect 532910 668866 533230 668898
rect 538840 669454 539160 669486
rect 538840 669218 538882 669454
rect 539118 669218 539160 669454
rect 538840 669134 539160 669218
rect 538840 668898 538882 669134
rect 539118 668898 539160 669134
rect 538840 668866 539160 668898
rect 544771 669454 545091 669486
rect 544771 669218 544813 669454
rect 545049 669218 545091 669454
rect 544771 669134 545091 669218
rect 544771 668898 544813 669134
rect 545049 668898 545091 669134
rect 544771 668866 545091 668898
rect 559794 669454 560414 686898
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 642454 11414 659898
rect 19794 661394 20414 662000
rect 19794 661158 19826 661394
rect 20062 661158 20146 661394
rect 20382 661158 20414 661394
rect 19794 661074 20414 661158
rect 19794 660838 19826 661074
rect 20062 660838 20146 661074
rect 20382 660838 20414 661074
rect 19794 659000 20414 660838
rect 28794 660454 29414 662000
rect 28794 660218 28826 660454
rect 29062 660218 29146 660454
rect 29382 660218 29414 660454
rect 28794 660134 29414 660218
rect 28794 659898 28826 660134
rect 29062 659898 29146 660134
rect 29382 659898 29414 660134
rect 28794 659000 29414 659898
rect 37794 661394 38414 662000
rect 37794 661158 37826 661394
rect 38062 661158 38146 661394
rect 38382 661158 38414 661394
rect 37794 661074 38414 661158
rect 37794 660838 37826 661074
rect 38062 660838 38146 661074
rect 38382 660838 38414 661074
rect 37794 659000 38414 660838
rect 46794 660454 47414 662000
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 659000 47414 659898
rect 55794 661394 56414 662000
rect 55794 661158 55826 661394
rect 56062 661158 56146 661394
rect 56382 661158 56414 661394
rect 55794 661074 56414 661158
rect 55794 660838 55826 661074
rect 56062 660838 56146 661074
rect 56382 660838 56414 661074
rect 55794 659000 56414 660838
rect 64794 660454 65414 662000
rect 64794 660218 64826 660454
rect 65062 660218 65146 660454
rect 65382 660218 65414 660454
rect 64794 660134 65414 660218
rect 64794 659898 64826 660134
rect 65062 659898 65146 660134
rect 65382 659898 65414 660134
rect 64794 659000 65414 659898
rect 73794 661394 74414 662000
rect 73794 661158 73826 661394
rect 74062 661158 74146 661394
rect 74382 661158 74414 661394
rect 73794 661074 74414 661158
rect 73794 660838 73826 661074
rect 74062 660838 74146 661074
rect 74382 660838 74414 661074
rect 73794 659000 74414 660838
rect 82794 660454 83414 662000
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 659000 83414 659898
rect 91794 661394 92414 662000
rect 91794 661158 91826 661394
rect 92062 661158 92146 661394
rect 92382 661158 92414 661394
rect 91794 661074 92414 661158
rect 91794 660838 91826 661074
rect 92062 660838 92146 661074
rect 92382 660838 92414 661074
rect 91794 659000 92414 660838
rect 100794 660454 101414 662000
rect 100794 660218 100826 660454
rect 101062 660218 101146 660454
rect 101382 660218 101414 660454
rect 100794 660134 101414 660218
rect 100794 659898 100826 660134
rect 101062 659898 101146 660134
rect 101382 659898 101414 660134
rect 100794 659000 101414 659898
rect 109794 661394 110414 662000
rect 109794 661158 109826 661394
rect 110062 661158 110146 661394
rect 110382 661158 110414 661394
rect 109794 661074 110414 661158
rect 109794 660838 109826 661074
rect 110062 660838 110146 661074
rect 110382 660838 110414 661074
rect 109794 659000 110414 660838
rect 118794 660454 119414 662000
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 659000 119414 659898
rect 127794 661394 128414 662000
rect 127794 661158 127826 661394
rect 128062 661158 128146 661394
rect 128382 661158 128414 661394
rect 127794 661074 128414 661158
rect 127794 660838 127826 661074
rect 128062 660838 128146 661074
rect 128382 660838 128414 661074
rect 127794 659000 128414 660838
rect 136794 660454 137414 662000
rect 136794 660218 136826 660454
rect 137062 660218 137146 660454
rect 137382 660218 137414 660454
rect 136794 660134 137414 660218
rect 136794 659898 136826 660134
rect 137062 659898 137146 660134
rect 137382 659898 137414 660134
rect 136794 659000 137414 659898
rect 145794 661394 146414 662000
rect 145794 661158 145826 661394
rect 146062 661158 146146 661394
rect 146382 661158 146414 661394
rect 145794 661074 146414 661158
rect 145794 660838 145826 661074
rect 146062 660838 146146 661074
rect 146382 660838 146414 661074
rect 145794 659000 146414 660838
rect 154794 660454 155414 662000
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 659000 155414 659898
rect 163794 661394 164414 662000
rect 163794 661158 163826 661394
rect 164062 661158 164146 661394
rect 164382 661158 164414 661394
rect 163794 661074 164414 661158
rect 163794 660838 163826 661074
rect 164062 660838 164146 661074
rect 164382 660838 164414 661074
rect 163794 659000 164414 660838
rect 172794 660454 173414 662000
rect 172794 660218 172826 660454
rect 173062 660218 173146 660454
rect 173382 660218 173414 660454
rect 172794 660134 173414 660218
rect 172794 659898 172826 660134
rect 173062 659898 173146 660134
rect 173382 659898 173414 660134
rect 172794 659000 173414 659898
rect 181794 661394 182414 662000
rect 181794 661158 181826 661394
rect 182062 661158 182146 661394
rect 182382 661158 182414 661394
rect 181794 661074 182414 661158
rect 181794 660838 181826 661074
rect 182062 660838 182146 661074
rect 182382 660838 182414 661074
rect 181794 659000 182414 660838
rect 190794 660454 191414 662000
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 659000 191414 659898
rect 199794 661394 200414 662000
rect 199794 661158 199826 661394
rect 200062 661158 200146 661394
rect 200382 661158 200414 661394
rect 199794 661074 200414 661158
rect 199794 660838 199826 661074
rect 200062 660838 200146 661074
rect 200382 660838 200414 661074
rect 199794 659000 200414 660838
rect 208794 660454 209414 662000
rect 208794 660218 208826 660454
rect 209062 660218 209146 660454
rect 209382 660218 209414 660454
rect 208794 660134 209414 660218
rect 208794 659898 208826 660134
rect 209062 659898 209146 660134
rect 209382 659898 209414 660134
rect 208794 659000 209414 659898
rect 217794 661394 218414 662000
rect 217794 661158 217826 661394
rect 218062 661158 218146 661394
rect 218382 661158 218414 661394
rect 217794 661074 218414 661158
rect 217794 660838 217826 661074
rect 218062 660838 218146 661074
rect 218382 660838 218414 661074
rect 217794 659000 218414 660838
rect 226794 660454 227414 662000
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 659000 227414 659898
rect 235794 661394 236414 662000
rect 235794 661158 235826 661394
rect 236062 661158 236146 661394
rect 236382 661158 236414 661394
rect 235794 661074 236414 661158
rect 235794 660838 235826 661074
rect 236062 660838 236146 661074
rect 236382 660838 236414 661074
rect 235794 659000 236414 660838
rect 244794 660454 245414 662000
rect 244794 660218 244826 660454
rect 245062 660218 245146 660454
rect 245382 660218 245414 660454
rect 244794 660134 245414 660218
rect 244794 659898 244826 660134
rect 245062 659898 245146 660134
rect 245382 659898 245414 660134
rect 244794 659000 245414 659898
rect 253794 661394 254414 662000
rect 253794 661158 253826 661394
rect 254062 661158 254146 661394
rect 254382 661158 254414 661394
rect 253794 661074 254414 661158
rect 253794 660838 253826 661074
rect 254062 660838 254146 661074
rect 254382 660838 254414 661074
rect 253794 659000 254414 660838
rect 262794 660454 263414 662000
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 659000 263414 659898
rect 271794 661394 272414 662000
rect 271794 661158 271826 661394
rect 272062 661158 272146 661394
rect 272382 661158 272414 661394
rect 271794 661074 272414 661158
rect 271794 660838 271826 661074
rect 272062 660838 272146 661074
rect 272382 660838 272414 661074
rect 271794 659000 272414 660838
rect 280794 660454 281414 662000
rect 280794 660218 280826 660454
rect 281062 660218 281146 660454
rect 281382 660218 281414 660454
rect 280794 660134 281414 660218
rect 280794 659898 280826 660134
rect 281062 659898 281146 660134
rect 281382 659898 281414 660134
rect 280794 659000 281414 659898
rect 289794 661394 290414 662000
rect 289794 661158 289826 661394
rect 290062 661158 290146 661394
rect 290382 661158 290414 661394
rect 289794 661074 290414 661158
rect 289794 660838 289826 661074
rect 290062 660838 290146 661074
rect 290382 660838 290414 661074
rect 289794 659000 290414 660838
rect 298794 660454 299414 662000
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 659000 299414 659898
rect 307794 661394 308414 662000
rect 307794 661158 307826 661394
rect 308062 661158 308146 661394
rect 308382 661158 308414 661394
rect 307794 661074 308414 661158
rect 307794 660838 307826 661074
rect 308062 660838 308146 661074
rect 308382 660838 308414 661074
rect 307794 659000 308414 660838
rect 316794 660454 317414 662000
rect 316794 660218 316826 660454
rect 317062 660218 317146 660454
rect 317382 660218 317414 660454
rect 316794 660134 317414 660218
rect 316794 659898 316826 660134
rect 317062 659898 317146 660134
rect 317382 659898 317414 660134
rect 316794 659000 317414 659898
rect 325794 661394 326414 662000
rect 325794 661158 325826 661394
rect 326062 661158 326146 661394
rect 326382 661158 326414 661394
rect 325794 661074 326414 661158
rect 325794 660838 325826 661074
rect 326062 660838 326146 661074
rect 326382 660838 326414 661074
rect 325794 659000 326414 660838
rect 334794 660454 335414 662000
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 659000 335414 659898
rect 343794 661394 344414 662000
rect 343794 661158 343826 661394
rect 344062 661158 344146 661394
rect 344382 661158 344414 661394
rect 343794 661074 344414 661158
rect 343794 660838 343826 661074
rect 344062 660838 344146 661074
rect 344382 660838 344414 661074
rect 343794 659000 344414 660838
rect 352794 660454 353414 662000
rect 352794 660218 352826 660454
rect 353062 660218 353146 660454
rect 353382 660218 353414 660454
rect 352794 660134 353414 660218
rect 352794 659898 352826 660134
rect 353062 659898 353146 660134
rect 353382 659898 353414 660134
rect 352794 659000 353414 659898
rect 361794 661394 362414 662000
rect 361794 661158 361826 661394
rect 362062 661158 362146 661394
rect 362382 661158 362414 661394
rect 361794 661074 362414 661158
rect 361794 660838 361826 661074
rect 362062 660838 362146 661074
rect 362382 660838 362414 661074
rect 361794 659000 362414 660838
rect 370794 660454 371414 662000
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 659000 371414 659898
rect 379794 661394 380414 662000
rect 379794 661158 379826 661394
rect 380062 661158 380146 661394
rect 380382 661158 380414 661394
rect 379794 661074 380414 661158
rect 379794 660838 379826 661074
rect 380062 660838 380146 661074
rect 380382 660838 380414 661074
rect 379794 659000 380414 660838
rect 388794 660454 389414 662000
rect 388794 660218 388826 660454
rect 389062 660218 389146 660454
rect 389382 660218 389414 660454
rect 388794 660134 389414 660218
rect 388794 659898 388826 660134
rect 389062 659898 389146 660134
rect 389382 659898 389414 660134
rect 388794 659000 389414 659898
rect 397794 661394 398414 662000
rect 397794 661158 397826 661394
rect 398062 661158 398146 661394
rect 398382 661158 398414 661394
rect 397794 661074 398414 661158
rect 397794 660838 397826 661074
rect 398062 660838 398146 661074
rect 398382 660838 398414 661074
rect 397794 659000 398414 660838
rect 406794 660454 407414 662000
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 659000 407414 659898
rect 415794 661394 416414 662000
rect 415794 661158 415826 661394
rect 416062 661158 416146 661394
rect 416382 661158 416414 661394
rect 415794 661074 416414 661158
rect 415794 660838 415826 661074
rect 416062 660838 416146 661074
rect 416382 660838 416414 661074
rect 415794 659000 416414 660838
rect 424794 660454 425414 662000
rect 424794 660218 424826 660454
rect 425062 660218 425146 660454
rect 425382 660218 425414 660454
rect 424794 660134 425414 660218
rect 424794 659898 424826 660134
rect 425062 659898 425146 660134
rect 425382 659898 425414 660134
rect 424794 659000 425414 659898
rect 433794 661394 434414 662000
rect 433794 661158 433826 661394
rect 434062 661158 434146 661394
rect 434382 661158 434414 661394
rect 433794 661074 434414 661158
rect 433794 660838 433826 661074
rect 434062 660838 434146 661074
rect 434382 660838 434414 661074
rect 433794 659000 434414 660838
rect 442794 660454 443414 662000
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 659000 443414 659898
rect 451794 661394 452414 662000
rect 451794 661158 451826 661394
rect 452062 661158 452146 661394
rect 452382 661158 452414 661394
rect 451794 661074 452414 661158
rect 451794 660838 451826 661074
rect 452062 660838 452146 661074
rect 452382 660838 452414 661074
rect 451794 659000 452414 660838
rect 460794 660454 461414 662000
rect 460794 660218 460826 660454
rect 461062 660218 461146 660454
rect 461382 660218 461414 660454
rect 460794 660134 461414 660218
rect 460794 659898 460826 660134
rect 461062 659898 461146 660134
rect 461382 659898 461414 660134
rect 460794 659000 461414 659898
rect 469794 661394 470414 662000
rect 469794 661158 469826 661394
rect 470062 661158 470146 661394
rect 470382 661158 470414 661394
rect 469794 661074 470414 661158
rect 469794 660838 469826 661074
rect 470062 660838 470146 661074
rect 470382 660838 470414 661074
rect 469794 659000 470414 660838
rect 478794 660454 479414 662000
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 659000 479414 659898
rect 487794 661394 488414 662000
rect 487794 661158 487826 661394
rect 488062 661158 488146 661394
rect 488382 661158 488414 661394
rect 487794 661074 488414 661158
rect 487794 660838 487826 661074
rect 488062 660838 488146 661074
rect 488382 660838 488414 661074
rect 487794 659000 488414 660838
rect 496794 660454 497414 662000
rect 496794 660218 496826 660454
rect 497062 660218 497146 660454
rect 497382 660218 497414 660454
rect 496794 660134 497414 660218
rect 496794 659898 496826 660134
rect 497062 659898 497146 660134
rect 497382 659898 497414 660134
rect 496794 659000 497414 659898
rect 505794 661394 506414 662000
rect 505794 661158 505826 661394
rect 506062 661158 506146 661394
rect 506382 661158 506414 661394
rect 505794 661074 506414 661158
rect 505794 660838 505826 661074
rect 506062 660838 506146 661074
rect 506382 660838 506414 661074
rect 505794 659000 506414 660838
rect 514794 660454 515414 662000
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 659000 515414 659898
rect 523794 661394 524414 662000
rect 523794 661158 523826 661394
rect 524062 661158 524146 661394
rect 524382 661158 524414 661394
rect 523794 661074 524414 661158
rect 523794 660838 523826 661074
rect 524062 660838 524146 661074
rect 524382 660838 524414 661074
rect 523794 659000 524414 660838
rect 532794 660454 533414 662000
rect 532794 660218 532826 660454
rect 533062 660218 533146 660454
rect 533382 660218 533414 660454
rect 532794 660134 533414 660218
rect 532794 659898 532826 660134
rect 533062 659898 533146 660134
rect 533382 659898 533414 660134
rect 532794 659000 533414 659898
rect 541794 661394 542414 662000
rect 541794 661158 541826 661394
rect 542062 661158 542146 661394
rect 542382 661158 542414 661394
rect 541794 661074 542414 661158
rect 541794 660838 541826 661074
rect 542062 660838 542146 661074
rect 542382 660838 542414 661074
rect 541794 659000 542414 660838
rect 550794 660454 551414 662000
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 659000 551414 659898
rect 19910 651454 20230 651486
rect 19910 651218 19952 651454
rect 20188 651218 20230 651454
rect 19910 651134 20230 651218
rect 19910 650898 19952 651134
rect 20188 650898 20230 651134
rect 19910 650866 20230 650898
rect 25840 651454 26160 651486
rect 25840 651218 25882 651454
rect 26118 651218 26160 651454
rect 25840 651134 26160 651218
rect 25840 650898 25882 651134
rect 26118 650898 26160 651134
rect 25840 650866 26160 650898
rect 31771 651454 32091 651486
rect 31771 651218 31813 651454
rect 32049 651218 32091 651454
rect 31771 651134 32091 651218
rect 31771 650898 31813 651134
rect 32049 650898 32091 651134
rect 31771 650866 32091 650898
rect 46910 651454 47230 651486
rect 46910 651218 46952 651454
rect 47188 651218 47230 651454
rect 46910 651134 47230 651218
rect 46910 650898 46952 651134
rect 47188 650898 47230 651134
rect 46910 650866 47230 650898
rect 52840 651454 53160 651486
rect 52840 651218 52882 651454
rect 53118 651218 53160 651454
rect 52840 651134 53160 651218
rect 52840 650898 52882 651134
rect 53118 650898 53160 651134
rect 52840 650866 53160 650898
rect 58771 651454 59091 651486
rect 58771 651218 58813 651454
rect 59049 651218 59091 651454
rect 58771 651134 59091 651218
rect 58771 650898 58813 651134
rect 59049 650898 59091 651134
rect 58771 650866 59091 650898
rect 73910 651454 74230 651486
rect 73910 651218 73952 651454
rect 74188 651218 74230 651454
rect 73910 651134 74230 651218
rect 73910 650898 73952 651134
rect 74188 650898 74230 651134
rect 73910 650866 74230 650898
rect 79840 651454 80160 651486
rect 79840 651218 79882 651454
rect 80118 651218 80160 651454
rect 79840 651134 80160 651218
rect 79840 650898 79882 651134
rect 80118 650898 80160 651134
rect 79840 650866 80160 650898
rect 85771 651454 86091 651486
rect 85771 651218 85813 651454
rect 86049 651218 86091 651454
rect 85771 651134 86091 651218
rect 85771 650898 85813 651134
rect 86049 650898 86091 651134
rect 85771 650866 86091 650898
rect 100910 651454 101230 651486
rect 100910 651218 100952 651454
rect 101188 651218 101230 651454
rect 100910 651134 101230 651218
rect 100910 650898 100952 651134
rect 101188 650898 101230 651134
rect 100910 650866 101230 650898
rect 106840 651454 107160 651486
rect 106840 651218 106882 651454
rect 107118 651218 107160 651454
rect 106840 651134 107160 651218
rect 106840 650898 106882 651134
rect 107118 650898 107160 651134
rect 106840 650866 107160 650898
rect 112771 651454 113091 651486
rect 112771 651218 112813 651454
rect 113049 651218 113091 651454
rect 112771 651134 113091 651218
rect 112771 650898 112813 651134
rect 113049 650898 113091 651134
rect 112771 650866 113091 650898
rect 127910 651454 128230 651486
rect 127910 651218 127952 651454
rect 128188 651218 128230 651454
rect 127910 651134 128230 651218
rect 127910 650898 127952 651134
rect 128188 650898 128230 651134
rect 127910 650866 128230 650898
rect 133840 651454 134160 651486
rect 133840 651218 133882 651454
rect 134118 651218 134160 651454
rect 133840 651134 134160 651218
rect 133840 650898 133882 651134
rect 134118 650898 134160 651134
rect 133840 650866 134160 650898
rect 139771 651454 140091 651486
rect 139771 651218 139813 651454
rect 140049 651218 140091 651454
rect 139771 651134 140091 651218
rect 139771 650898 139813 651134
rect 140049 650898 140091 651134
rect 139771 650866 140091 650898
rect 154910 651454 155230 651486
rect 154910 651218 154952 651454
rect 155188 651218 155230 651454
rect 154910 651134 155230 651218
rect 154910 650898 154952 651134
rect 155188 650898 155230 651134
rect 154910 650866 155230 650898
rect 160840 651454 161160 651486
rect 160840 651218 160882 651454
rect 161118 651218 161160 651454
rect 160840 651134 161160 651218
rect 160840 650898 160882 651134
rect 161118 650898 161160 651134
rect 160840 650866 161160 650898
rect 166771 651454 167091 651486
rect 166771 651218 166813 651454
rect 167049 651218 167091 651454
rect 166771 651134 167091 651218
rect 166771 650898 166813 651134
rect 167049 650898 167091 651134
rect 166771 650866 167091 650898
rect 181910 651454 182230 651486
rect 181910 651218 181952 651454
rect 182188 651218 182230 651454
rect 181910 651134 182230 651218
rect 181910 650898 181952 651134
rect 182188 650898 182230 651134
rect 181910 650866 182230 650898
rect 187840 651454 188160 651486
rect 187840 651218 187882 651454
rect 188118 651218 188160 651454
rect 187840 651134 188160 651218
rect 187840 650898 187882 651134
rect 188118 650898 188160 651134
rect 187840 650866 188160 650898
rect 193771 651454 194091 651486
rect 193771 651218 193813 651454
rect 194049 651218 194091 651454
rect 193771 651134 194091 651218
rect 193771 650898 193813 651134
rect 194049 650898 194091 651134
rect 193771 650866 194091 650898
rect 208910 651454 209230 651486
rect 208910 651218 208952 651454
rect 209188 651218 209230 651454
rect 208910 651134 209230 651218
rect 208910 650898 208952 651134
rect 209188 650898 209230 651134
rect 208910 650866 209230 650898
rect 214840 651454 215160 651486
rect 214840 651218 214882 651454
rect 215118 651218 215160 651454
rect 214840 651134 215160 651218
rect 214840 650898 214882 651134
rect 215118 650898 215160 651134
rect 214840 650866 215160 650898
rect 220771 651454 221091 651486
rect 220771 651218 220813 651454
rect 221049 651218 221091 651454
rect 220771 651134 221091 651218
rect 220771 650898 220813 651134
rect 221049 650898 221091 651134
rect 220771 650866 221091 650898
rect 235910 651454 236230 651486
rect 235910 651218 235952 651454
rect 236188 651218 236230 651454
rect 235910 651134 236230 651218
rect 235910 650898 235952 651134
rect 236188 650898 236230 651134
rect 235910 650866 236230 650898
rect 241840 651454 242160 651486
rect 241840 651218 241882 651454
rect 242118 651218 242160 651454
rect 241840 651134 242160 651218
rect 241840 650898 241882 651134
rect 242118 650898 242160 651134
rect 241840 650866 242160 650898
rect 247771 651454 248091 651486
rect 247771 651218 247813 651454
rect 248049 651218 248091 651454
rect 247771 651134 248091 651218
rect 247771 650898 247813 651134
rect 248049 650898 248091 651134
rect 247771 650866 248091 650898
rect 262910 651454 263230 651486
rect 262910 651218 262952 651454
rect 263188 651218 263230 651454
rect 262910 651134 263230 651218
rect 262910 650898 262952 651134
rect 263188 650898 263230 651134
rect 262910 650866 263230 650898
rect 268840 651454 269160 651486
rect 268840 651218 268882 651454
rect 269118 651218 269160 651454
rect 268840 651134 269160 651218
rect 268840 650898 268882 651134
rect 269118 650898 269160 651134
rect 268840 650866 269160 650898
rect 274771 651454 275091 651486
rect 274771 651218 274813 651454
rect 275049 651218 275091 651454
rect 274771 651134 275091 651218
rect 274771 650898 274813 651134
rect 275049 650898 275091 651134
rect 274771 650866 275091 650898
rect 289910 651454 290230 651486
rect 289910 651218 289952 651454
rect 290188 651218 290230 651454
rect 289910 651134 290230 651218
rect 289910 650898 289952 651134
rect 290188 650898 290230 651134
rect 289910 650866 290230 650898
rect 295840 651454 296160 651486
rect 295840 651218 295882 651454
rect 296118 651218 296160 651454
rect 295840 651134 296160 651218
rect 295840 650898 295882 651134
rect 296118 650898 296160 651134
rect 295840 650866 296160 650898
rect 301771 651454 302091 651486
rect 301771 651218 301813 651454
rect 302049 651218 302091 651454
rect 301771 651134 302091 651218
rect 301771 650898 301813 651134
rect 302049 650898 302091 651134
rect 301771 650866 302091 650898
rect 316910 651454 317230 651486
rect 316910 651218 316952 651454
rect 317188 651218 317230 651454
rect 316910 651134 317230 651218
rect 316910 650898 316952 651134
rect 317188 650898 317230 651134
rect 316910 650866 317230 650898
rect 322840 651454 323160 651486
rect 322840 651218 322882 651454
rect 323118 651218 323160 651454
rect 322840 651134 323160 651218
rect 322840 650898 322882 651134
rect 323118 650898 323160 651134
rect 322840 650866 323160 650898
rect 328771 651454 329091 651486
rect 328771 651218 328813 651454
rect 329049 651218 329091 651454
rect 328771 651134 329091 651218
rect 328771 650898 328813 651134
rect 329049 650898 329091 651134
rect 328771 650866 329091 650898
rect 343910 651454 344230 651486
rect 343910 651218 343952 651454
rect 344188 651218 344230 651454
rect 343910 651134 344230 651218
rect 343910 650898 343952 651134
rect 344188 650898 344230 651134
rect 343910 650866 344230 650898
rect 349840 651454 350160 651486
rect 349840 651218 349882 651454
rect 350118 651218 350160 651454
rect 349840 651134 350160 651218
rect 349840 650898 349882 651134
rect 350118 650898 350160 651134
rect 349840 650866 350160 650898
rect 355771 651454 356091 651486
rect 355771 651218 355813 651454
rect 356049 651218 356091 651454
rect 355771 651134 356091 651218
rect 355771 650898 355813 651134
rect 356049 650898 356091 651134
rect 355771 650866 356091 650898
rect 370910 651454 371230 651486
rect 370910 651218 370952 651454
rect 371188 651218 371230 651454
rect 370910 651134 371230 651218
rect 370910 650898 370952 651134
rect 371188 650898 371230 651134
rect 370910 650866 371230 650898
rect 376840 651454 377160 651486
rect 376840 651218 376882 651454
rect 377118 651218 377160 651454
rect 376840 651134 377160 651218
rect 376840 650898 376882 651134
rect 377118 650898 377160 651134
rect 376840 650866 377160 650898
rect 382771 651454 383091 651486
rect 382771 651218 382813 651454
rect 383049 651218 383091 651454
rect 382771 651134 383091 651218
rect 382771 650898 382813 651134
rect 383049 650898 383091 651134
rect 382771 650866 383091 650898
rect 397910 651454 398230 651486
rect 397910 651218 397952 651454
rect 398188 651218 398230 651454
rect 397910 651134 398230 651218
rect 397910 650898 397952 651134
rect 398188 650898 398230 651134
rect 397910 650866 398230 650898
rect 403840 651454 404160 651486
rect 403840 651218 403882 651454
rect 404118 651218 404160 651454
rect 403840 651134 404160 651218
rect 403840 650898 403882 651134
rect 404118 650898 404160 651134
rect 403840 650866 404160 650898
rect 409771 651454 410091 651486
rect 409771 651218 409813 651454
rect 410049 651218 410091 651454
rect 409771 651134 410091 651218
rect 409771 650898 409813 651134
rect 410049 650898 410091 651134
rect 409771 650866 410091 650898
rect 424910 651454 425230 651486
rect 424910 651218 424952 651454
rect 425188 651218 425230 651454
rect 424910 651134 425230 651218
rect 424910 650898 424952 651134
rect 425188 650898 425230 651134
rect 424910 650866 425230 650898
rect 430840 651454 431160 651486
rect 430840 651218 430882 651454
rect 431118 651218 431160 651454
rect 430840 651134 431160 651218
rect 430840 650898 430882 651134
rect 431118 650898 431160 651134
rect 430840 650866 431160 650898
rect 436771 651454 437091 651486
rect 436771 651218 436813 651454
rect 437049 651218 437091 651454
rect 436771 651134 437091 651218
rect 436771 650898 436813 651134
rect 437049 650898 437091 651134
rect 436771 650866 437091 650898
rect 451910 651454 452230 651486
rect 451910 651218 451952 651454
rect 452188 651218 452230 651454
rect 451910 651134 452230 651218
rect 451910 650898 451952 651134
rect 452188 650898 452230 651134
rect 451910 650866 452230 650898
rect 457840 651454 458160 651486
rect 457840 651218 457882 651454
rect 458118 651218 458160 651454
rect 457840 651134 458160 651218
rect 457840 650898 457882 651134
rect 458118 650898 458160 651134
rect 457840 650866 458160 650898
rect 463771 651454 464091 651486
rect 463771 651218 463813 651454
rect 464049 651218 464091 651454
rect 463771 651134 464091 651218
rect 463771 650898 463813 651134
rect 464049 650898 464091 651134
rect 463771 650866 464091 650898
rect 478910 651454 479230 651486
rect 478910 651218 478952 651454
rect 479188 651218 479230 651454
rect 478910 651134 479230 651218
rect 478910 650898 478952 651134
rect 479188 650898 479230 651134
rect 478910 650866 479230 650898
rect 484840 651454 485160 651486
rect 484840 651218 484882 651454
rect 485118 651218 485160 651454
rect 484840 651134 485160 651218
rect 484840 650898 484882 651134
rect 485118 650898 485160 651134
rect 484840 650866 485160 650898
rect 490771 651454 491091 651486
rect 490771 651218 490813 651454
rect 491049 651218 491091 651454
rect 490771 651134 491091 651218
rect 490771 650898 490813 651134
rect 491049 650898 491091 651134
rect 490771 650866 491091 650898
rect 505910 651454 506230 651486
rect 505910 651218 505952 651454
rect 506188 651218 506230 651454
rect 505910 651134 506230 651218
rect 505910 650898 505952 651134
rect 506188 650898 506230 651134
rect 505910 650866 506230 650898
rect 511840 651454 512160 651486
rect 511840 651218 511882 651454
rect 512118 651218 512160 651454
rect 511840 651134 512160 651218
rect 511840 650898 511882 651134
rect 512118 650898 512160 651134
rect 511840 650866 512160 650898
rect 517771 651454 518091 651486
rect 517771 651218 517813 651454
rect 518049 651218 518091 651454
rect 517771 651134 518091 651218
rect 517771 650898 517813 651134
rect 518049 650898 518091 651134
rect 517771 650866 518091 650898
rect 532910 651454 533230 651486
rect 532910 651218 532952 651454
rect 533188 651218 533230 651454
rect 532910 651134 533230 651218
rect 532910 650898 532952 651134
rect 533188 650898 533230 651134
rect 532910 650866 533230 650898
rect 538840 651454 539160 651486
rect 538840 651218 538882 651454
rect 539118 651218 539160 651454
rect 538840 651134 539160 651218
rect 538840 650898 538882 651134
rect 539118 650898 539160 651134
rect 538840 650866 539160 650898
rect 544771 651454 545091 651486
rect 544771 651218 544813 651454
rect 545049 651218 545091 651454
rect 544771 651134 545091 651218
rect 544771 650898 544813 651134
rect 545049 650898 545091 651134
rect 544771 650866 545091 650898
rect 559794 651454 560414 668898
rect 559794 651218 559826 651454
rect 560062 651218 560146 651454
rect 560382 651218 560414 651454
rect 559794 651134 560414 651218
rect 559794 650898 559826 651134
rect 560062 650898 560146 651134
rect 560382 650898 560414 651134
rect 10794 642218 10826 642454
rect 11062 642218 11146 642454
rect 11382 642218 11414 642454
rect 10794 642134 11414 642218
rect 10794 641898 10826 642134
rect 11062 641898 11146 642134
rect 11382 641898 11414 642134
rect 10794 624454 11414 641898
rect 22874 642454 23194 642486
rect 22874 642218 22916 642454
rect 23152 642218 23194 642454
rect 22874 642134 23194 642218
rect 22874 641898 22916 642134
rect 23152 641898 23194 642134
rect 22874 641866 23194 641898
rect 28805 642454 29125 642486
rect 28805 642218 28847 642454
rect 29083 642218 29125 642454
rect 28805 642134 29125 642218
rect 28805 641898 28847 642134
rect 29083 641898 29125 642134
rect 28805 641866 29125 641898
rect 49874 642454 50194 642486
rect 49874 642218 49916 642454
rect 50152 642218 50194 642454
rect 49874 642134 50194 642218
rect 49874 641898 49916 642134
rect 50152 641898 50194 642134
rect 49874 641866 50194 641898
rect 55805 642454 56125 642486
rect 55805 642218 55847 642454
rect 56083 642218 56125 642454
rect 55805 642134 56125 642218
rect 55805 641898 55847 642134
rect 56083 641898 56125 642134
rect 55805 641866 56125 641898
rect 76874 642454 77194 642486
rect 76874 642218 76916 642454
rect 77152 642218 77194 642454
rect 76874 642134 77194 642218
rect 76874 641898 76916 642134
rect 77152 641898 77194 642134
rect 76874 641866 77194 641898
rect 82805 642454 83125 642486
rect 82805 642218 82847 642454
rect 83083 642218 83125 642454
rect 82805 642134 83125 642218
rect 82805 641898 82847 642134
rect 83083 641898 83125 642134
rect 82805 641866 83125 641898
rect 103874 642454 104194 642486
rect 103874 642218 103916 642454
rect 104152 642218 104194 642454
rect 103874 642134 104194 642218
rect 103874 641898 103916 642134
rect 104152 641898 104194 642134
rect 103874 641866 104194 641898
rect 109805 642454 110125 642486
rect 109805 642218 109847 642454
rect 110083 642218 110125 642454
rect 109805 642134 110125 642218
rect 109805 641898 109847 642134
rect 110083 641898 110125 642134
rect 109805 641866 110125 641898
rect 130874 642454 131194 642486
rect 130874 642218 130916 642454
rect 131152 642218 131194 642454
rect 130874 642134 131194 642218
rect 130874 641898 130916 642134
rect 131152 641898 131194 642134
rect 130874 641866 131194 641898
rect 136805 642454 137125 642486
rect 136805 642218 136847 642454
rect 137083 642218 137125 642454
rect 136805 642134 137125 642218
rect 136805 641898 136847 642134
rect 137083 641898 137125 642134
rect 136805 641866 137125 641898
rect 157874 642454 158194 642486
rect 157874 642218 157916 642454
rect 158152 642218 158194 642454
rect 157874 642134 158194 642218
rect 157874 641898 157916 642134
rect 158152 641898 158194 642134
rect 157874 641866 158194 641898
rect 163805 642454 164125 642486
rect 163805 642218 163847 642454
rect 164083 642218 164125 642454
rect 163805 642134 164125 642218
rect 163805 641898 163847 642134
rect 164083 641898 164125 642134
rect 163805 641866 164125 641898
rect 184874 642454 185194 642486
rect 184874 642218 184916 642454
rect 185152 642218 185194 642454
rect 184874 642134 185194 642218
rect 184874 641898 184916 642134
rect 185152 641898 185194 642134
rect 184874 641866 185194 641898
rect 190805 642454 191125 642486
rect 190805 642218 190847 642454
rect 191083 642218 191125 642454
rect 190805 642134 191125 642218
rect 190805 641898 190847 642134
rect 191083 641898 191125 642134
rect 190805 641866 191125 641898
rect 211874 642454 212194 642486
rect 211874 642218 211916 642454
rect 212152 642218 212194 642454
rect 211874 642134 212194 642218
rect 211874 641898 211916 642134
rect 212152 641898 212194 642134
rect 211874 641866 212194 641898
rect 217805 642454 218125 642486
rect 217805 642218 217847 642454
rect 218083 642218 218125 642454
rect 217805 642134 218125 642218
rect 217805 641898 217847 642134
rect 218083 641898 218125 642134
rect 217805 641866 218125 641898
rect 238874 642454 239194 642486
rect 238874 642218 238916 642454
rect 239152 642218 239194 642454
rect 238874 642134 239194 642218
rect 238874 641898 238916 642134
rect 239152 641898 239194 642134
rect 238874 641866 239194 641898
rect 244805 642454 245125 642486
rect 244805 642218 244847 642454
rect 245083 642218 245125 642454
rect 244805 642134 245125 642218
rect 244805 641898 244847 642134
rect 245083 641898 245125 642134
rect 244805 641866 245125 641898
rect 265874 642454 266194 642486
rect 265874 642218 265916 642454
rect 266152 642218 266194 642454
rect 265874 642134 266194 642218
rect 265874 641898 265916 642134
rect 266152 641898 266194 642134
rect 265874 641866 266194 641898
rect 271805 642454 272125 642486
rect 271805 642218 271847 642454
rect 272083 642218 272125 642454
rect 271805 642134 272125 642218
rect 271805 641898 271847 642134
rect 272083 641898 272125 642134
rect 271805 641866 272125 641898
rect 292874 642454 293194 642486
rect 292874 642218 292916 642454
rect 293152 642218 293194 642454
rect 292874 642134 293194 642218
rect 292874 641898 292916 642134
rect 293152 641898 293194 642134
rect 292874 641866 293194 641898
rect 298805 642454 299125 642486
rect 298805 642218 298847 642454
rect 299083 642218 299125 642454
rect 298805 642134 299125 642218
rect 298805 641898 298847 642134
rect 299083 641898 299125 642134
rect 298805 641866 299125 641898
rect 319874 642454 320194 642486
rect 319874 642218 319916 642454
rect 320152 642218 320194 642454
rect 319874 642134 320194 642218
rect 319874 641898 319916 642134
rect 320152 641898 320194 642134
rect 319874 641866 320194 641898
rect 325805 642454 326125 642486
rect 325805 642218 325847 642454
rect 326083 642218 326125 642454
rect 325805 642134 326125 642218
rect 325805 641898 325847 642134
rect 326083 641898 326125 642134
rect 325805 641866 326125 641898
rect 346874 642454 347194 642486
rect 346874 642218 346916 642454
rect 347152 642218 347194 642454
rect 346874 642134 347194 642218
rect 346874 641898 346916 642134
rect 347152 641898 347194 642134
rect 346874 641866 347194 641898
rect 352805 642454 353125 642486
rect 352805 642218 352847 642454
rect 353083 642218 353125 642454
rect 352805 642134 353125 642218
rect 352805 641898 352847 642134
rect 353083 641898 353125 642134
rect 352805 641866 353125 641898
rect 373874 642454 374194 642486
rect 373874 642218 373916 642454
rect 374152 642218 374194 642454
rect 373874 642134 374194 642218
rect 373874 641898 373916 642134
rect 374152 641898 374194 642134
rect 373874 641866 374194 641898
rect 379805 642454 380125 642486
rect 379805 642218 379847 642454
rect 380083 642218 380125 642454
rect 379805 642134 380125 642218
rect 379805 641898 379847 642134
rect 380083 641898 380125 642134
rect 379805 641866 380125 641898
rect 400874 642454 401194 642486
rect 400874 642218 400916 642454
rect 401152 642218 401194 642454
rect 400874 642134 401194 642218
rect 400874 641898 400916 642134
rect 401152 641898 401194 642134
rect 400874 641866 401194 641898
rect 406805 642454 407125 642486
rect 406805 642218 406847 642454
rect 407083 642218 407125 642454
rect 406805 642134 407125 642218
rect 406805 641898 406847 642134
rect 407083 641898 407125 642134
rect 406805 641866 407125 641898
rect 427874 642454 428194 642486
rect 427874 642218 427916 642454
rect 428152 642218 428194 642454
rect 427874 642134 428194 642218
rect 427874 641898 427916 642134
rect 428152 641898 428194 642134
rect 427874 641866 428194 641898
rect 433805 642454 434125 642486
rect 433805 642218 433847 642454
rect 434083 642218 434125 642454
rect 433805 642134 434125 642218
rect 433805 641898 433847 642134
rect 434083 641898 434125 642134
rect 433805 641866 434125 641898
rect 454874 642454 455194 642486
rect 454874 642218 454916 642454
rect 455152 642218 455194 642454
rect 454874 642134 455194 642218
rect 454874 641898 454916 642134
rect 455152 641898 455194 642134
rect 454874 641866 455194 641898
rect 460805 642454 461125 642486
rect 460805 642218 460847 642454
rect 461083 642218 461125 642454
rect 460805 642134 461125 642218
rect 460805 641898 460847 642134
rect 461083 641898 461125 642134
rect 460805 641866 461125 641898
rect 481874 642454 482194 642486
rect 481874 642218 481916 642454
rect 482152 642218 482194 642454
rect 481874 642134 482194 642218
rect 481874 641898 481916 642134
rect 482152 641898 482194 642134
rect 481874 641866 482194 641898
rect 487805 642454 488125 642486
rect 487805 642218 487847 642454
rect 488083 642218 488125 642454
rect 487805 642134 488125 642218
rect 487805 641898 487847 642134
rect 488083 641898 488125 642134
rect 487805 641866 488125 641898
rect 508874 642454 509194 642486
rect 508874 642218 508916 642454
rect 509152 642218 509194 642454
rect 508874 642134 509194 642218
rect 508874 641898 508916 642134
rect 509152 641898 509194 642134
rect 508874 641866 509194 641898
rect 514805 642454 515125 642486
rect 514805 642218 514847 642454
rect 515083 642218 515125 642454
rect 514805 642134 515125 642218
rect 514805 641898 514847 642134
rect 515083 641898 515125 642134
rect 514805 641866 515125 641898
rect 535874 642454 536194 642486
rect 535874 642218 535916 642454
rect 536152 642218 536194 642454
rect 535874 642134 536194 642218
rect 535874 641898 535916 642134
rect 536152 641898 536194 642134
rect 535874 641866 536194 641898
rect 541805 642454 542125 642486
rect 541805 642218 541847 642454
rect 542083 642218 542125 642454
rect 541805 642134 542125 642218
rect 541805 641898 541847 642134
rect 542083 641898 542125 642134
rect 541805 641866 542125 641898
rect 19794 633454 20414 635000
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 632000 20414 632898
rect 28794 634394 29414 635000
rect 28794 634158 28826 634394
rect 29062 634158 29146 634394
rect 29382 634158 29414 634394
rect 28794 634074 29414 634158
rect 28794 633838 28826 634074
rect 29062 633838 29146 634074
rect 29382 633838 29414 634074
rect 28794 632000 29414 633838
rect 37794 633454 38414 635000
rect 37794 633218 37826 633454
rect 38062 633218 38146 633454
rect 38382 633218 38414 633454
rect 37794 633134 38414 633218
rect 37794 632898 37826 633134
rect 38062 632898 38146 633134
rect 38382 632898 38414 633134
rect 37794 632000 38414 632898
rect 46794 634394 47414 635000
rect 46794 634158 46826 634394
rect 47062 634158 47146 634394
rect 47382 634158 47414 634394
rect 46794 634074 47414 634158
rect 46794 633838 46826 634074
rect 47062 633838 47146 634074
rect 47382 633838 47414 634074
rect 46794 632000 47414 633838
rect 55794 633454 56414 635000
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 632000 56414 632898
rect 64794 634394 65414 635000
rect 64794 634158 64826 634394
rect 65062 634158 65146 634394
rect 65382 634158 65414 634394
rect 64794 634074 65414 634158
rect 64794 633838 64826 634074
rect 65062 633838 65146 634074
rect 65382 633838 65414 634074
rect 64794 632000 65414 633838
rect 73794 633454 74414 635000
rect 73794 633218 73826 633454
rect 74062 633218 74146 633454
rect 74382 633218 74414 633454
rect 73794 633134 74414 633218
rect 73794 632898 73826 633134
rect 74062 632898 74146 633134
rect 74382 632898 74414 633134
rect 73794 632000 74414 632898
rect 82794 634394 83414 635000
rect 82794 634158 82826 634394
rect 83062 634158 83146 634394
rect 83382 634158 83414 634394
rect 82794 634074 83414 634158
rect 82794 633838 82826 634074
rect 83062 633838 83146 634074
rect 83382 633838 83414 634074
rect 82794 632000 83414 633838
rect 91794 633454 92414 635000
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 632000 92414 632898
rect 100794 634394 101414 635000
rect 100794 634158 100826 634394
rect 101062 634158 101146 634394
rect 101382 634158 101414 634394
rect 100794 634074 101414 634158
rect 100794 633838 100826 634074
rect 101062 633838 101146 634074
rect 101382 633838 101414 634074
rect 100794 632000 101414 633838
rect 109794 633454 110414 635000
rect 109794 633218 109826 633454
rect 110062 633218 110146 633454
rect 110382 633218 110414 633454
rect 109794 633134 110414 633218
rect 109794 632898 109826 633134
rect 110062 632898 110146 633134
rect 110382 632898 110414 633134
rect 109794 632000 110414 632898
rect 118794 634394 119414 635000
rect 118794 634158 118826 634394
rect 119062 634158 119146 634394
rect 119382 634158 119414 634394
rect 118794 634074 119414 634158
rect 118794 633838 118826 634074
rect 119062 633838 119146 634074
rect 119382 633838 119414 634074
rect 118794 632000 119414 633838
rect 127794 633454 128414 635000
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 632000 128414 632898
rect 136794 634394 137414 635000
rect 136794 634158 136826 634394
rect 137062 634158 137146 634394
rect 137382 634158 137414 634394
rect 136794 634074 137414 634158
rect 136794 633838 136826 634074
rect 137062 633838 137146 634074
rect 137382 633838 137414 634074
rect 136794 632000 137414 633838
rect 145794 633454 146414 635000
rect 145794 633218 145826 633454
rect 146062 633218 146146 633454
rect 146382 633218 146414 633454
rect 145794 633134 146414 633218
rect 145794 632898 145826 633134
rect 146062 632898 146146 633134
rect 146382 632898 146414 633134
rect 145794 632000 146414 632898
rect 154794 634394 155414 635000
rect 154794 634158 154826 634394
rect 155062 634158 155146 634394
rect 155382 634158 155414 634394
rect 154794 634074 155414 634158
rect 154794 633838 154826 634074
rect 155062 633838 155146 634074
rect 155382 633838 155414 634074
rect 154794 632000 155414 633838
rect 163794 633454 164414 635000
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 632000 164414 632898
rect 172794 634394 173414 635000
rect 172794 634158 172826 634394
rect 173062 634158 173146 634394
rect 173382 634158 173414 634394
rect 172794 634074 173414 634158
rect 172794 633838 172826 634074
rect 173062 633838 173146 634074
rect 173382 633838 173414 634074
rect 172794 632000 173414 633838
rect 181794 633454 182414 635000
rect 181794 633218 181826 633454
rect 182062 633218 182146 633454
rect 182382 633218 182414 633454
rect 181794 633134 182414 633218
rect 181794 632898 181826 633134
rect 182062 632898 182146 633134
rect 182382 632898 182414 633134
rect 181794 632000 182414 632898
rect 190794 634394 191414 635000
rect 190794 634158 190826 634394
rect 191062 634158 191146 634394
rect 191382 634158 191414 634394
rect 190794 634074 191414 634158
rect 190794 633838 190826 634074
rect 191062 633838 191146 634074
rect 191382 633838 191414 634074
rect 190794 632000 191414 633838
rect 199794 633454 200414 635000
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 632000 200414 632898
rect 208794 634394 209414 635000
rect 208794 634158 208826 634394
rect 209062 634158 209146 634394
rect 209382 634158 209414 634394
rect 208794 634074 209414 634158
rect 208794 633838 208826 634074
rect 209062 633838 209146 634074
rect 209382 633838 209414 634074
rect 208794 632000 209414 633838
rect 217794 633454 218414 635000
rect 217794 633218 217826 633454
rect 218062 633218 218146 633454
rect 218382 633218 218414 633454
rect 217794 633134 218414 633218
rect 217794 632898 217826 633134
rect 218062 632898 218146 633134
rect 218382 632898 218414 633134
rect 217794 632000 218414 632898
rect 226794 634394 227414 635000
rect 226794 634158 226826 634394
rect 227062 634158 227146 634394
rect 227382 634158 227414 634394
rect 226794 634074 227414 634158
rect 226794 633838 226826 634074
rect 227062 633838 227146 634074
rect 227382 633838 227414 634074
rect 226794 632000 227414 633838
rect 235794 633454 236414 635000
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 632000 236414 632898
rect 244794 634394 245414 635000
rect 244794 634158 244826 634394
rect 245062 634158 245146 634394
rect 245382 634158 245414 634394
rect 244794 634074 245414 634158
rect 244794 633838 244826 634074
rect 245062 633838 245146 634074
rect 245382 633838 245414 634074
rect 244794 632000 245414 633838
rect 253794 633454 254414 635000
rect 253794 633218 253826 633454
rect 254062 633218 254146 633454
rect 254382 633218 254414 633454
rect 253794 633134 254414 633218
rect 253794 632898 253826 633134
rect 254062 632898 254146 633134
rect 254382 632898 254414 633134
rect 253794 632000 254414 632898
rect 262794 634394 263414 635000
rect 262794 634158 262826 634394
rect 263062 634158 263146 634394
rect 263382 634158 263414 634394
rect 262794 634074 263414 634158
rect 262794 633838 262826 634074
rect 263062 633838 263146 634074
rect 263382 633838 263414 634074
rect 262794 632000 263414 633838
rect 271794 633454 272414 635000
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 632000 272414 632898
rect 280794 634394 281414 635000
rect 280794 634158 280826 634394
rect 281062 634158 281146 634394
rect 281382 634158 281414 634394
rect 280794 634074 281414 634158
rect 280794 633838 280826 634074
rect 281062 633838 281146 634074
rect 281382 633838 281414 634074
rect 280794 632000 281414 633838
rect 289794 633454 290414 635000
rect 289794 633218 289826 633454
rect 290062 633218 290146 633454
rect 290382 633218 290414 633454
rect 289794 633134 290414 633218
rect 289794 632898 289826 633134
rect 290062 632898 290146 633134
rect 290382 632898 290414 633134
rect 289794 632000 290414 632898
rect 298794 634394 299414 635000
rect 298794 634158 298826 634394
rect 299062 634158 299146 634394
rect 299382 634158 299414 634394
rect 298794 634074 299414 634158
rect 298794 633838 298826 634074
rect 299062 633838 299146 634074
rect 299382 633838 299414 634074
rect 298794 632000 299414 633838
rect 307794 633454 308414 635000
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 632000 308414 632898
rect 316794 634394 317414 635000
rect 316794 634158 316826 634394
rect 317062 634158 317146 634394
rect 317382 634158 317414 634394
rect 316794 634074 317414 634158
rect 316794 633838 316826 634074
rect 317062 633838 317146 634074
rect 317382 633838 317414 634074
rect 316794 632000 317414 633838
rect 325794 633454 326414 635000
rect 325794 633218 325826 633454
rect 326062 633218 326146 633454
rect 326382 633218 326414 633454
rect 325794 633134 326414 633218
rect 325794 632898 325826 633134
rect 326062 632898 326146 633134
rect 326382 632898 326414 633134
rect 325794 632000 326414 632898
rect 334794 634394 335414 635000
rect 334794 634158 334826 634394
rect 335062 634158 335146 634394
rect 335382 634158 335414 634394
rect 334794 634074 335414 634158
rect 334794 633838 334826 634074
rect 335062 633838 335146 634074
rect 335382 633838 335414 634074
rect 334794 632000 335414 633838
rect 343794 633454 344414 635000
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 632000 344414 632898
rect 352794 634394 353414 635000
rect 352794 634158 352826 634394
rect 353062 634158 353146 634394
rect 353382 634158 353414 634394
rect 352794 634074 353414 634158
rect 352794 633838 352826 634074
rect 353062 633838 353146 634074
rect 353382 633838 353414 634074
rect 352794 632000 353414 633838
rect 361794 633454 362414 635000
rect 361794 633218 361826 633454
rect 362062 633218 362146 633454
rect 362382 633218 362414 633454
rect 361794 633134 362414 633218
rect 361794 632898 361826 633134
rect 362062 632898 362146 633134
rect 362382 632898 362414 633134
rect 361794 632000 362414 632898
rect 370794 634394 371414 635000
rect 370794 634158 370826 634394
rect 371062 634158 371146 634394
rect 371382 634158 371414 634394
rect 370794 634074 371414 634158
rect 370794 633838 370826 634074
rect 371062 633838 371146 634074
rect 371382 633838 371414 634074
rect 370794 632000 371414 633838
rect 379794 633454 380414 635000
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 632000 380414 632898
rect 388794 634394 389414 635000
rect 388794 634158 388826 634394
rect 389062 634158 389146 634394
rect 389382 634158 389414 634394
rect 388794 634074 389414 634158
rect 388794 633838 388826 634074
rect 389062 633838 389146 634074
rect 389382 633838 389414 634074
rect 388794 632000 389414 633838
rect 397794 633454 398414 635000
rect 397794 633218 397826 633454
rect 398062 633218 398146 633454
rect 398382 633218 398414 633454
rect 397794 633134 398414 633218
rect 397794 632898 397826 633134
rect 398062 632898 398146 633134
rect 398382 632898 398414 633134
rect 397794 632000 398414 632898
rect 406794 634394 407414 635000
rect 406794 634158 406826 634394
rect 407062 634158 407146 634394
rect 407382 634158 407414 634394
rect 406794 634074 407414 634158
rect 406794 633838 406826 634074
rect 407062 633838 407146 634074
rect 407382 633838 407414 634074
rect 406794 632000 407414 633838
rect 415794 633454 416414 635000
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 632000 416414 632898
rect 424794 634394 425414 635000
rect 424794 634158 424826 634394
rect 425062 634158 425146 634394
rect 425382 634158 425414 634394
rect 424794 634074 425414 634158
rect 424794 633838 424826 634074
rect 425062 633838 425146 634074
rect 425382 633838 425414 634074
rect 424794 632000 425414 633838
rect 433794 633454 434414 635000
rect 433794 633218 433826 633454
rect 434062 633218 434146 633454
rect 434382 633218 434414 633454
rect 433794 633134 434414 633218
rect 433794 632898 433826 633134
rect 434062 632898 434146 633134
rect 434382 632898 434414 633134
rect 433794 632000 434414 632898
rect 442794 634394 443414 635000
rect 442794 634158 442826 634394
rect 443062 634158 443146 634394
rect 443382 634158 443414 634394
rect 442794 634074 443414 634158
rect 442794 633838 442826 634074
rect 443062 633838 443146 634074
rect 443382 633838 443414 634074
rect 442794 632000 443414 633838
rect 451794 633454 452414 635000
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 632000 452414 632898
rect 460794 634394 461414 635000
rect 460794 634158 460826 634394
rect 461062 634158 461146 634394
rect 461382 634158 461414 634394
rect 460794 634074 461414 634158
rect 460794 633838 460826 634074
rect 461062 633838 461146 634074
rect 461382 633838 461414 634074
rect 460794 632000 461414 633838
rect 469794 633454 470414 635000
rect 469794 633218 469826 633454
rect 470062 633218 470146 633454
rect 470382 633218 470414 633454
rect 469794 633134 470414 633218
rect 469794 632898 469826 633134
rect 470062 632898 470146 633134
rect 470382 632898 470414 633134
rect 469794 632000 470414 632898
rect 478794 634394 479414 635000
rect 478794 634158 478826 634394
rect 479062 634158 479146 634394
rect 479382 634158 479414 634394
rect 478794 634074 479414 634158
rect 478794 633838 478826 634074
rect 479062 633838 479146 634074
rect 479382 633838 479414 634074
rect 478794 632000 479414 633838
rect 487794 633454 488414 635000
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 632000 488414 632898
rect 496794 634394 497414 635000
rect 496794 634158 496826 634394
rect 497062 634158 497146 634394
rect 497382 634158 497414 634394
rect 496794 634074 497414 634158
rect 496794 633838 496826 634074
rect 497062 633838 497146 634074
rect 497382 633838 497414 634074
rect 496794 632000 497414 633838
rect 505794 633454 506414 635000
rect 505794 633218 505826 633454
rect 506062 633218 506146 633454
rect 506382 633218 506414 633454
rect 505794 633134 506414 633218
rect 505794 632898 505826 633134
rect 506062 632898 506146 633134
rect 506382 632898 506414 633134
rect 505794 632000 506414 632898
rect 514794 634394 515414 635000
rect 514794 634158 514826 634394
rect 515062 634158 515146 634394
rect 515382 634158 515414 634394
rect 514794 634074 515414 634158
rect 514794 633838 514826 634074
rect 515062 633838 515146 634074
rect 515382 633838 515414 634074
rect 514794 632000 515414 633838
rect 523794 633454 524414 635000
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 632000 524414 632898
rect 532794 634394 533414 635000
rect 532794 634158 532826 634394
rect 533062 634158 533146 634394
rect 533382 634158 533414 634394
rect 532794 634074 533414 634158
rect 532794 633838 532826 634074
rect 533062 633838 533146 634074
rect 533382 633838 533414 634074
rect 532794 632000 533414 633838
rect 541794 633454 542414 635000
rect 541794 633218 541826 633454
rect 542062 633218 542146 633454
rect 542382 633218 542414 633454
rect 541794 633134 542414 633218
rect 541794 632898 541826 633134
rect 542062 632898 542146 633134
rect 542382 632898 542414 633134
rect 541794 632000 542414 632898
rect 550794 634394 551414 635000
rect 550794 634158 550826 634394
rect 551062 634158 551146 634394
rect 551382 634158 551414 634394
rect 550794 634074 551414 634158
rect 550794 633838 550826 634074
rect 551062 633838 551146 634074
rect 551382 633838 551414 634074
rect 550794 632000 551414 633838
rect 559794 633454 560414 650898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 606454 11414 623898
rect 22874 624454 23194 624486
rect 22874 624218 22916 624454
rect 23152 624218 23194 624454
rect 22874 624134 23194 624218
rect 22874 623898 22916 624134
rect 23152 623898 23194 624134
rect 22874 623866 23194 623898
rect 28805 624454 29125 624486
rect 28805 624218 28847 624454
rect 29083 624218 29125 624454
rect 28805 624134 29125 624218
rect 28805 623898 28847 624134
rect 29083 623898 29125 624134
rect 28805 623866 29125 623898
rect 49874 624454 50194 624486
rect 49874 624218 49916 624454
rect 50152 624218 50194 624454
rect 49874 624134 50194 624218
rect 49874 623898 49916 624134
rect 50152 623898 50194 624134
rect 49874 623866 50194 623898
rect 55805 624454 56125 624486
rect 55805 624218 55847 624454
rect 56083 624218 56125 624454
rect 55805 624134 56125 624218
rect 55805 623898 55847 624134
rect 56083 623898 56125 624134
rect 55805 623866 56125 623898
rect 76874 624454 77194 624486
rect 76874 624218 76916 624454
rect 77152 624218 77194 624454
rect 76874 624134 77194 624218
rect 76874 623898 76916 624134
rect 77152 623898 77194 624134
rect 76874 623866 77194 623898
rect 82805 624454 83125 624486
rect 82805 624218 82847 624454
rect 83083 624218 83125 624454
rect 82805 624134 83125 624218
rect 82805 623898 82847 624134
rect 83083 623898 83125 624134
rect 82805 623866 83125 623898
rect 103874 624454 104194 624486
rect 103874 624218 103916 624454
rect 104152 624218 104194 624454
rect 103874 624134 104194 624218
rect 103874 623898 103916 624134
rect 104152 623898 104194 624134
rect 103874 623866 104194 623898
rect 109805 624454 110125 624486
rect 109805 624218 109847 624454
rect 110083 624218 110125 624454
rect 109805 624134 110125 624218
rect 109805 623898 109847 624134
rect 110083 623898 110125 624134
rect 109805 623866 110125 623898
rect 130874 624454 131194 624486
rect 130874 624218 130916 624454
rect 131152 624218 131194 624454
rect 130874 624134 131194 624218
rect 130874 623898 130916 624134
rect 131152 623898 131194 624134
rect 130874 623866 131194 623898
rect 136805 624454 137125 624486
rect 136805 624218 136847 624454
rect 137083 624218 137125 624454
rect 136805 624134 137125 624218
rect 136805 623898 136847 624134
rect 137083 623898 137125 624134
rect 136805 623866 137125 623898
rect 157874 624454 158194 624486
rect 157874 624218 157916 624454
rect 158152 624218 158194 624454
rect 157874 624134 158194 624218
rect 157874 623898 157916 624134
rect 158152 623898 158194 624134
rect 157874 623866 158194 623898
rect 163805 624454 164125 624486
rect 163805 624218 163847 624454
rect 164083 624218 164125 624454
rect 163805 624134 164125 624218
rect 163805 623898 163847 624134
rect 164083 623898 164125 624134
rect 163805 623866 164125 623898
rect 184874 624454 185194 624486
rect 184874 624218 184916 624454
rect 185152 624218 185194 624454
rect 184874 624134 185194 624218
rect 184874 623898 184916 624134
rect 185152 623898 185194 624134
rect 184874 623866 185194 623898
rect 190805 624454 191125 624486
rect 190805 624218 190847 624454
rect 191083 624218 191125 624454
rect 190805 624134 191125 624218
rect 190805 623898 190847 624134
rect 191083 623898 191125 624134
rect 190805 623866 191125 623898
rect 211874 624454 212194 624486
rect 211874 624218 211916 624454
rect 212152 624218 212194 624454
rect 211874 624134 212194 624218
rect 211874 623898 211916 624134
rect 212152 623898 212194 624134
rect 211874 623866 212194 623898
rect 217805 624454 218125 624486
rect 217805 624218 217847 624454
rect 218083 624218 218125 624454
rect 217805 624134 218125 624218
rect 217805 623898 217847 624134
rect 218083 623898 218125 624134
rect 217805 623866 218125 623898
rect 238874 624454 239194 624486
rect 238874 624218 238916 624454
rect 239152 624218 239194 624454
rect 238874 624134 239194 624218
rect 238874 623898 238916 624134
rect 239152 623898 239194 624134
rect 238874 623866 239194 623898
rect 244805 624454 245125 624486
rect 244805 624218 244847 624454
rect 245083 624218 245125 624454
rect 244805 624134 245125 624218
rect 244805 623898 244847 624134
rect 245083 623898 245125 624134
rect 244805 623866 245125 623898
rect 265874 624454 266194 624486
rect 265874 624218 265916 624454
rect 266152 624218 266194 624454
rect 265874 624134 266194 624218
rect 265874 623898 265916 624134
rect 266152 623898 266194 624134
rect 265874 623866 266194 623898
rect 271805 624454 272125 624486
rect 271805 624218 271847 624454
rect 272083 624218 272125 624454
rect 271805 624134 272125 624218
rect 271805 623898 271847 624134
rect 272083 623898 272125 624134
rect 271805 623866 272125 623898
rect 292874 624454 293194 624486
rect 292874 624218 292916 624454
rect 293152 624218 293194 624454
rect 292874 624134 293194 624218
rect 292874 623898 292916 624134
rect 293152 623898 293194 624134
rect 292874 623866 293194 623898
rect 298805 624454 299125 624486
rect 298805 624218 298847 624454
rect 299083 624218 299125 624454
rect 298805 624134 299125 624218
rect 298805 623898 298847 624134
rect 299083 623898 299125 624134
rect 298805 623866 299125 623898
rect 319874 624454 320194 624486
rect 319874 624218 319916 624454
rect 320152 624218 320194 624454
rect 319874 624134 320194 624218
rect 319874 623898 319916 624134
rect 320152 623898 320194 624134
rect 319874 623866 320194 623898
rect 325805 624454 326125 624486
rect 325805 624218 325847 624454
rect 326083 624218 326125 624454
rect 325805 624134 326125 624218
rect 325805 623898 325847 624134
rect 326083 623898 326125 624134
rect 325805 623866 326125 623898
rect 346874 624454 347194 624486
rect 346874 624218 346916 624454
rect 347152 624218 347194 624454
rect 346874 624134 347194 624218
rect 346874 623898 346916 624134
rect 347152 623898 347194 624134
rect 346874 623866 347194 623898
rect 352805 624454 353125 624486
rect 352805 624218 352847 624454
rect 353083 624218 353125 624454
rect 352805 624134 353125 624218
rect 352805 623898 352847 624134
rect 353083 623898 353125 624134
rect 352805 623866 353125 623898
rect 373874 624454 374194 624486
rect 373874 624218 373916 624454
rect 374152 624218 374194 624454
rect 373874 624134 374194 624218
rect 373874 623898 373916 624134
rect 374152 623898 374194 624134
rect 373874 623866 374194 623898
rect 379805 624454 380125 624486
rect 379805 624218 379847 624454
rect 380083 624218 380125 624454
rect 379805 624134 380125 624218
rect 379805 623898 379847 624134
rect 380083 623898 380125 624134
rect 379805 623866 380125 623898
rect 400874 624454 401194 624486
rect 400874 624218 400916 624454
rect 401152 624218 401194 624454
rect 400874 624134 401194 624218
rect 400874 623898 400916 624134
rect 401152 623898 401194 624134
rect 400874 623866 401194 623898
rect 406805 624454 407125 624486
rect 406805 624218 406847 624454
rect 407083 624218 407125 624454
rect 406805 624134 407125 624218
rect 406805 623898 406847 624134
rect 407083 623898 407125 624134
rect 406805 623866 407125 623898
rect 427874 624454 428194 624486
rect 427874 624218 427916 624454
rect 428152 624218 428194 624454
rect 427874 624134 428194 624218
rect 427874 623898 427916 624134
rect 428152 623898 428194 624134
rect 427874 623866 428194 623898
rect 433805 624454 434125 624486
rect 433805 624218 433847 624454
rect 434083 624218 434125 624454
rect 433805 624134 434125 624218
rect 433805 623898 433847 624134
rect 434083 623898 434125 624134
rect 433805 623866 434125 623898
rect 454874 624454 455194 624486
rect 454874 624218 454916 624454
rect 455152 624218 455194 624454
rect 454874 624134 455194 624218
rect 454874 623898 454916 624134
rect 455152 623898 455194 624134
rect 454874 623866 455194 623898
rect 460805 624454 461125 624486
rect 460805 624218 460847 624454
rect 461083 624218 461125 624454
rect 460805 624134 461125 624218
rect 460805 623898 460847 624134
rect 461083 623898 461125 624134
rect 460805 623866 461125 623898
rect 481874 624454 482194 624486
rect 481874 624218 481916 624454
rect 482152 624218 482194 624454
rect 481874 624134 482194 624218
rect 481874 623898 481916 624134
rect 482152 623898 482194 624134
rect 481874 623866 482194 623898
rect 487805 624454 488125 624486
rect 487805 624218 487847 624454
rect 488083 624218 488125 624454
rect 487805 624134 488125 624218
rect 487805 623898 487847 624134
rect 488083 623898 488125 624134
rect 487805 623866 488125 623898
rect 508874 624454 509194 624486
rect 508874 624218 508916 624454
rect 509152 624218 509194 624454
rect 508874 624134 509194 624218
rect 508874 623898 508916 624134
rect 509152 623898 509194 624134
rect 508874 623866 509194 623898
rect 514805 624454 515125 624486
rect 514805 624218 514847 624454
rect 515083 624218 515125 624454
rect 514805 624134 515125 624218
rect 514805 623898 514847 624134
rect 515083 623898 515125 624134
rect 514805 623866 515125 623898
rect 535874 624454 536194 624486
rect 535874 624218 535916 624454
rect 536152 624218 536194 624454
rect 535874 624134 536194 624218
rect 535874 623898 535916 624134
rect 536152 623898 536194 624134
rect 535874 623866 536194 623898
rect 541805 624454 542125 624486
rect 541805 624218 541847 624454
rect 542083 624218 542125 624454
rect 541805 624134 542125 624218
rect 541805 623898 541847 624134
rect 542083 623898 542125 624134
rect 541805 623866 542125 623898
rect 19910 615454 20230 615486
rect 19910 615218 19952 615454
rect 20188 615218 20230 615454
rect 19910 615134 20230 615218
rect 19910 614898 19952 615134
rect 20188 614898 20230 615134
rect 19910 614866 20230 614898
rect 25840 615454 26160 615486
rect 25840 615218 25882 615454
rect 26118 615218 26160 615454
rect 25840 615134 26160 615218
rect 25840 614898 25882 615134
rect 26118 614898 26160 615134
rect 25840 614866 26160 614898
rect 31771 615454 32091 615486
rect 31771 615218 31813 615454
rect 32049 615218 32091 615454
rect 31771 615134 32091 615218
rect 31771 614898 31813 615134
rect 32049 614898 32091 615134
rect 31771 614866 32091 614898
rect 46910 615454 47230 615486
rect 46910 615218 46952 615454
rect 47188 615218 47230 615454
rect 46910 615134 47230 615218
rect 46910 614898 46952 615134
rect 47188 614898 47230 615134
rect 46910 614866 47230 614898
rect 52840 615454 53160 615486
rect 52840 615218 52882 615454
rect 53118 615218 53160 615454
rect 52840 615134 53160 615218
rect 52840 614898 52882 615134
rect 53118 614898 53160 615134
rect 52840 614866 53160 614898
rect 58771 615454 59091 615486
rect 58771 615218 58813 615454
rect 59049 615218 59091 615454
rect 58771 615134 59091 615218
rect 58771 614898 58813 615134
rect 59049 614898 59091 615134
rect 58771 614866 59091 614898
rect 73910 615454 74230 615486
rect 73910 615218 73952 615454
rect 74188 615218 74230 615454
rect 73910 615134 74230 615218
rect 73910 614898 73952 615134
rect 74188 614898 74230 615134
rect 73910 614866 74230 614898
rect 79840 615454 80160 615486
rect 79840 615218 79882 615454
rect 80118 615218 80160 615454
rect 79840 615134 80160 615218
rect 79840 614898 79882 615134
rect 80118 614898 80160 615134
rect 79840 614866 80160 614898
rect 85771 615454 86091 615486
rect 85771 615218 85813 615454
rect 86049 615218 86091 615454
rect 85771 615134 86091 615218
rect 85771 614898 85813 615134
rect 86049 614898 86091 615134
rect 85771 614866 86091 614898
rect 100910 615454 101230 615486
rect 100910 615218 100952 615454
rect 101188 615218 101230 615454
rect 100910 615134 101230 615218
rect 100910 614898 100952 615134
rect 101188 614898 101230 615134
rect 100910 614866 101230 614898
rect 106840 615454 107160 615486
rect 106840 615218 106882 615454
rect 107118 615218 107160 615454
rect 106840 615134 107160 615218
rect 106840 614898 106882 615134
rect 107118 614898 107160 615134
rect 106840 614866 107160 614898
rect 112771 615454 113091 615486
rect 112771 615218 112813 615454
rect 113049 615218 113091 615454
rect 112771 615134 113091 615218
rect 112771 614898 112813 615134
rect 113049 614898 113091 615134
rect 112771 614866 113091 614898
rect 127910 615454 128230 615486
rect 127910 615218 127952 615454
rect 128188 615218 128230 615454
rect 127910 615134 128230 615218
rect 127910 614898 127952 615134
rect 128188 614898 128230 615134
rect 127910 614866 128230 614898
rect 133840 615454 134160 615486
rect 133840 615218 133882 615454
rect 134118 615218 134160 615454
rect 133840 615134 134160 615218
rect 133840 614898 133882 615134
rect 134118 614898 134160 615134
rect 133840 614866 134160 614898
rect 139771 615454 140091 615486
rect 139771 615218 139813 615454
rect 140049 615218 140091 615454
rect 139771 615134 140091 615218
rect 139771 614898 139813 615134
rect 140049 614898 140091 615134
rect 139771 614866 140091 614898
rect 154910 615454 155230 615486
rect 154910 615218 154952 615454
rect 155188 615218 155230 615454
rect 154910 615134 155230 615218
rect 154910 614898 154952 615134
rect 155188 614898 155230 615134
rect 154910 614866 155230 614898
rect 160840 615454 161160 615486
rect 160840 615218 160882 615454
rect 161118 615218 161160 615454
rect 160840 615134 161160 615218
rect 160840 614898 160882 615134
rect 161118 614898 161160 615134
rect 160840 614866 161160 614898
rect 166771 615454 167091 615486
rect 166771 615218 166813 615454
rect 167049 615218 167091 615454
rect 166771 615134 167091 615218
rect 166771 614898 166813 615134
rect 167049 614898 167091 615134
rect 166771 614866 167091 614898
rect 181910 615454 182230 615486
rect 181910 615218 181952 615454
rect 182188 615218 182230 615454
rect 181910 615134 182230 615218
rect 181910 614898 181952 615134
rect 182188 614898 182230 615134
rect 181910 614866 182230 614898
rect 187840 615454 188160 615486
rect 187840 615218 187882 615454
rect 188118 615218 188160 615454
rect 187840 615134 188160 615218
rect 187840 614898 187882 615134
rect 188118 614898 188160 615134
rect 187840 614866 188160 614898
rect 193771 615454 194091 615486
rect 193771 615218 193813 615454
rect 194049 615218 194091 615454
rect 193771 615134 194091 615218
rect 193771 614898 193813 615134
rect 194049 614898 194091 615134
rect 193771 614866 194091 614898
rect 208910 615454 209230 615486
rect 208910 615218 208952 615454
rect 209188 615218 209230 615454
rect 208910 615134 209230 615218
rect 208910 614898 208952 615134
rect 209188 614898 209230 615134
rect 208910 614866 209230 614898
rect 214840 615454 215160 615486
rect 214840 615218 214882 615454
rect 215118 615218 215160 615454
rect 214840 615134 215160 615218
rect 214840 614898 214882 615134
rect 215118 614898 215160 615134
rect 214840 614866 215160 614898
rect 220771 615454 221091 615486
rect 220771 615218 220813 615454
rect 221049 615218 221091 615454
rect 220771 615134 221091 615218
rect 220771 614898 220813 615134
rect 221049 614898 221091 615134
rect 220771 614866 221091 614898
rect 235910 615454 236230 615486
rect 235910 615218 235952 615454
rect 236188 615218 236230 615454
rect 235910 615134 236230 615218
rect 235910 614898 235952 615134
rect 236188 614898 236230 615134
rect 235910 614866 236230 614898
rect 241840 615454 242160 615486
rect 241840 615218 241882 615454
rect 242118 615218 242160 615454
rect 241840 615134 242160 615218
rect 241840 614898 241882 615134
rect 242118 614898 242160 615134
rect 241840 614866 242160 614898
rect 247771 615454 248091 615486
rect 247771 615218 247813 615454
rect 248049 615218 248091 615454
rect 247771 615134 248091 615218
rect 247771 614898 247813 615134
rect 248049 614898 248091 615134
rect 247771 614866 248091 614898
rect 262910 615454 263230 615486
rect 262910 615218 262952 615454
rect 263188 615218 263230 615454
rect 262910 615134 263230 615218
rect 262910 614898 262952 615134
rect 263188 614898 263230 615134
rect 262910 614866 263230 614898
rect 268840 615454 269160 615486
rect 268840 615218 268882 615454
rect 269118 615218 269160 615454
rect 268840 615134 269160 615218
rect 268840 614898 268882 615134
rect 269118 614898 269160 615134
rect 268840 614866 269160 614898
rect 274771 615454 275091 615486
rect 274771 615218 274813 615454
rect 275049 615218 275091 615454
rect 274771 615134 275091 615218
rect 274771 614898 274813 615134
rect 275049 614898 275091 615134
rect 274771 614866 275091 614898
rect 289910 615454 290230 615486
rect 289910 615218 289952 615454
rect 290188 615218 290230 615454
rect 289910 615134 290230 615218
rect 289910 614898 289952 615134
rect 290188 614898 290230 615134
rect 289910 614866 290230 614898
rect 295840 615454 296160 615486
rect 295840 615218 295882 615454
rect 296118 615218 296160 615454
rect 295840 615134 296160 615218
rect 295840 614898 295882 615134
rect 296118 614898 296160 615134
rect 295840 614866 296160 614898
rect 301771 615454 302091 615486
rect 301771 615218 301813 615454
rect 302049 615218 302091 615454
rect 301771 615134 302091 615218
rect 301771 614898 301813 615134
rect 302049 614898 302091 615134
rect 301771 614866 302091 614898
rect 316910 615454 317230 615486
rect 316910 615218 316952 615454
rect 317188 615218 317230 615454
rect 316910 615134 317230 615218
rect 316910 614898 316952 615134
rect 317188 614898 317230 615134
rect 316910 614866 317230 614898
rect 322840 615454 323160 615486
rect 322840 615218 322882 615454
rect 323118 615218 323160 615454
rect 322840 615134 323160 615218
rect 322840 614898 322882 615134
rect 323118 614898 323160 615134
rect 322840 614866 323160 614898
rect 328771 615454 329091 615486
rect 328771 615218 328813 615454
rect 329049 615218 329091 615454
rect 328771 615134 329091 615218
rect 328771 614898 328813 615134
rect 329049 614898 329091 615134
rect 328771 614866 329091 614898
rect 343910 615454 344230 615486
rect 343910 615218 343952 615454
rect 344188 615218 344230 615454
rect 343910 615134 344230 615218
rect 343910 614898 343952 615134
rect 344188 614898 344230 615134
rect 343910 614866 344230 614898
rect 349840 615454 350160 615486
rect 349840 615218 349882 615454
rect 350118 615218 350160 615454
rect 349840 615134 350160 615218
rect 349840 614898 349882 615134
rect 350118 614898 350160 615134
rect 349840 614866 350160 614898
rect 355771 615454 356091 615486
rect 355771 615218 355813 615454
rect 356049 615218 356091 615454
rect 355771 615134 356091 615218
rect 355771 614898 355813 615134
rect 356049 614898 356091 615134
rect 355771 614866 356091 614898
rect 370910 615454 371230 615486
rect 370910 615218 370952 615454
rect 371188 615218 371230 615454
rect 370910 615134 371230 615218
rect 370910 614898 370952 615134
rect 371188 614898 371230 615134
rect 370910 614866 371230 614898
rect 376840 615454 377160 615486
rect 376840 615218 376882 615454
rect 377118 615218 377160 615454
rect 376840 615134 377160 615218
rect 376840 614898 376882 615134
rect 377118 614898 377160 615134
rect 376840 614866 377160 614898
rect 382771 615454 383091 615486
rect 382771 615218 382813 615454
rect 383049 615218 383091 615454
rect 382771 615134 383091 615218
rect 382771 614898 382813 615134
rect 383049 614898 383091 615134
rect 382771 614866 383091 614898
rect 397910 615454 398230 615486
rect 397910 615218 397952 615454
rect 398188 615218 398230 615454
rect 397910 615134 398230 615218
rect 397910 614898 397952 615134
rect 398188 614898 398230 615134
rect 397910 614866 398230 614898
rect 403840 615454 404160 615486
rect 403840 615218 403882 615454
rect 404118 615218 404160 615454
rect 403840 615134 404160 615218
rect 403840 614898 403882 615134
rect 404118 614898 404160 615134
rect 403840 614866 404160 614898
rect 409771 615454 410091 615486
rect 409771 615218 409813 615454
rect 410049 615218 410091 615454
rect 409771 615134 410091 615218
rect 409771 614898 409813 615134
rect 410049 614898 410091 615134
rect 409771 614866 410091 614898
rect 424910 615454 425230 615486
rect 424910 615218 424952 615454
rect 425188 615218 425230 615454
rect 424910 615134 425230 615218
rect 424910 614898 424952 615134
rect 425188 614898 425230 615134
rect 424910 614866 425230 614898
rect 430840 615454 431160 615486
rect 430840 615218 430882 615454
rect 431118 615218 431160 615454
rect 430840 615134 431160 615218
rect 430840 614898 430882 615134
rect 431118 614898 431160 615134
rect 430840 614866 431160 614898
rect 436771 615454 437091 615486
rect 436771 615218 436813 615454
rect 437049 615218 437091 615454
rect 436771 615134 437091 615218
rect 436771 614898 436813 615134
rect 437049 614898 437091 615134
rect 436771 614866 437091 614898
rect 451910 615454 452230 615486
rect 451910 615218 451952 615454
rect 452188 615218 452230 615454
rect 451910 615134 452230 615218
rect 451910 614898 451952 615134
rect 452188 614898 452230 615134
rect 451910 614866 452230 614898
rect 457840 615454 458160 615486
rect 457840 615218 457882 615454
rect 458118 615218 458160 615454
rect 457840 615134 458160 615218
rect 457840 614898 457882 615134
rect 458118 614898 458160 615134
rect 457840 614866 458160 614898
rect 463771 615454 464091 615486
rect 463771 615218 463813 615454
rect 464049 615218 464091 615454
rect 463771 615134 464091 615218
rect 463771 614898 463813 615134
rect 464049 614898 464091 615134
rect 463771 614866 464091 614898
rect 478910 615454 479230 615486
rect 478910 615218 478952 615454
rect 479188 615218 479230 615454
rect 478910 615134 479230 615218
rect 478910 614898 478952 615134
rect 479188 614898 479230 615134
rect 478910 614866 479230 614898
rect 484840 615454 485160 615486
rect 484840 615218 484882 615454
rect 485118 615218 485160 615454
rect 484840 615134 485160 615218
rect 484840 614898 484882 615134
rect 485118 614898 485160 615134
rect 484840 614866 485160 614898
rect 490771 615454 491091 615486
rect 490771 615218 490813 615454
rect 491049 615218 491091 615454
rect 490771 615134 491091 615218
rect 490771 614898 490813 615134
rect 491049 614898 491091 615134
rect 490771 614866 491091 614898
rect 505910 615454 506230 615486
rect 505910 615218 505952 615454
rect 506188 615218 506230 615454
rect 505910 615134 506230 615218
rect 505910 614898 505952 615134
rect 506188 614898 506230 615134
rect 505910 614866 506230 614898
rect 511840 615454 512160 615486
rect 511840 615218 511882 615454
rect 512118 615218 512160 615454
rect 511840 615134 512160 615218
rect 511840 614898 511882 615134
rect 512118 614898 512160 615134
rect 511840 614866 512160 614898
rect 517771 615454 518091 615486
rect 517771 615218 517813 615454
rect 518049 615218 518091 615454
rect 517771 615134 518091 615218
rect 517771 614898 517813 615134
rect 518049 614898 518091 615134
rect 517771 614866 518091 614898
rect 532910 615454 533230 615486
rect 532910 615218 532952 615454
rect 533188 615218 533230 615454
rect 532910 615134 533230 615218
rect 532910 614898 532952 615134
rect 533188 614898 533230 615134
rect 532910 614866 533230 614898
rect 538840 615454 539160 615486
rect 538840 615218 538882 615454
rect 539118 615218 539160 615454
rect 538840 615134 539160 615218
rect 538840 614898 538882 615134
rect 539118 614898 539160 615134
rect 538840 614866 539160 614898
rect 544771 615454 545091 615486
rect 544771 615218 544813 615454
rect 545049 615218 545091 615454
rect 544771 615134 545091 615218
rect 544771 614898 544813 615134
rect 545049 614898 545091 615134
rect 544771 614866 545091 614898
rect 559794 615454 560414 632898
rect 559794 615218 559826 615454
rect 560062 615218 560146 615454
rect 560382 615218 560414 615454
rect 559794 615134 560414 615218
rect 559794 614898 559826 615134
rect 560062 614898 560146 615134
rect 560382 614898 560414 615134
rect 10794 606218 10826 606454
rect 11062 606218 11146 606454
rect 11382 606218 11414 606454
rect 10794 606134 11414 606218
rect 10794 605898 10826 606134
rect 11062 605898 11146 606134
rect 11382 605898 11414 606134
rect 10794 588454 11414 605898
rect 19794 607394 20414 608000
rect 19794 607158 19826 607394
rect 20062 607158 20146 607394
rect 20382 607158 20414 607394
rect 19794 607074 20414 607158
rect 19794 606838 19826 607074
rect 20062 606838 20146 607074
rect 20382 606838 20414 607074
rect 19794 605000 20414 606838
rect 28794 606454 29414 608000
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 605000 29414 605898
rect 37794 607394 38414 608000
rect 37794 607158 37826 607394
rect 38062 607158 38146 607394
rect 38382 607158 38414 607394
rect 37794 607074 38414 607158
rect 37794 606838 37826 607074
rect 38062 606838 38146 607074
rect 38382 606838 38414 607074
rect 37794 605000 38414 606838
rect 46794 606454 47414 608000
rect 46794 606218 46826 606454
rect 47062 606218 47146 606454
rect 47382 606218 47414 606454
rect 46794 606134 47414 606218
rect 46794 605898 46826 606134
rect 47062 605898 47146 606134
rect 47382 605898 47414 606134
rect 46794 605000 47414 605898
rect 55794 607394 56414 608000
rect 55794 607158 55826 607394
rect 56062 607158 56146 607394
rect 56382 607158 56414 607394
rect 55794 607074 56414 607158
rect 55794 606838 55826 607074
rect 56062 606838 56146 607074
rect 56382 606838 56414 607074
rect 55794 605000 56414 606838
rect 64794 606454 65414 608000
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 605000 65414 605898
rect 73794 607394 74414 608000
rect 73794 607158 73826 607394
rect 74062 607158 74146 607394
rect 74382 607158 74414 607394
rect 73794 607074 74414 607158
rect 73794 606838 73826 607074
rect 74062 606838 74146 607074
rect 74382 606838 74414 607074
rect 73794 605000 74414 606838
rect 82794 606454 83414 608000
rect 82794 606218 82826 606454
rect 83062 606218 83146 606454
rect 83382 606218 83414 606454
rect 82794 606134 83414 606218
rect 82794 605898 82826 606134
rect 83062 605898 83146 606134
rect 83382 605898 83414 606134
rect 82794 605000 83414 605898
rect 91794 607394 92414 608000
rect 91794 607158 91826 607394
rect 92062 607158 92146 607394
rect 92382 607158 92414 607394
rect 91794 607074 92414 607158
rect 91794 606838 91826 607074
rect 92062 606838 92146 607074
rect 92382 606838 92414 607074
rect 91794 605000 92414 606838
rect 100794 606454 101414 608000
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 605000 101414 605898
rect 109794 607394 110414 608000
rect 109794 607158 109826 607394
rect 110062 607158 110146 607394
rect 110382 607158 110414 607394
rect 109794 607074 110414 607158
rect 109794 606838 109826 607074
rect 110062 606838 110146 607074
rect 110382 606838 110414 607074
rect 109794 605000 110414 606838
rect 118794 606454 119414 608000
rect 118794 606218 118826 606454
rect 119062 606218 119146 606454
rect 119382 606218 119414 606454
rect 118794 606134 119414 606218
rect 118794 605898 118826 606134
rect 119062 605898 119146 606134
rect 119382 605898 119414 606134
rect 118794 605000 119414 605898
rect 127794 607394 128414 608000
rect 127794 607158 127826 607394
rect 128062 607158 128146 607394
rect 128382 607158 128414 607394
rect 127794 607074 128414 607158
rect 127794 606838 127826 607074
rect 128062 606838 128146 607074
rect 128382 606838 128414 607074
rect 127794 605000 128414 606838
rect 136794 606454 137414 608000
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 605000 137414 605898
rect 145794 607394 146414 608000
rect 145794 607158 145826 607394
rect 146062 607158 146146 607394
rect 146382 607158 146414 607394
rect 145794 607074 146414 607158
rect 145794 606838 145826 607074
rect 146062 606838 146146 607074
rect 146382 606838 146414 607074
rect 145794 605000 146414 606838
rect 154794 606454 155414 608000
rect 154794 606218 154826 606454
rect 155062 606218 155146 606454
rect 155382 606218 155414 606454
rect 154794 606134 155414 606218
rect 154794 605898 154826 606134
rect 155062 605898 155146 606134
rect 155382 605898 155414 606134
rect 154794 605000 155414 605898
rect 163794 607394 164414 608000
rect 163794 607158 163826 607394
rect 164062 607158 164146 607394
rect 164382 607158 164414 607394
rect 163794 607074 164414 607158
rect 163794 606838 163826 607074
rect 164062 606838 164146 607074
rect 164382 606838 164414 607074
rect 163794 605000 164414 606838
rect 172794 606454 173414 608000
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 605000 173414 605898
rect 181794 607394 182414 608000
rect 181794 607158 181826 607394
rect 182062 607158 182146 607394
rect 182382 607158 182414 607394
rect 181794 607074 182414 607158
rect 181794 606838 181826 607074
rect 182062 606838 182146 607074
rect 182382 606838 182414 607074
rect 181794 605000 182414 606838
rect 190794 606454 191414 608000
rect 190794 606218 190826 606454
rect 191062 606218 191146 606454
rect 191382 606218 191414 606454
rect 190794 606134 191414 606218
rect 190794 605898 190826 606134
rect 191062 605898 191146 606134
rect 191382 605898 191414 606134
rect 190794 605000 191414 605898
rect 199794 607394 200414 608000
rect 199794 607158 199826 607394
rect 200062 607158 200146 607394
rect 200382 607158 200414 607394
rect 199794 607074 200414 607158
rect 199794 606838 199826 607074
rect 200062 606838 200146 607074
rect 200382 606838 200414 607074
rect 199794 605000 200414 606838
rect 208794 606454 209414 608000
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 605000 209414 605898
rect 217794 607394 218414 608000
rect 217794 607158 217826 607394
rect 218062 607158 218146 607394
rect 218382 607158 218414 607394
rect 217794 607074 218414 607158
rect 217794 606838 217826 607074
rect 218062 606838 218146 607074
rect 218382 606838 218414 607074
rect 217794 605000 218414 606838
rect 226794 606454 227414 608000
rect 226794 606218 226826 606454
rect 227062 606218 227146 606454
rect 227382 606218 227414 606454
rect 226794 606134 227414 606218
rect 226794 605898 226826 606134
rect 227062 605898 227146 606134
rect 227382 605898 227414 606134
rect 226794 605000 227414 605898
rect 235794 607394 236414 608000
rect 235794 607158 235826 607394
rect 236062 607158 236146 607394
rect 236382 607158 236414 607394
rect 235794 607074 236414 607158
rect 235794 606838 235826 607074
rect 236062 606838 236146 607074
rect 236382 606838 236414 607074
rect 235794 605000 236414 606838
rect 244794 606454 245414 608000
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 605000 245414 605898
rect 253794 607394 254414 608000
rect 253794 607158 253826 607394
rect 254062 607158 254146 607394
rect 254382 607158 254414 607394
rect 253794 607074 254414 607158
rect 253794 606838 253826 607074
rect 254062 606838 254146 607074
rect 254382 606838 254414 607074
rect 253794 605000 254414 606838
rect 262794 606454 263414 608000
rect 262794 606218 262826 606454
rect 263062 606218 263146 606454
rect 263382 606218 263414 606454
rect 262794 606134 263414 606218
rect 262794 605898 262826 606134
rect 263062 605898 263146 606134
rect 263382 605898 263414 606134
rect 262794 605000 263414 605898
rect 271794 607394 272414 608000
rect 271794 607158 271826 607394
rect 272062 607158 272146 607394
rect 272382 607158 272414 607394
rect 271794 607074 272414 607158
rect 271794 606838 271826 607074
rect 272062 606838 272146 607074
rect 272382 606838 272414 607074
rect 271794 605000 272414 606838
rect 280794 606454 281414 608000
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 605000 281414 605898
rect 289794 607394 290414 608000
rect 289794 607158 289826 607394
rect 290062 607158 290146 607394
rect 290382 607158 290414 607394
rect 289794 607074 290414 607158
rect 289794 606838 289826 607074
rect 290062 606838 290146 607074
rect 290382 606838 290414 607074
rect 289794 605000 290414 606838
rect 298794 606454 299414 608000
rect 298794 606218 298826 606454
rect 299062 606218 299146 606454
rect 299382 606218 299414 606454
rect 298794 606134 299414 606218
rect 298794 605898 298826 606134
rect 299062 605898 299146 606134
rect 299382 605898 299414 606134
rect 298794 605000 299414 605898
rect 307794 607394 308414 608000
rect 307794 607158 307826 607394
rect 308062 607158 308146 607394
rect 308382 607158 308414 607394
rect 307794 607074 308414 607158
rect 307794 606838 307826 607074
rect 308062 606838 308146 607074
rect 308382 606838 308414 607074
rect 307794 605000 308414 606838
rect 316794 606454 317414 608000
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 605000 317414 605898
rect 325794 607394 326414 608000
rect 325794 607158 325826 607394
rect 326062 607158 326146 607394
rect 326382 607158 326414 607394
rect 325794 607074 326414 607158
rect 325794 606838 325826 607074
rect 326062 606838 326146 607074
rect 326382 606838 326414 607074
rect 325794 605000 326414 606838
rect 334794 606454 335414 608000
rect 334794 606218 334826 606454
rect 335062 606218 335146 606454
rect 335382 606218 335414 606454
rect 334794 606134 335414 606218
rect 334794 605898 334826 606134
rect 335062 605898 335146 606134
rect 335382 605898 335414 606134
rect 334794 605000 335414 605898
rect 343794 607394 344414 608000
rect 343794 607158 343826 607394
rect 344062 607158 344146 607394
rect 344382 607158 344414 607394
rect 343794 607074 344414 607158
rect 343794 606838 343826 607074
rect 344062 606838 344146 607074
rect 344382 606838 344414 607074
rect 343794 605000 344414 606838
rect 352794 606454 353414 608000
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 605000 353414 605898
rect 361794 607394 362414 608000
rect 361794 607158 361826 607394
rect 362062 607158 362146 607394
rect 362382 607158 362414 607394
rect 361794 607074 362414 607158
rect 361794 606838 361826 607074
rect 362062 606838 362146 607074
rect 362382 606838 362414 607074
rect 361794 605000 362414 606838
rect 370794 606454 371414 608000
rect 370794 606218 370826 606454
rect 371062 606218 371146 606454
rect 371382 606218 371414 606454
rect 370794 606134 371414 606218
rect 370794 605898 370826 606134
rect 371062 605898 371146 606134
rect 371382 605898 371414 606134
rect 370794 605000 371414 605898
rect 379794 607394 380414 608000
rect 379794 607158 379826 607394
rect 380062 607158 380146 607394
rect 380382 607158 380414 607394
rect 379794 607074 380414 607158
rect 379794 606838 379826 607074
rect 380062 606838 380146 607074
rect 380382 606838 380414 607074
rect 379794 605000 380414 606838
rect 388794 606454 389414 608000
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 605000 389414 605898
rect 397794 607394 398414 608000
rect 397794 607158 397826 607394
rect 398062 607158 398146 607394
rect 398382 607158 398414 607394
rect 397794 607074 398414 607158
rect 397794 606838 397826 607074
rect 398062 606838 398146 607074
rect 398382 606838 398414 607074
rect 397794 605000 398414 606838
rect 406794 606454 407414 608000
rect 406794 606218 406826 606454
rect 407062 606218 407146 606454
rect 407382 606218 407414 606454
rect 406794 606134 407414 606218
rect 406794 605898 406826 606134
rect 407062 605898 407146 606134
rect 407382 605898 407414 606134
rect 406794 605000 407414 605898
rect 415794 607394 416414 608000
rect 415794 607158 415826 607394
rect 416062 607158 416146 607394
rect 416382 607158 416414 607394
rect 415794 607074 416414 607158
rect 415794 606838 415826 607074
rect 416062 606838 416146 607074
rect 416382 606838 416414 607074
rect 415794 605000 416414 606838
rect 424794 606454 425414 608000
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 605000 425414 605898
rect 433794 607394 434414 608000
rect 433794 607158 433826 607394
rect 434062 607158 434146 607394
rect 434382 607158 434414 607394
rect 433794 607074 434414 607158
rect 433794 606838 433826 607074
rect 434062 606838 434146 607074
rect 434382 606838 434414 607074
rect 433794 605000 434414 606838
rect 442794 606454 443414 608000
rect 442794 606218 442826 606454
rect 443062 606218 443146 606454
rect 443382 606218 443414 606454
rect 442794 606134 443414 606218
rect 442794 605898 442826 606134
rect 443062 605898 443146 606134
rect 443382 605898 443414 606134
rect 442794 605000 443414 605898
rect 451794 607394 452414 608000
rect 451794 607158 451826 607394
rect 452062 607158 452146 607394
rect 452382 607158 452414 607394
rect 451794 607074 452414 607158
rect 451794 606838 451826 607074
rect 452062 606838 452146 607074
rect 452382 606838 452414 607074
rect 451794 605000 452414 606838
rect 460794 606454 461414 608000
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 605000 461414 605898
rect 469794 607394 470414 608000
rect 469794 607158 469826 607394
rect 470062 607158 470146 607394
rect 470382 607158 470414 607394
rect 469794 607074 470414 607158
rect 469794 606838 469826 607074
rect 470062 606838 470146 607074
rect 470382 606838 470414 607074
rect 469794 605000 470414 606838
rect 478794 606454 479414 608000
rect 478794 606218 478826 606454
rect 479062 606218 479146 606454
rect 479382 606218 479414 606454
rect 478794 606134 479414 606218
rect 478794 605898 478826 606134
rect 479062 605898 479146 606134
rect 479382 605898 479414 606134
rect 478794 605000 479414 605898
rect 487794 607394 488414 608000
rect 487794 607158 487826 607394
rect 488062 607158 488146 607394
rect 488382 607158 488414 607394
rect 487794 607074 488414 607158
rect 487794 606838 487826 607074
rect 488062 606838 488146 607074
rect 488382 606838 488414 607074
rect 487794 605000 488414 606838
rect 496794 606454 497414 608000
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 605000 497414 605898
rect 505794 607394 506414 608000
rect 505794 607158 505826 607394
rect 506062 607158 506146 607394
rect 506382 607158 506414 607394
rect 505794 607074 506414 607158
rect 505794 606838 505826 607074
rect 506062 606838 506146 607074
rect 506382 606838 506414 607074
rect 505794 605000 506414 606838
rect 514794 606454 515414 608000
rect 514794 606218 514826 606454
rect 515062 606218 515146 606454
rect 515382 606218 515414 606454
rect 514794 606134 515414 606218
rect 514794 605898 514826 606134
rect 515062 605898 515146 606134
rect 515382 605898 515414 606134
rect 514794 605000 515414 605898
rect 523794 607394 524414 608000
rect 523794 607158 523826 607394
rect 524062 607158 524146 607394
rect 524382 607158 524414 607394
rect 523794 607074 524414 607158
rect 523794 606838 523826 607074
rect 524062 606838 524146 607074
rect 524382 606838 524414 607074
rect 523794 605000 524414 606838
rect 532794 606454 533414 608000
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 605000 533414 605898
rect 541794 607394 542414 608000
rect 541794 607158 541826 607394
rect 542062 607158 542146 607394
rect 542382 607158 542414 607394
rect 541794 607074 542414 607158
rect 541794 606838 541826 607074
rect 542062 606838 542146 607074
rect 542382 606838 542414 607074
rect 541794 605000 542414 606838
rect 550794 606454 551414 608000
rect 550794 606218 550826 606454
rect 551062 606218 551146 606454
rect 551382 606218 551414 606454
rect 550794 606134 551414 606218
rect 550794 605898 550826 606134
rect 551062 605898 551146 606134
rect 551382 605898 551414 606134
rect 550794 605000 551414 605898
rect 19910 597454 20230 597486
rect 19910 597218 19952 597454
rect 20188 597218 20230 597454
rect 19910 597134 20230 597218
rect 19910 596898 19952 597134
rect 20188 596898 20230 597134
rect 19910 596866 20230 596898
rect 25840 597454 26160 597486
rect 25840 597218 25882 597454
rect 26118 597218 26160 597454
rect 25840 597134 26160 597218
rect 25840 596898 25882 597134
rect 26118 596898 26160 597134
rect 25840 596866 26160 596898
rect 31771 597454 32091 597486
rect 31771 597218 31813 597454
rect 32049 597218 32091 597454
rect 31771 597134 32091 597218
rect 31771 596898 31813 597134
rect 32049 596898 32091 597134
rect 31771 596866 32091 596898
rect 46910 597454 47230 597486
rect 46910 597218 46952 597454
rect 47188 597218 47230 597454
rect 46910 597134 47230 597218
rect 46910 596898 46952 597134
rect 47188 596898 47230 597134
rect 46910 596866 47230 596898
rect 52840 597454 53160 597486
rect 52840 597218 52882 597454
rect 53118 597218 53160 597454
rect 52840 597134 53160 597218
rect 52840 596898 52882 597134
rect 53118 596898 53160 597134
rect 52840 596866 53160 596898
rect 58771 597454 59091 597486
rect 58771 597218 58813 597454
rect 59049 597218 59091 597454
rect 58771 597134 59091 597218
rect 58771 596898 58813 597134
rect 59049 596898 59091 597134
rect 58771 596866 59091 596898
rect 73910 597454 74230 597486
rect 73910 597218 73952 597454
rect 74188 597218 74230 597454
rect 73910 597134 74230 597218
rect 73910 596898 73952 597134
rect 74188 596898 74230 597134
rect 73910 596866 74230 596898
rect 79840 597454 80160 597486
rect 79840 597218 79882 597454
rect 80118 597218 80160 597454
rect 79840 597134 80160 597218
rect 79840 596898 79882 597134
rect 80118 596898 80160 597134
rect 79840 596866 80160 596898
rect 85771 597454 86091 597486
rect 85771 597218 85813 597454
rect 86049 597218 86091 597454
rect 85771 597134 86091 597218
rect 85771 596898 85813 597134
rect 86049 596898 86091 597134
rect 85771 596866 86091 596898
rect 100910 597454 101230 597486
rect 100910 597218 100952 597454
rect 101188 597218 101230 597454
rect 100910 597134 101230 597218
rect 100910 596898 100952 597134
rect 101188 596898 101230 597134
rect 100910 596866 101230 596898
rect 106840 597454 107160 597486
rect 106840 597218 106882 597454
rect 107118 597218 107160 597454
rect 106840 597134 107160 597218
rect 106840 596898 106882 597134
rect 107118 596898 107160 597134
rect 106840 596866 107160 596898
rect 112771 597454 113091 597486
rect 112771 597218 112813 597454
rect 113049 597218 113091 597454
rect 112771 597134 113091 597218
rect 112771 596898 112813 597134
rect 113049 596898 113091 597134
rect 112771 596866 113091 596898
rect 127910 597454 128230 597486
rect 127910 597218 127952 597454
rect 128188 597218 128230 597454
rect 127910 597134 128230 597218
rect 127910 596898 127952 597134
rect 128188 596898 128230 597134
rect 127910 596866 128230 596898
rect 133840 597454 134160 597486
rect 133840 597218 133882 597454
rect 134118 597218 134160 597454
rect 133840 597134 134160 597218
rect 133840 596898 133882 597134
rect 134118 596898 134160 597134
rect 133840 596866 134160 596898
rect 139771 597454 140091 597486
rect 139771 597218 139813 597454
rect 140049 597218 140091 597454
rect 139771 597134 140091 597218
rect 139771 596898 139813 597134
rect 140049 596898 140091 597134
rect 139771 596866 140091 596898
rect 154910 597454 155230 597486
rect 154910 597218 154952 597454
rect 155188 597218 155230 597454
rect 154910 597134 155230 597218
rect 154910 596898 154952 597134
rect 155188 596898 155230 597134
rect 154910 596866 155230 596898
rect 160840 597454 161160 597486
rect 160840 597218 160882 597454
rect 161118 597218 161160 597454
rect 160840 597134 161160 597218
rect 160840 596898 160882 597134
rect 161118 596898 161160 597134
rect 160840 596866 161160 596898
rect 166771 597454 167091 597486
rect 166771 597218 166813 597454
rect 167049 597218 167091 597454
rect 166771 597134 167091 597218
rect 166771 596898 166813 597134
rect 167049 596898 167091 597134
rect 166771 596866 167091 596898
rect 181910 597454 182230 597486
rect 181910 597218 181952 597454
rect 182188 597218 182230 597454
rect 181910 597134 182230 597218
rect 181910 596898 181952 597134
rect 182188 596898 182230 597134
rect 181910 596866 182230 596898
rect 187840 597454 188160 597486
rect 187840 597218 187882 597454
rect 188118 597218 188160 597454
rect 187840 597134 188160 597218
rect 187840 596898 187882 597134
rect 188118 596898 188160 597134
rect 187840 596866 188160 596898
rect 193771 597454 194091 597486
rect 193771 597218 193813 597454
rect 194049 597218 194091 597454
rect 193771 597134 194091 597218
rect 193771 596898 193813 597134
rect 194049 596898 194091 597134
rect 193771 596866 194091 596898
rect 208910 597454 209230 597486
rect 208910 597218 208952 597454
rect 209188 597218 209230 597454
rect 208910 597134 209230 597218
rect 208910 596898 208952 597134
rect 209188 596898 209230 597134
rect 208910 596866 209230 596898
rect 214840 597454 215160 597486
rect 214840 597218 214882 597454
rect 215118 597218 215160 597454
rect 214840 597134 215160 597218
rect 214840 596898 214882 597134
rect 215118 596898 215160 597134
rect 214840 596866 215160 596898
rect 220771 597454 221091 597486
rect 220771 597218 220813 597454
rect 221049 597218 221091 597454
rect 220771 597134 221091 597218
rect 220771 596898 220813 597134
rect 221049 596898 221091 597134
rect 220771 596866 221091 596898
rect 235910 597454 236230 597486
rect 235910 597218 235952 597454
rect 236188 597218 236230 597454
rect 235910 597134 236230 597218
rect 235910 596898 235952 597134
rect 236188 596898 236230 597134
rect 235910 596866 236230 596898
rect 241840 597454 242160 597486
rect 241840 597218 241882 597454
rect 242118 597218 242160 597454
rect 241840 597134 242160 597218
rect 241840 596898 241882 597134
rect 242118 596898 242160 597134
rect 241840 596866 242160 596898
rect 247771 597454 248091 597486
rect 247771 597218 247813 597454
rect 248049 597218 248091 597454
rect 247771 597134 248091 597218
rect 247771 596898 247813 597134
rect 248049 596898 248091 597134
rect 247771 596866 248091 596898
rect 262910 597454 263230 597486
rect 262910 597218 262952 597454
rect 263188 597218 263230 597454
rect 262910 597134 263230 597218
rect 262910 596898 262952 597134
rect 263188 596898 263230 597134
rect 262910 596866 263230 596898
rect 268840 597454 269160 597486
rect 268840 597218 268882 597454
rect 269118 597218 269160 597454
rect 268840 597134 269160 597218
rect 268840 596898 268882 597134
rect 269118 596898 269160 597134
rect 268840 596866 269160 596898
rect 274771 597454 275091 597486
rect 274771 597218 274813 597454
rect 275049 597218 275091 597454
rect 274771 597134 275091 597218
rect 274771 596898 274813 597134
rect 275049 596898 275091 597134
rect 274771 596866 275091 596898
rect 289910 597454 290230 597486
rect 289910 597218 289952 597454
rect 290188 597218 290230 597454
rect 289910 597134 290230 597218
rect 289910 596898 289952 597134
rect 290188 596898 290230 597134
rect 289910 596866 290230 596898
rect 295840 597454 296160 597486
rect 295840 597218 295882 597454
rect 296118 597218 296160 597454
rect 295840 597134 296160 597218
rect 295840 596898 295882 597134
rect 296118 596898 296160 597134
rect 295840 596866 296160 596898
rect 301771 597454 302091 597486
rect 301771 597218 301813 597454
rect 302049 597218 302091 597454
rect 301771 597134 302091 597218
rect 301771 596898 301813 597134
rect 302049 596898 302091 597134
rect 301771 596866 302091 596898
rect 316910 597454 317230 597486
rect 316910 597218 316952 597454
rect 317188 597218 317230 597454
rect 316910 597134 317230 597218
rect 316910 596898 316952 597134
rect 317188 596898 317230 597134
rect 316910 596866 317230 596898
rect 322840 597454 323160 597486
rect 322840 597218 322882 597454
rect 323118 597218 323160 597454
rect 322840 597134 323160 597218
rect 322840 596898 322882 597134
rect 323118 596898 323160 597134
rect 322840 596866 323160 596898
rect 328771 597454 329091 597486
rect 328771 597218 328813 597454
rect 329049 597218 329091 597454
rect 328771 597134 329091 597218
rect 328771 596898 328813 597134
rect 329049 596898 329091 597134
rect 328771 596866 329091 596898
rect 343910 597454 344230 597486
rect 343910 597218 343952 597454
rect 344188 597218 344230 597454
rect 343910 597134 344230 597218
rect 343910 596898 343952 597134
rect 344188 596898 344230 597134
rect 343910 596866 344230 596898
rect 349840 597454 350160 597486
rect 349840 597218 349882 597454
rect 350118 597218 350160 597454
rect 349840 597134 350160 597218
rect 349840 596898 349882 597134
rect 350118 596898 350160 597134
rect 349840 596866 350160 596898
rect 355771 597454 356091 597486
rect 355771 597218 355813 597454
rect 356049 597218 356091 597454
rect 355771 597134 356091 597218
rect 355771 596898 355813 597134
rect 356049 596898 356091 597134
rect 355771 596866 356091 596898
rect 370910 597454 371230 597486
rect 370910 597218 370952 597454
rect 371188 597218 371230 597454
rect 370910 597134 371230 597218
rect 370910 596898 370952 597134
rect 371188 596898 371230 597134
rect 370910 596866 371230 596898
rect 376840 597454 377160 597486
rect 376840 597218 376882 597454
rect 377118 597218 377160 597454
rect 376840 597134 377160 597218
rect 376840 596898 376882 597134
rect 377118 596898 377160 597134
rect 376840 596866 377160 596898
rect 382771 597454 383091 597486
rect 382771 597218 382813 597454
rect 383049 597218 383091 597454
rect 382771 597134 383091 597218
rect 382771 596898 382813 597134
rect 383049 596898 383091 597134
rect 382771 596866 383091 596898
rect 397910 597454 398230 597486
rect 397910 597218 397952 597454
rect 398188 597218 398230 597454
rect 397910 597134 398230 597218
rect 397910 596898 397952 597134
rect 398188 596898 398230 597134
rect 397910 596866 398230 596898
rect 403840 597454 404160 597486
rect 403840 597218 403882 597454
rect 404118 597218 404160 597454
rect 403840 597134 404160 597218
rect 403840 596898 403882 597134
rect 404118 596898 404160 597134
rect 403840 596866 404160 596898
rect 409771 597454 410091 597486
rect 409771 597218 409813 597454
rect 410049 597218 410091 597454
rect 409771 597134 410091 597218
rect 409771 596898 409813 597134
rect 410049 596898 410091 597134
rect 409771 596866 410091 596898
rect 424910 597454 425230 597486
rect 424910 597218 424952 597454
rect 425188 597218 425230 597454
rect 424910 597134 425230 597218
rect 424910 596898 424952 597134
rect 425188 596898 425230 597134
rect 424910 596866 425230 596898
rect 430840 597454 431160 597486
rect 430840 597218 430882 597454
rect 431118 597218 431160 597454
rect 430840 597134 431160 597218
rect 430840 596898 430882 597134
rect 431118 596898 431160 597134
rect 430840 596866 431160 596898
rect 436771 597454 437091 597486
rect 436771 597218 436813 597454
rect 437049 597218 437091 597454
rect 436771 597134 437091 597218
rect 436771 596898 436813 597134
rect 437049 596898 437091 597134
rect 436771 596866 437091 596898
rect 451910 597454 452230 597486
rect 451910 597218 451952 597454
rect 452188 597218 452230 597454
rect 451910 597134 452230 597218
rect 451910 596898 451952 597134
rect 452188 596898 452230 597134
rect 451910 596866 452230 596898
rect 457840 597454 458160 597486
rect 457840 597218 457882 597454
rect 458118 597218 458160 597454
rect 457840 597134 458160 597218
rect 457840 596898 457882 597134
rect 458118 596898 458160 597134
rect 457840 596866 458160 596898
rect 463771 597454 464091 597486
rect 463771 597218 463813 597454
rect 464049 597218 464091 597454
rect 463771 597134 464091 597218
rect 463771 596898 463813 597134
rect 464049 596898 464091 597134
rect 463771 596866 464091 596898
rect 478910 597454 479230 597486
rect 478910 597218 478952 597454
rect 479188 597218 479230 597454
rect 478910 597134 479230 597218
rect 478910 596898 478952 597134
rect 479188 596898 479230 597134
rect 478910 596866 479230 596898
rect 484840 597454 485160 597486
rect 484840 597218 484882 597454
rect 485118 597218 485160 597454
rect 484840 597134 485160 597218
rect 484840 596898 484882 597134
rect 485118 596898 485160 597134
rect 484840 596866 485160 596898
rect 490771 597454 491091 597486
rect 490771 597218 490813 597454
rect 491049 597218 491091 597454
rect 490771 597134 491091 597218
rect 490771 596898 490813 597134
rect 491049 596898 491091 597134
rect 490771 596866 491091 596898
rect 505910 597454 506230 597486
rect 505910 597218 505952 597454
rect 506188 597218 506230 597454
rect 505910 597134 506230 597218
rect 505910 596898 505952 597134
rect 506188 596898 506230 597134
rect 505910 596866 506230 596898
rect 511840 597454 512160 597486
rect 511840 597218 511882 597454
rect 512118 597218 512160 597454
rect 511840 597134 512160 597218
rect 511840 596898 511882 597134
rect 512118 596898 512160 597134
rect 511840 596866 512160 596898
rect 517771 597454 518091 597486
rect 517771 597218 517813 597454
rect 518049 597218 518091 597454
rect 517771 597134 518091 597218
rect 517771 596898 517813 597134
rect 518049 596898 518091 597134
rect 517771 596866 518091 596898
rect 532910 597454 533230 597486
rect 532910 597218 532952 597454
rect 533188 597218 533230 597454
rect 532910 597134 533230 597218
rect 532910 596898 532952 597134
rect 533188 596898 533230 597134
rect 532910 596866 533230 596898
rect 538840 597454 539160 597486
rect 538840 597218 538882 597454
rect 539118 597218 539160 597454
rect 538840 597134 539160 597218
rect 538840 596898 538882 597134
rect 539118 596898 539160 597134
rect 538840 596866 539160 596898
rect 544771 597454 545091 597486
rect 544771 597218 544813 597454
rect 545049 597218 545091 597454
rect 544771 597134 545091 597218
rect 544771 596898 544813 597134
rect 545049 596898 545091 597134
rect 544771 596866 545091 596898
rect 559794 597454 560414 614898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 570454 11414 587898
rect 22874 588454 23194 588486
rect 22874 588218 22916 588454
rect 23152 588218 23194 588454
rect 22874 588134 23194 588218
rect 22874 587898 22916 588134
rect 23152 587898 23194 588134
rect 22874 587866 23194 587898
rect 28805 588454 29125 588486
rect 28805 588218 28847 588454
rect 29083 588218 29125 588454
rect 28805 588134 29125 588218
rect 28805 587898 28847 588134
rect 29083 587898 29125 588134
rect 28805 587866 29125 587898
rect 49874 588454 50194 588486
rect 49874 588218 49916 588454
rect 50152 588218 50194 588454
rect 49874 588134 50194 588218
rect 49874 587898 49916 588134
rect 50152 587898 50194 588134
rect 49874 587866 50194 587898
rect 55805 588454 56125 588486
rect 55805 588218 55847 588454
rect 56083 588218 56125 588454
rect 55805 588134 56125 588218
rect 55805 587898 55847 588134
rect 56083 587898 56125 588134
rect 55805 587866 56125 587898
rect 76874 588454 77194 588486
rect 76874 588218 76916 588454
rect 77152 588218 77194 588454
rect 76874 588134 77194 588218
rect 76874 587898 76916 588134
rect 77152 587898 77194 588134
rect 76874 587866 77194 587898
rect 82805 588454 83125 588486
rect 82805 588218 82847 588454
rect 83083 588218 83125 588454
rect 82805 588134 83125 588218
rect 82805 587898 82847 588134
rect 83083 587898 83125 588134
rect 82805 587866 83125 587898
rect 103874 588454 104194 588486
rect 103874 588218 103916 588454
rect 104152 588218 104194 588454
rect 103874 588134 104194 588218
rect 103874 587898 103916 588134
rect 104152 587898 104194 588134
rect 103874 587866 104194 587898
rect 109805 588454 110125 588486
rect 109805 588218 109847 588454
rect 110083 588218 110125 588454
rect 109805 588134 110125 588218
rect 109805 587898 109847 588134
rect 110083 587898 110125 588134
rect 109805 587866 110125 587898
rect 130874 588454 131194 588486
rect 130874 588218 130916 588454
rect 131152 588218 131194 588454
rect 130874 588134 131194 588218
rect 130874 587898 130916 588134
rect 131152 587898 131194 588134
rect 130874 587866 131194 587898
rect 136805 588454 137125 588486
rect 136805 588218 136847 588454
rect 137083 588218 137125 588454
rect 136805 588134 137125 588218
rect 136805 587898 136847 588134
rect 137083 587898 137125 588134
rect 136805 587866 137125 587898
rect 157874 588454 158194 588486
rect 157874 588218 157916 588454
rect 158152 588218 158194 588454
rect 157874 588134 158194 588218
rect 157874 587898 157916 588134
rect 158152 587898 158194 588134
rect 157874 587866 158194 587898
rect 163805 588454 164125 588486
rect 163805 588218 163847 588454
rect 164083 588218 164125 588454
rect 163805 588134 164125 588218
rect 163805 587898 163847 588134
rect 164083 587898 164125 588134
rect 163805 587866 164125 587898
rect 184874 588454 185194 588486
rect 184874 588218 184916 588454
rect 185152 588218 185194 588454
rect 184874 588134 185194 588218
rect 184874 587898 184916 588134
rect 185152 587898 185194 588134
rect 184874 587866 185194 587898
rect 190805 588454 191125 588486
rect 190805 588218 190847 588454
rect 191083 588218 191125 588454
rect 190805 588134 191125 588218
rect 190805 587898 190847 588134
rect 191083 587898 191125 588134
rect 190805 587866 191125 587898
rect 211874 588454 212194 588486
rect 211874 588218 211916 588454
rect 212152 588218 212194 588454
rect 211874 588134 212194 588218
rect 211874 587898 211916 588134
rect 212152 587898 212194 588134
rect 211874 587866 212194 587898
rect 217805 588454 218125 588486
rect 217805 588218 217847 588454
rect 218083 588218 218125 588454
rect 217805 588134 218125 588218
rect 217805 587898 217847 588134
rect 218083 587898 218125 588134
rect 217805 587866 218125 587898
rect 238874 588454 239194 588486
rect 238874 588218 238916 588454
rect 239152 588218 239194 588454
rect 238874 588134 239194 588218
rect 238874 587898 238916 588134
rect 239152 587898 239194 588134
rect 238874 587866 239194 587898
rect 244805 588454 245125 588486
rect 244805 588218 244847 588454
rect 245083 588218 245125 588454
rect 244805 588134 245125 588218
rect 244805 587898 244847 588134
rect 245083 587898 245125 588134
rect 244805 587866 245125 587898
rect 265874 588454 266194 588486
rect 265874 588218 265916 588454
rect 266152 588218 266194 588454
rect 265874 588134 266194 588218
rect 265874 587898 265916 588134
rect 266152 587898 266194 588134
rect 265874 587866 266194 587898
rect 271805 588454 272125 588486
rect 271805 588218 271847 588454
rect 272083 588218 272125 588454
rect 271805 588134 272125 588218
rect 271805 587898 271847 588134
rect 272083 587898 272125 588134
rect 271805 587866 272125 587898
rect 292874 588454 293194 588486
rect 292874 588218 292916 588454
rect 293152 588218 293194 588454
rect 292874 588134 293194 588218
rect 292874 587898 292916 588134
rect 293152 587898 293194 588134
rect 292874 587866 293194 587898
rect 298805 588454 299125 588486
rect 298805 588218 298847 588454
rect 299083 588218 299125 588454
rect 298805 588134 299125 588218
rect 298805 587898 298847 588134
rect 299083 587898 299125 588134
rect 298805 587866 299125 587898
rect 319874 588454 320194 588486
rect 319874 588218 319916 588454
rect 320152 588218 320194 588454
rect 319874 588134 320194 588218
rect 319874 587898 319916 588134
rect 320152 587898 320194 588134
rect 319874 587866 320194 587898
rect 325805 588454 326125 588486
rect 325805 588218 325847 588454
rect 326083 588218 326125 588454
rect 325805 588134 326125 588218
rect 325805 587898 325847 588134
rect 326083 587898 326125 588134
rect 325805 587866 326125 587898
rect 346874 588454 347194 588486
rect 346874 588218 346916 588454
rect 347152 588218 347194 588454
rect 346874 588134 347194 588218
rect 346874 587898 346916 588134
rect 347152 587898 347194 588134
rect 346874 587866 347194 587898
rect 352805 588454 353125 588486
rect 352805 588218 352847 588454
rect 353083 588218 353125 588454
rect 352805 588134 353125 588218
rect 352805 587898 352847 588134
rect 353083 587898 353125 588134
rect 352805 587866 353125 587898
rect 373874 588454 374194 588486
rect 373874 588218 373916 588454
rect 374152 588218 374194 588454
rect 373874 588134 374194 588218
rect 373874 587898 373916 588134
rect 374152 587898 374194 588134
rect 373874 587866 374194 587898
rect 379805 588454 380125 588486
rect 379805 588218 379847 588454
rect 380083 588218 380125 588454
rect 379805 588134 380125 588218
rect 379805 587898 379847 588134
rect 380083 587898 380125 588134
rect 379805 587866 380125 587898
rect 400874 588454 401194 588486
rect 400874 588218 400916 588454
rect 401152 588218 401194 588454
rect 400874 588134 401194 588218
rect 400874 587898 400916 588134
rect 401152 587898 401194 588134
rect 400874 587866 401194 587898
rect 406805 588454 407125 588486
rect 406805 588218 406847 588454
rect 407083 588218 407125 588454
rect 406805 588134 407125 588218
rect 406805 587898 406847 588134
rect 407083 587898 407125 588134
rect 406805 587866 407125 587898
rect 427874 588454 428194 588486
rect 427874 588218 427916 588454
rect 428152 588218 428194 588454
rect 427874 588134 428194 588218
rect 427874 587898 427916 588134
rect 428152 587898 428194 588134
rect 427874 587866 428194 587898
rect 433805 588454 434125 588486
rect 433805 588218 433847 588454
rect 434083 588218 434125 588454
rect 433805 588134 434125 588218
rect 433805 587898 433847 588134
rect 434083 587898 434125 588134
rect 433805 587866 434125 587898
rect 454874 588454 455194 588486
rect 454874 588218 454916 588454
rect 455152 588218 455194 588454
rect 454874 588134 455194 588218
rect 454874 587898 454916 588134
rect 455152 587898 455194 588134
rect 454874 587866 455194 587898
rect 460805 588454 461125 588486
rect 460805 588218 460847 588454
rect 461083 588218 461125 588454
rect 460805 588134 461125 588218
rect 460805 587898 460847 588134
rect 461083 587898 461125 588134
rect 460805 587866 461125 587898
rect 481874 588454 482194 588486
rect 481874 588218 481916 588454
rect 482152 588218 482194 588454
rect 481874 588134 482194 588218
rect 481874 587898 481916 588134
rect 482152 587898 482194 588134
rect 481874 587866 482194 587898
rect 487805 588454 488125 588486
rect 487805 588218 487847 588454
rect 488083 588218 488125 588454
rect 487805 588134 488125 588218
rect 487805 587898 487847 588134
rect 488083 587898 488125 588134
rect 487805 587866 488125 587898
rect 508874 588454 509194 588486
rect 508874 588218 508916 588454
rect 509152 588218 509194 588454
rect 508874 588134 509194 588218
rect 508874 587898 508916 588134
rect 509152 587898 509194 588134
rect 508874 587866 509194 587898
rect 514805 588454 515125 588486
rect 514805 588218 514847 588454
rect 515083 588218 515125 588454
rect 514805 588134 515125 588218
rect 514805 587898 514847 588134
rect 515083 587898 515125 588134
rect 514805 587866 515125 587898
rect 535874 588454 536194 588486
rect 535874 588218 535916 588454
rect 536152 588218 536194 588454
rect 535874 588134 536194 588218
rect 535874 587898 535916 588134
rect 536152 587898 536194 588134
rect 535874 587866 536194 587898
rect 541805 588454 542125 588486
rect 541805 588218 541847 588454
rect 542083 588218 542125 588454
rect 541805 588134 542125 588218
rect 541805 587898 541847 588134
rect 542083 587898 542125 588134
rect 541805 587866 542125 587898
rect 19794 579454 20414 581000
rect 19794 579218 19826 579454
rect 20062 579218 20146 579454
rect 20382 579218 20414 579454
rect 19794 579134 20414 579218
rect 19794 578898 19826 579134
rect 20062 578898 20146 579134
rect 20382 578898 20414 579134
rect 19794 578000 20414 578898
rect 28794 580394 29414 581000
rect 28794 580158 28826 580394
rect 29062 580158 29146 580394
rect 29382 580158 29414 580394
rect 28794 580074 29414 580158
rect 28794 579838 28826 580074
rect 29062 579838 29146 580074
rect 29382 579838 29414 580074
rect 28794 578000 29414 579838
rect 37794 579454 38414 581000
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 578000 38414 578898
rect 46794 580394 47414 581000
rect 46794 580158 46826 580394
rect 47062 580158 47146 580394
rect 47382 580158 47414 580394
rect 46794 580074 47414 580158
rect 46794 579838 46826 580074
rect 47062 579838 47146 580074
rect 47382 579838 47414 580074
rect 46794 578000 47414 579838
rect 55794 579454 56414 581000
rect 55794 579218 55826 579454
rect 56062 579218 56146 579454
rect 56382 579218 56414 579454
rect 55794 579134 56414 579218
rect 55794 578898 55826 579134
rect 56062 578898 56146 579134
rect 56382 578898 56414 579134
rect 55794 578000 56414 578898
rect 64794 580394 65414 581000
rect 64794 580158 64826 580394
rect 65062 580158 65146 580394
rect 65382 580158 65414 580394
rect 64794 580074 65414 580158
rect 64794 579838 64826 580074
rect 65062 579838 65146 580074
rect 65382 579838 65414 580074
rect 64794 578000 65414 579838
rect 73794 579454 74414 581000
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 578000 74414 578898
rect 82794 580394 83414 581000
rect 82794 580158 82826 580394
rect 83062 580158 83146 580394
rect 83382 580158 83414 580394
rect 82794 580074 83414 580158
rect 82794 579838 82826 580074
rect 83062 579838 83146 580074
rect 83382 579838 83414 580074
rect 82794 578000 83414 579838
rect 91794 579454 92414 581000
rect 91794 579218 91826 579454
rect 92062 579218 92146 579454
rect 92382 579218 92414 579454
rect 91794 579134 92414 579218
rect 91794 578898 91826 579134
rect 92062 578898 92146 579134
rect 92382 578898 92414 579134
rect 91794 578000 92414 578898
rect 100794 580394 101414 581000
rect 100794 580158 100826 580394
rect 101062 580158 101146 580394
rect 101382 580158 101414 580394
rect 100794 580074 101414 580158
rect 100794 579838 100826 580074
rect 101062 579838 101146 580074
rect 101382 579838 101414 580074
rect 100794 578000 101414 579838
rect 109794 579454 110414 581000
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 578000 110414 578898
rect 118794 580394 119414 581000
rect 118794 580158 118826 580394
rect 119062 580158 119146 580394
rect 119382 580158 119414 580394
rect 118794 580074 119414 580158
rect 118794 579838 118826 580074
rect 119062 579838 119146 580074
rect 119382 579838 119414 580074
rect 118794 578000 119414 579838
rect 127794 579454 128414 581000
rect 127794 579218 127826 579454
rect 128062 579218 128146 579454
rect 128382 579218 128414 579454
rect 127794 579134 128414 579218
rect 127794 578898 127826 579134
rect 128062 578898 128146 579134
rect 128382 578898 128414 579134
rect 127794 578000 128414 578898
rect 136794 580394 137414 581000
rect 136794 580158 136826 580394
rect 137062 580158 137146 580394
rect 137382 580158 137414 580394
rect 136794 580074 137414 580158
rect 136794 579838 136826 580074
rect 137062 579838 137146 580074
rect 137382 579838 137414 580074
rect 136794 578000 137414 579838
rect 145794 579454 146414 581000
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 578000 146414 578898
rect 154794 580394 155414 581000
rect 154794 580158 154826 580394
rect 155062 580158 155146 580394
rect 155382 580158 155414 580394
rect 154794 580074 155414 580158
rect 154794 579838 154826 580074
rect 155062 579838 155146 580074
rect 155382 579838 155414 580074
rect 154794 578000 155414 579838
rect 163794 579454 164414 581000
rect 163794 579218 163826 579454
rect 164062 579218 164146 579454
rect 164382 579218 164414 579454
rect 163794 579134 164414 579218
rect 163794 578898 163826 579134
rect 164062 578898 164146 579134
rect 164382 578898 164414 579134
rect 163794 578000 164414 578898
rect 172794 580394 173414 581000
rect 172794 580158 172826 580394
rect 173062 580158 173146 580394
rect 173382 580158 173414 580394
rect 172794 580074 173414 580158
rect 172794 579838 172826 580074
rect 173062 579838 173146 580074
rect 173382 579838 173414 580074
rect 172794 578000 173414 579838
rect 181794 579454 182414 581000
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 578000 182414 578898
rect 190794 580394 191414 581000
rect 190794 580158 190826 580394
rect 191062 580158 191146 580394
rect 191382 580158 191414 580394
rect 190794 580074 191414 580158
rect 190794 579838 190826 580074
rect 191062 579838 191146 580074
rect 191382 579838 191414 580074
rect 190794 578000 191414 579838
rect 199794 579454 200414 581000
rect 199794 579218 199826 579454
rect 200062 579218 200146 579454
rect 200382 579218 200414 579454
rect 199794 579134 200414 579218
rect 199794 578898 199826 579134
rect 200062 578898 200146 579134
rect 200382 578898 200414 579134
rect 199794 578000 200414 578898
rect 208794 580394 209414 581000
rect 208794 580158 208826 580394
rect 209062 580158 209146 580394
rect 209382 580158 209414 580394
rect 208794 580074 209414 580158
rect 208794 579838 208826 580074
rect 209062 579838 209146 580074
rect 209382 579838 209414 580074
rect 208794 578000 209414 579838
rect 217794 579454 218414 581000
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 578000 218414 578898
rect 226794 580394 227414 581000
rect 226794 580158 226826 580394
rect 227062 580158 227146 580394
rect 227382 580158 227414 580394
rect 226794 580074 227414 580158
rect 226794 579838 226826 580074
rect 227062 579838 227146 580074
rect 227382 579838 227414 580074
rect 226794 578000 227414 579838
rect 235794 579454 236414 581000
rect 235794 579218 235826 579454
rect 236062 579218 236146 579454
rect 236382 579218 236414 579454
rect 235794 579134 236414 579218
rect 235794 578898 235826 579134
rect 236062 578898 236146 579134
rect 236382 578898 236414 579134
rect 235794 578000 236414 578898
rect 244794 580394 245414 581000
rect 244794 580158 244826 580394
rect 245062 580158 245146 580394
rect 245382 580158 245414 580394
rect 244794 580074 245414 580158
rect 244794 579838 244826 580074
rect 245062 579838 245146 580074
rect 245382 579838 245414 580074
rect 244794 578000 245414 579838
rect 253794 579454 254414 581000
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 578000 254414 578898
rect 262794 580394 263414 581000
rect 262794 580158 262826 580394
rect 263062 580158 263146 580394
rect 263382 580158 263414 580394
rect 262794 580074 263414 580158
rect 262794 579838 262826 580074
rect 263062 579838 263146 580074
rect 263382 579838 263414 580074
rect 262794 578000 263414 579838
rect 271794 579454 272414 581000
rect 271794 579218 271826 579454
rect 272062 579218 272146 579454
rect 272382 579218 272414 579454
rect 271794 579134 272414 579218
rect 271794 578898 271826 579134
rect 272062 578898 272146 579134
rect 272382 578898 272414 579134
rect 271794 578000 272414 578898
rect 280794 580394 281414 581000
rect 280794 580158 280826 580394
rect 281062 580158 281146 580394
rect 281382 580158 281414 580394
rect 280794 580074 281414 580158
rect 280794 579838 280826 580074
rect 281062 579838 281146 580074
rect 281382 579838 281414 580074
rect 280794 578000 281414 579838
rect 289794 579454 290414 581000
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 578000 290414 578898
rect 298794 580394 299414 581000
rect 298794 580158 298826 580394
rect 299062 580158 299146 580394
rect 299382 580158 299414 580394
rect 298794 580074 299414 580158
rect 298794 579838 298826 580074
rect 299062 579838 299146 580074
rect 299382 579838 299414 580074
rect 298794 578000 299414 579838
rect 307794 579454 308414 581000
rect 307794 579218 307826 579454
rect 308062 579218 308146 579454
rect 308382 579218 308414 579454
rect 307794 579134 308414 579218
rect 307794 578898 307826 579134
rect 308062 578898 308146 579134
rect 308382 578898 308414 579134
rect 307794 578000 308414 578898
rect 316794 580394 317414 581000
rect 316794 580158 316826 580394
rect 317062 580158 317146 580394
rect 317382 580158 317414 580394
rect 316794 580074 317414 580158
rect 316794 579838 316826 580074
rect 317062 579838 317146 580074
rect 317382 579838 317414 580074
rect 316794 578000 317414 579838
rect 325794 579454 326414 581000
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 578000 326414 578898
rect 334794 580394 335414 581000
rect 334794 580158 334826 580394
rect 335062 580158 335146 580394
rect 335382 580158 335414 580394
rect 334794 580074 335414 580158
rect 334794 579838 334826 580074
rect 335062 579838 335146 580074
rect 335382 579838 335414 580074
rect 334794 578000 335414 579838
rect 343794 579454 344414 581000
rect 343794 579218 343826 579454
rect 344062 579218 344146 579454
rect 344382 579218 344414 579454
rect 343794 579134 344414 579218
rect 343794 578898 343826 579134
rect 344062 578898 344146 579134
rect 344382 578898 344414 579134
rect 343794 578000 344414 578898
rect 352794 580394 353414 581000
rect 352794 580158 352826 580394
rect 353062 580158 353146 580394
rect 353382 580158 353414 580394
rect 352794 580074 353414 580158
rect 352794 579838 352826 580074
rect 353062 579838 353146 580074
rect 353382 579838 353414 580074
rect 352794 578000 353414 579838
rect 361794 579454 362414 581000
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 578000 362414 578898
rect 370794 580394 371414 581000
rect 370794 580158 370826 580394
rect 371062 580158 371146 580394
rect 371382 580158 371414 580394
rect 370794 580074 371414 580158
rect 370794 579838 370826 580074
rect 371062 579838 371146 580074
rect 371382 579838 371414 580074
rect 370794 578000 371414 579838
rect 379794 579454 380414 581000
rect 379794 579218 379826 579454
rect 380062 579218 380146 579454
rect 380382 579218 380414 579454
rect 379794 579134 380414 579218
rect 379794 578898 379826 579134
rect 380062 578898 380146 579134
rect 380382 578898 380414 579134
rect 379794 578000 380414 578898
rect 388794 580394 389414 581000
rect 388794 580158 388826 580394
rect 389062 580158 389146 580394
rect 389382 580158 389414 580394
rect 388794 580074 389414 580158
rect 388794 579838 388826 580074
rect 389062 579838 389146 580074
rect 389382 579838 389414 580074
rect 388794 578000 389414 579838
rect 397794 579454 398414 581000
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 578000 398414 578898
rect 406794 580394 407414 581000
rect 406794 580158 406826 580394
rect 407062 580158 407146 580394
rect 407382 580158 407414 580394
rect 406794 580074 407414 580158
rect 406794 579838 406826 580074
rect 407062 579838 407146 580074
rect 407382 579838 407414 580074
rect 406794 578000 407414 579838
rect 415794 579454 416414 581000
rect 415794 579218 415826 579454
rect 416062 579218 416146 579454
rect 416382 579218 416414 579454
rect 415794 579134 416414 579218
rect 415794 578898 415826 579134
rect 416062 578898 416146 579134
rect 416382 578898 416414 579134
rect 415794 578000 416414 578898
rect 424794 580394 425414 581000
rect 424794 580158 424826 580394
rect 425062 580158 425146 580394
rect 425382 580158 425414 580394
rect 424794 580074 425414 580158
rect 424794 579838 424826 580074
rect 425062 579838 425146 580074
rect 425382 579838 425414 580074
rect 424794 578000 425414 579838
rect 433794 579454 434414 581000
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 578000 434414 578898
rect 442794 580394 443414 581000
rect 442794 580158 442826 580394
rect 443062 580158 443146 580394
rect 443382 580158 443414 580394
rect 442794 580074 443414 580158
rect 442794 579838 442826 580074
rect 443062 579838 443146 580074
rect 443382 579838 443414 580074
rect 442794 578000 443414 579838
rect 451794 579454 452414 581000
rect 451794 579218 451826 579454
rect 452062 579218 452146 579454
rect 452382 579218 452414 579454
rect 451794 579134 452414 579218
rect 451794 578898 451826 579134
rect 452062 578898 452146 579134
rect 452382 578898 452414 579134
rect 451794 578000 452414 578898
rect 460794 580394 461414 581000
rect 460794 580158 460826 580394
rect 461062 580158 461146 580394
rect 461382 580158 461414 580394
rect 460794 580074 461414 580158
rect 460794 579838 460826 580074
rect 461062 579838 461146 580074
rect 461382 579838 461414 580074
rect 460794 578000 461414 579838
rect 469794 579454 470414 581000
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 578000 470414 578898
rect 478794 580394 479414 581000
rect 478794 580158 478826 580394
rect 479062 580158 479146 580394
rect 479382 580158 479414 580394
rect 478794 580074 479414 580158
rect 478794 579838 478826 580074
rect 479062 579838 479146 580074
rect 479382 579838 479414 580074
rect 478794 578000 479414 579838
rect 487794 579454 488414 581000
rect 487794 579218 487826 579454
rect 488062 579218 488146 579454
rect 488382 579218 488414 579454
rect 487794 579134 488414 579218
rect 487794 578898 487826 579134
rect 488062 578898 488146 579134
rect 488382 578898 488414 579134
rect 487794 578000 488414 578898
rect 496794 580394 497414 581000
rect 496794 580158 496826 580394
rect 497062 580158 497146 580394
rect 497382 580158 497414 580394
rect 496794 580074 497414 580158
rect 496794 579838 496826 580074
rect 497062 579838 497146 580074
rect 497382 579838 497414 580074
rect 496794 578000 497414 579838
rect 505794 579454 506414 581000
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 578000 506414 578898
rect 514794 580394 515414 581000
rect 514794 580158 514826 580394
rect 515062 580158 515146 580394
rect 515382 580158 515414 580394
rect 514794 580074 515414 580158
rect 514794 579838 514826 580074
rect 515062 579838 515146 580074
rect 515382 579838 515414 580074
rect 514794 578000 515414 579838
rect 523794 579454 524414 581000
rect 523794 579218 523826 579454
rect 524062 579218 524146 579454
rect 524382 579218 524414 579454
rect 523794 579134 524414 579218
rect 523794 578898 523826 579134
rect 524062 578898 524146 579134
rect 524382 578898 524414 579134
rect 523794 578000 524414 578898
rect 532794 580394 533414 581000
rect 532794 580158 532826 580394
rect 533062 580158 533146 580394
rect 533382 580158 533414 580394
rect 532794 580074 533414 580158
rect 532794 579838 532826 580074
rect 533062 579838 533146 580074
rect 533382 579838 533414 580074
rect 532794 578000 533414 579838
rect 541794 579454 542414 581000
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 578000 542414 578898
rect 550794 580394 551414 581000
rect 550794 580158 550826 580394
rect 551062 580158 551146 580394
rect 551382 580158 551414 580394
rect 550794 580074 551414 580158
rect 550794 579838 550826 580074
rect 551062 579838 551146 580074
rect 551382 579838 551414 580074
rect 550794 578000 551414 579838
rect 559794 579454 560414 596898
rect 559794 579218 559826 579454
rect 560062 579218 560146 579454
rect 560382 579218 560414 579454
rect 559794 579134 560414 579218
rect 559794 578898 559826 579134
rect 560062 578898 560146 579134
rect 560382 578898 560414 579134
rect 10794 570218 10826 570454
rect 11062 570218 11146 570454
rect 11382 570218 11414 570454
rect 10794 570134 11414 570218
rect 10794 569898 10826 570134
rect 11062 569898 11146 570134
rect 11382 569898 11414 570134
rect 10794 552454 11414 569898
rect 22874 570454 23194 570486
rect 22874 570218 22916 570454
rect 23152 570218 23194 570454
rect 22874 570134 23194 570218
rect 22874 569898 22916 570134
rect 23152 569898 23194 570134
rect 22874 569866 23194 569898
rect 28805 570454 29125 570486
rect 28805 570218 28847 570454
rect 29083 570218 29125 570454
rect 28805 570134 29125 570218
rect 28805 569898 28847 570134
rect 29083 569898 29125 570134
rect 28805 569866 29125 569898
rect 49874 570454 50194 570486
rect 49874 570218 49916 570454
rect 50152 570218 50194 570454
rect 49874 570134 50194 570218
rect 49874 569898 49916 570134
rect 50152 569898 50194 570134
rect 49874 569866 50194 569898
rect 55805 570454 56125 570486
rect 55805 570218 55847 570454
rect 56083 570218 56125 570454
rect 55805 570134 56125 570218
rect 55805 569898 55847 570134
rect 56083 569898 56125 570134
rect 55805 569866 56125 569898
rect 76874 570454 77194 570486
rect 76874 570218 76916 570454
rect 77152 570218 77194 570454
rect 76874 570134 77194 570218
rect 76874 569898 76916 570134
rect 77152 569898 77194 570134
rect 76874 569866 77194 569898
rect 82805 570454 83125 570486
rect 82805 570218 82847 570454
rect 83083 570218 83125 570454
rect 82805 570134 83125 570218
rect 82805 569898 82847 570134
rect 83083 569898 83125 570134
rect 82805 569866 83125 569898
rect 103874 570454 104194 570486
rect 103874 570218 103916 570454
rect 104152 570218 104194 570454
rect 103874 570134 104194 570218
rect 103874 569898 103916 570134
rect 104152 569898 104194 570134
rect 103874 569866 104194 569898
rect 109805 570454 110125 570486
rect 109805 570218 109847 570454
rect 110083 570218 110125 570454
rect 109805 570134 110125 570218
rect 109805 569898 109847 570134
rect 110083 569898 110125 570134
rect 109805 569866 110125 569898
rect 130874 570454 131194 570486
rect 130874 570218 130916 570454
rect 131152 570218 131194 570454
rect 130874 570134 131194 570218
rect 130874 569898 130916 570134
rect 131152 569898 131194 570134
rect 130874 569866 131194 569898
rect 136805 570454 137125 570486
rect 136805 570218 136847 570454
rect 137083 570218 137125 570454
rect 136805 570134 137125 570218
rect 136805 569898 136847 570134
rect 137083 569898 137125 570134
rect 136805 569866 137125 569898
rect 157874 570454 158194 570486
rect 157874 570218 157916 570454
rect 158152 570218 158194 570454
rect 157874 570134 158194 570218
rect 157874 569898 157916 570134
rect 158152 569898 158194 570134
rect 157874 569866 158194 569898
rect 163805 570454 164125 570486
rect 163805 570218 163847 570454
rect 164083 570218 164125 570454
rect 163805 570134 164125 570218
rect 163805 569898 163847 570134
rect 164083 569898 164125 570134
rect 163805 569866 164125 569898
rect 184874 570454 185194 570486
rect 184874 570218 184916 570454
rect 185152 570218 185194 570454
rect 184874 570134 185194 570218
rect 184874 569898 184916 570134
rect 185152 569898 185194 570134
rect 184874 569866 185194 569898
rect 190805 570454 191125 570486
rect 190805 570218 190847 570454
rect 191083 570218 191125 570454
rect 190805 570134 191125 570218
rect 190805 569898 190847 570134
rect 191083 569898 191125 570134
rect 190805 569866 191125 569898
rect 211874 570454 212194 570486
rect 211874 570218 211916 570454
rect 212152 570218 212194 570454
rect 211874 570134 212194 570218
rect 211874 569898 211916 570134
rect 212152 569898 212194 570134
rect 211874 569866 212194 569898
rect 217805 570454 218125 570486
rect 217805 570218 217847 570454
rect 218083 570218 218125 570454
rect 217805 570134 218125 570218
rect 217805 569898 217847 570134
rect 218083 569898 218125 570134
rect 217805 569866 218125 569898
rect 238874 570454 239194 570486
rect 238874 570218 238916 570454
rect 239152 570218 239194 570454
rect 238874 570134 239194 570218
rect 238874 569898 238916 570134
rect 239152 569898 239194 570134
rect 238874 569866 239194 569898
rect 244805 570454 245125 570486
rect 244805 570218 244847 570454
rect 245083 570218 245125 570454
rect 244805 570134 245125 570218
rect 244805 569898 244847 570134
rect 245083 569898 245125 570134
rect 244805 569866 245125 569898
rect 265874 570454 266194 570486
rect 265874 570218 265916 570454
rect 266152 570218 266194 570454
rect 265874 570134 266194 570218
rect 265874 569898 265916 570134
rect 266152 569898 266194 570134
rect 265874 569866 266194 569898
rect 271805 570454 272125 570486
rect 271805 570218 271847 570454
rect 272083 570218 272125 570454
rect 271805 570134 272125 570218
rect 271805 569898 271847 570134
rect 272083 569898 272125 570134
rect 271805 569866 272125 569898
rect 292874 570454 293194 570486
rect 292874 570218 292916 570454
rect 293152 570218 293194 570454
rect 292874 570134 293194 570218
rect 292874 569898 292916 570134
rect 293152 569898 293194 570134
rect 292874 569866 293194 569898
rect 298805 570454 299125 570486
rect 298805 570218 298847 570454
rect 299083 570218 299125 570454
rect 298805 570134 299125 570218
rect 298805 569898 298847 570134
rect 299083 569898 299125 570134
rect 298805 569866 299125 569898
rect 319874 570454 320194 570486
rect 319874 570218 319916 570454
rect 320152 570218 320194 570454
rect 319874 570134 320194 570218
rect 319874 569898 319916 570134
rect 320152 569898 320194 570134
rect 319874 569866 320194 569898
rect 325805 570454 326125 570486
rect 325805 570218 325847 570454
rect 326083 570218 326125 570454
rect 325805 570134 326125 570218
rect 325805 569898 325847 570134
rect 326083 569898 326125 570134
rect 325805 569866 326125 569898
rect 346874 570454 347194 570486
rect 346874 570218 346916 570454
rect 347152 570218 347194 570454
rect 346874 570134 347194 570218
rect 346874 569898 346916 570134
rect 347152 569898 347194 570134
rect 346874 569866 347194 569898
rect 352805 570454 353125 570486
rect 352805 570218 352847 570454
rect 353083 570218 353125 570454
rect 352805 570134 353125 570218
rect 352805 569898 352847 570134
rect 353083 569898 353125 570134
rect 352805 569866 353125 569898
rect 373874 570454 374194 570486
rect 373874 570218 373916 570454
rect 374152 570218 374194 570454
rect 373874 570134 374194 570218
rect 373874 569898 373916 570134
rect 374152 569898 374194 570134
rect 373874 569866 374194 569898
rect 379805 570454 380125 570486
rect 379805 570218 379847 570454
rect 380083 570218 380125 570454
rect 379805 570134 380125 570218
rect 379805 569898 379847 570134
rect 380083 569898 380125 570134
rect 379805 569866 380125 569898
rect 400874 570454 401194 570486
rect 400874 570218 400916 570454
rect 401152 570218 401194 570454
rect 400874 570134 401194 570218
rect 400874 569898 400916 570134
rect 401152 569898 401194 570134
rect 400874 569866 401194 569898
rect 406805 570454 407125 570486
rect 406805 570218 406847 570454
rect 407083 570218 407125 570454
rect 406805 570134 407125 570218
rect 406805 569898 406847 570134
rect 407083 569898 407125 570134
rect 406805 569866 407125 569898
rect 427874 570454 428194 570486
rect 427874 570218 427916 570454
rect 428152 570218 428194 570454
rect 427874 570134 428194 570218
rect 427874 569898 427916 570134
rect 428152 569898 428194 570134
rect 427874 569866 428194 569898
rect 433805 570454 434125 570486
rect 433805 570218 433847 570454
rect 434083 570218 434125 570454
rect 433805 570134 434125 570218
rect 433805 569898 433847 570134
rect 434083 569898 434125 570134
rect 433805 569866 434125 569898
rect 454874 570454 455194 570486
rect 454874 570218 454916 570454
rect 455152 570218 455194 570454
rect 454874 570134 455194 570218
rect 454874 569898 454916 570134
rect 455152 569898 455194 570134
rect 454874 569866 455194 569898
rect 460805 570454 461125 570486
rect 460805 570218 460847 570454
rect 461083 570218 461125 570454
rect 460805 570134 461125 570218
rect 460805 569898 460847 570134
rect 461083 569898 461125 570134
rect 460805 569866 461125 569898
rect 481874 570454 482194 570486
rect 481874 570218 481916 570454
rect 482152 570218 482194 570454
rect 481874 570134 482194 570218
rect 481874 569898 481916 570134
rect 482152 569898 482194 570134
rect 481874 569866 482194 569898
rect 487805 570454 488125 570486
rect 487805 570218 487847 570454
rect 488083 570218 488125 570454
rect 487805 570134 488125 570218
rect 487805 569898 487847 570134
rect 488083 569898 488125 570134
rect 487805 569866 488125 569898
rect 508874 570454 509194 570486
rect 508874 570218 508916 570454
rect 509152 570218 509194 570454
rect 508874 570134 509194 570218
rect 508874 569898 508916 570134
rect 509152 569898 509194 570134
rect 508874 569866 509194 569898
rect 514805 570454 515125 570486
rect 514805 570218 514847 570454
rect 515083 570218 515125 570454
rect 514805 570134 515125 570218
rect 514805 569898 514847 570134
rect 515083 569898 515125 570134
rect 514805 569866 515125 569898
rect 535874 570454 536194 570486
rect 535874 570218 535916 570454
rect 536152 570218 536194 570454
rect 535874 570134 536194 570218
rect 535874 569898 535916 570134
rect 536152 569898 536194 570134
rect 535874 569866 536194 569898
rect 541805 570454 542125 570486
rect 541805 570218 541847 570454
rect 542083 570218 542125 570454
rect 541805 570134 542125 570218
rect 541805 569898 541847 570134
rect 542083 569898 542125 570134
rect 541805 569866 542125 569898
rect 19910 561454 20230 561486
rect 19910 561218 19952 561454
rect 20188 561218 20230 561454
rect 19910 561134 20230 561218
rect 19910 560898 19952 561134
rect 20188 560898 20230 561134
rect 19910 560866 20230 560898
rect 25840 561454 26160 561486
rect 25840 561218 25882 561454
rect 26118 561218 26160 561454
rect 25840 561134 26160 561218
rect 25840 560898 25882 561134
rect 26118 560898 26160 561134
rect 25840 560866 26160 560898
rect 31771 561454 32091 561486
rect 31771 561218 31813 561454
rect 32049 561218 32091 561454
rect 31771 561134 32091 561218
rect 31771 560898 31813 561134
rect 32049 560898 32091 561134
rect 31771 560866 32091 560898
rect 46910 561454 47230 561486
rect 46910 561218 46952 561454
rect 47188 561218 47230 561454
rect 46910 561134 47230 561218
rect 46910 560898 46952 561134
rect 47188 560898 47230 561134
rect 46910 560866 47230 560898
rect 52840 561454 53160 561486
rect 52840 561218 52882 561454
rect 53118 561218 53160 561454
rect 52840 561134 53160 561218
rect 52840 560898 52882 561134
rect 53118 560898 53160 561134
rect 52840 560866 53160 560898
rect 58771 561454 59091 561486
rect 58771 561218 58813 561454
rect 59049 561218 59091 561454
rect 58771 561134 59091 561218
rect 58771 560898 58813 561134
rect 59049 560898 59091 561134
rect 58771 560866 59091 560898
rect 73910 561454 74230 561486
rect 73910 561218 73952 561454
rect 74188 561218 74230 561454
rect 73910 561134 74230 561218
rect 73910 560898 73952 561134
rect 74188 560898 74230 561134
rect 73910 560866 74230 560898
rect 79840 561454 80160 561486
rect 79840 561218 79882 561454
rect 80118 561218 80160 561454
rect 79840 561134 80160 561218
rect 79840 560898 79882 561134
rect 80118 560898 80160 561134
rect 79840 560866 80160 560898
rect 85771 561454 86091 561486
rect 85771 561218 85813 561454
rect 86049 561218 86091 561454
rect 85771 561134 86091 561218
rect 85771 560898 85813 561134
rect 86049 560898 86091 561134
rect 85771 560866 86091 560898
rect 100910 561454 101230 561486
rect 100910 561218 100952 561454
rect 101188 561218 101230 561454
rect 100910 561134 101230 561218
rect 100910 560898 100952 561134
rect 101188 560898 101230 561134
rect 100910 560866 101230 560898
rect 106840 561454 107160 561486
rect 106840 561218 106882 561454
rect 107118 561218 107160 561454
rect 106840 561134 107160 561218
rect 106840 560898 106882 561134
rect 107118 560898 107160 561134
rect 106840 560866 107160 560898
rect 112771 561454 113091 561486
rect 112771 561218 112813 561454
rect 113049 561218 113091 561454
rect 112771 561134 113091 561218
rect 112771 560898 112813 561134
rect 113049 560898 113091 561134
rect 112771 560866 113091 560898
rect 127910 561454 128230 561486
rect 127910 561218 127952 561454
rect 128188 561218 128230 561454
rect 127910 561134 128230 561218
rect 127910 560898 127952 561134
rect 128188 560898 128230 561134
rect 127910 560866 128230 560898
rect 133840 561454 134160 561486
rect 133840 561218 133882 561454
rect 134118 561218 134160 561454
rect 133840 561134 134160 561218
rect 133840 560898 133882 561134
rect 134118 560898 134160 561134
rect 133840 560866 134160 560898
rect 139771 561454 140091 561486
rect 139771 561218 139813 561454
rect 140049 561218 140091 561454
rect 139771 561134 140091 561218
rect 139771 560898 139813 561134
rect 140049 560898 140091 561134
rect 139771 560866 140091 560898
rect 154910 561454 155230 561486
rect 154910 561218 154952 561454
rect 155188 561218 155230 561454
rect 154910 561134 155230 561218
rect 154910 560898 154952 561134
rect 155188 560898 155230 561134
rect 154910 560866 155230 560898
rect 160840 561454 161160 561486
rect 160840 561218 160882 561454
rect 161118 561218 161160 561454
rect 160840 561134 161160 561218
rect 160840 560898 160882 561134
rect 161118 560898 161160 561134
rect 160840 560866 161160 560898
rect 166771 561454 167091 561486
rect 166771 561218 166813 561454
rect 167049 561218 167091 561454
rect 166771 561134 167091 561218
rect 166771 560898 166813 561134
rect 167049 560898 167091 561134
rect 166771 560866 167091 560898
rect 181910 561454 182230 561486
rect 181910 561218 181952 561454
rect 182188 561218 182230 561454
rect 181910 561134 182230 561218
rect 181910 560898 181952 561134
rect 182188 560898 182230 561134
rect 181910 560866 182230 560898
rect 187840 561454 188160 561486
rect 187840 561218 187882 561454
rect 188118 561218 188160 561454
rect 187840 561134 188160 561218
rect 187840 560898 187882 561134
rect 188118 560898 188160 561134
rect 187840 560866 188160 560898
rect 193771 561454 194091 561486
rect 193771 561218 193813 561454
rect 194049 561218 194091 561454
rect 193771 561134 194091 561218
rect 193771 560898 193813 561134
rect 194049 560898 194091 561134
rect 193771 560866 194091 560898
rect 208910 561454 209230 561486
rect 208910 561218 208952 561454
rect 209188 561218 209230 561454
rect 208910 561134 209230 561218
rect 208910 560898 208952 561134
rect 209188 560898 209230 561134
rect 208910 560866 209230 560898
rect 214840 561454 215160 561486
rect 214840 561218 214882 561454
rect 215118 561218 215160 561454
rect 214840 561134 215160 561218
rect 214840 560898 214882 561134
rect 215118 560898 215160 561134
rect 214840 560866 215160 560898
rect 220771 561454 221091 561486
rect 220771 561218 220813 561454
rect 221049 561218 221091 561454
rect 220771 561134 221091 561218
rect 220771 560898 220813 561134
rect 221049 560898 221091 561134
rect 220771 560866 221091 560898
rect 235910 561454 236230 561486
rect 235910 561218 235952 561454
rect 236188 561218 236230 561454
rect 235910 561134 236230 561218
rect 235910 560898 235952 561134
rect 236188 560898 236230 561134
rect 235910 560866 236230 560898
rect 241840 561454 242160 561486
rect 241840 561218 241882 561454
rect 242118 561218 242160 561454
rect 241840 561134 242160 561218
rect 241840 560898 241882 561134
rect 242118 560898 242160 561134
rect 241840 560866 242160 560898
rect 247771 561454 248091 561486
rect 247771 561218 247813 561454
rect 248049 561218 248091 561454
rect 247771 561134 248091 561218
rect 247771 560898 247813 561134
rect 248049 560898 248091 561134
rect 247771 560866 248091 560898
rect 262910 561454 263230 561486
rect 262910 561218 262952 561454
rect 263188 561218 263230 561454
rect 262910 561134 263230 561218
rect 262910 560898 262952 561134
rect 263188 560898 263230 561134
rect 262910 560866 263230 560898
rect 268840 561454 269160 561486
rect 268840 561218 268882 561454
rect 269118 561218 269160 561454
rect 268840 561134 269160 561218
rect 268840 560898 268882 561134
rect 269118 560898 269160 561134
rect 268840 560866 269160 560898
rect 274771 561454 275091 561486
rect 274771 561218 274813 561454
rect 275049 561218 275091 561454
rect 274771 561134 275091 561218
rect 274771 560898 274813 561134
rect 275049 560898 275091 561134
rect 274771 560866 275091 560898
rect 289910 561454 290230 561486
rect 289910 561218 289952 561454
rect 290188 561218 290230 561454
rect 289910 561134 290230 561218
rect 289910 560898 289952 561134
rect 290188 560898 290230 561134
rect 289910 560866 290230 560898
rect 295840 561454 296160 561486
rect 295840 561218 295882 561454
rect 296118 561218 296160 561454
rect 295840 561134 296160 561218
rect 295840 560898 295882 561134
rect 296118 560898 296160 561134
rect 295840 560866 296160 560898
rect 301771 561454 302091 561486
rect 301771 561218 301813 561454
rect 302049 561218 302091 561454
rect 301771 561134 302091 561218
rect 301771 560898 301813 561134
rect 302049 560898 302091 561134
rect 301771 560866 302091 560898
rect 316910 561454 317230 561486
rect 316910 561218 316952 561454
rect 317188 561218 317230 561454
rect 316910 561134 317230 561218
rect 316910 560898 316952 561134
rect 317188 560898 317230 561134
rect 316910 560866 317230 560898
rect 322840 561454 323160 561486
rect 322840 561218 322882 561454
rect 323118 561218 323160 561454
rect 322840 561134 323160 561218
rect 322840 560898 322882 561134
rect 323118 560898 323160 561134
rect 322840 560866 323160 560898
rect 328771 561454 329091 561486
rect 328771 561218 328813 561454
rect 329049 561218 329091 561454
rect 328771 561134 329091 561218
rect 328771 560898 328813 561134
rect 329049 560898 329091 561134
rect 328771 560866 329091 560898
rect 343910 561454 344230 561486
rect 343910 561218 343952 561454
rect 344188 561218 344230 561454
rect 343910 561134 344230 561218
rect 343910 560898 343952 561134
rect 344188 560898 344230 561134
rect 343910 560866 344230 560898
rect 349840 561454 350160 561486
rect 349840 561218 349882 561454
rect 350118 561218 350160 561454
rect 349840 561134 350160 561218
rect 349840 560898 349882 561134
rect 350118 560898 350160 561134
rect 349840 560866 350160 560898
rect 355771 561454 356091 561486
rect 355771 561218 355813 561454
rect 356049 561218 356091 561454
rect 355771 561134 356091 561218
rect 355771 560898 355813 561134
rect 356049 560898 356091 561134
rect 355771 560866 356091 560898
rect 370910 561454 371230 561486
rect 370910 561218 370952 561454
rect 371188 561218 371230 561454
rect 370910 561134 371230 561218
rect 370910 560898 370952 561134
rect 371188 560898 371230 561134
rect 370910 560866 371230 560898
rect 376840 561454 377160 561486
rect 376840 561218 376882 561454
rect 377118 561218 377160 561454
rect 376840 561134 377160 561218
rect 376840 560898 376882 561134
rect 377118 560898 377160 561134
rect 376840 560866 377160 560898
rect 382771 561454 383091 561486
rect 382771 561218 382813 561454
rect 383049 561218 383091 561454
rect 382771 561134 383091 561218
rect 382771 560898 382813 561134
rect 383049 560898 383091 561134
rect 382771 560866 383091 560898
rect 397910 561454 398230 561486
rect 397910 561218 397952 561454
rect 398188 561218 398230 561454
rect 397910 561134 398230 561218
rect 397910 560898 397952 561134
rect 398188 560898 398230 561134
rect 397910 560866 398230 560898
rect 403840 561454 404160 561486
rect 403840 561218 403882 561454
rect 404118 561218 404160 561454
rect 403840 561134 404160 561218
rect 403840 560898 403882 561134
rect 404118 560898 404160 561134
rect 403840 560866 404160 560898
rect 409771 561454 410091 561486
rect 409771 561218 409813 561454
rect 410049 561218 410091 561454
rect 409771 561134 410091 561218
rect 409771 560898 409813 561134
rect 410049 560898 410091 561134
rect 409771 560866 410091 560898
rect 424910 561454 425230 561486
rect 424910 561218 424952 561454
rect 425188 561218 425230 561454
rect 424910 561134 425230 561218
rect 424910 560898 424952 561134
rect 425188 560898 425230 561134
rect 424910 560866 425230 560898
rect 430840 561454 431160 561486
rect 430840 561218 430882 561454
rect 431118 561218 431160 561454
rect 430840 561134 431160 561218
rect 430840 560898 430882 561134
rect 431118 560898 431160 561134
rect 430840 560866 431160 560898
rect 436771 561454 437091 561486
rect 436771 561218 436813 561454
rect 437049 561218 437091 561454
rect 436771 561134 437091 561218
rect 436771 560898 436813 561134
rect 437049 560898 437091 561134
rect 436771 560866 437091 560898
rect 451910 561454 452230 561486
rect 451910 561218 451952 561454
rect 452188 561218 452230 561454
rect 451910 561134 452230 561218
rect 451910 560898 451952 561134
rect 452188 560898 452230 561134
rect 451910 560866 452230 560898
rect 457840 561454 458160 561486
rect 457840 561218 457882 561454
rect 458118 561218 458160 561454
rect 457840 561134 458160 561218
rect 457840 560898 457882 561134
rect 458118 560898 458160 561134
rect 457840 560866 458160 560898
rect 463771 561454 464091 561486
rect 463771 561218 463813 561454
rect 464049 561218 464091 561454
rect 463771 561134 464091 561218
rect 463771 560898 463813 561134
rect 464049 560898 464091 561134
rect 463771 560866 464091 560898
rect 478910 561454 479230 561486
rect 478910 561218 478952 561454
rect 479188 561218 479230 561454
rect 478910 561134 479230 561218
rect 478910 560898 478952 561134
rect 479188 560898 479230 561134
rect 478910 560866 479230 560898
rect 484840 561454 485160 561486
rect 484840 561218 484882 561454
rect 485118 561218 485160 561454
rect 484840 561134 485160 561218
rect 484840 560898 484882 561134
rect 485118 560898 485160 561134
rect 484840 560866 485160 560898
rect 490771 561454 491091 561486
rect 490771 561218 490813 561454
rect 491049 561218 491091 561454
rect 490771 561134 491091 561218
rect 490771 560898 490813 561134
rect 491049 560898 491091 561134
rect 490771 560866 491091 560898
rect 505910 561454 506230 561486
rect 505910 561218 505952 561454
rect 506188 561218 506230 561454
rect 505910 561134 506230 561218
rect 505910 560898 505952 561134
rect 506188 560898 506230 561134
rect 505910 560866 506230 560898
rect 511840 561454 512160 561486
rect 511840 561218 511882 561454
rect 512118 561218 512160 561454
rect 511840 561134 512160 561218
rect 511840 560898 511882 561134
rect 512118 560898 512160 561134
rect 511840 560866 512160 560898
rect 517771 561454 518091 561486
rect 517771 561218 517813 561454
rect 518049 561218 518091 561454
rect 517771 561134 518091 561218
rect 517771 560898 517813 561134
rect 518049 560898 518091 561134
rect 517771 560866 518091 560898
rect 532910 561454 533230 561486
rect 532910 561218 532952 561454
rect 533188 561218 533230 561454
rect 532910 561134 533230 561218
rect 532910 560898 532952 561134
rect 533188 560898 533230 561134
rect 532910 560866 533230 560898
rect 538840 561454 539160 561486
rect 538840 561218 538882 561454
rect 539118 561218 539160 561454
rect 538840 561134 539160 561218
rect 538840 560898 538882 561134
rect 539118 560898 539160 561134
rect 538840 560866 539160 560898
rect 544771 561454 545091 561486
rect 544771 561218 544813 561454
rect 545049 561218 545091 561454
rect 544771 561134 545091 561218
rect 544771 560898 544813 561134
rect 545049 560898 545091 561134
rect 544771 560866 545091 560898
rect 559794 561454 560414 578898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 534454 11414 551898
rect 19794 553394 20414 554000
rect 19794 553158 19826 553394
rect 20062 553158 20146 553394
rect 20382 553158 20414 553394
rect 19794 553074 20414 553158
rect 19794 552838 19826 553074
rect 20062 552838 20146 553074
rect 20382 552838 20414 553074
rect 19794 551000 20414 552838
rect 28794 552454 29414 554000
rect 28794 552218 28826 552454
rect 29062 552218 29146 552454
rect 29382 552218 29414 552454
rect 28794 552134 29414 552218
rect 28794 551898 28826 552134
rect 29062 551898 29146 552134
rect 29382 551898 29414 552134
rect 28794 551000 29414 551898
rect 37794 553394 38414 554000
rect 37794 553158 37826 553394
rect 38062 553158 38146 553394
rect 38382 553158 38414 553394
rect 37794 553074 38414 553158
rect 37794 552838 37826 553074
rect 38062 552838 38146 553074
rect 38382 552838 38414 553074
rect 37794 551000 38414 552838
rect 46794 552454 47414 554000
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 551000 47414 551898
rect 55794 553394 56414 554000
rect 55794 553158 55826 553394
rect 56062 553158 56146 553394
rect 56382 553158 56414 553394
rect 55794 553074 56414 553158
rect 55794 552838 55826 553074
rect 56062 552838 56146 553074
rect 56382 552838 56414 553074
rect 55794 551000 56414 552838
rect 64794 552454 65414 554000
rect 64794 552218 64826 552454
rect 65062 552218 65146 552454
rect 65382 552218 65414 552454
rect 64794 552134 65414 552218
rect 64794 551898 64826 552134
rect 65062 551898 65146 552134
rect 65382 551898 65414 552134
rect 64794 551000 65414 551898
rect 73794 553394 74414 554000
rect 73794 553158 73826 553394
rect 74062 553158 74146 553394
rect 74382 553158 74414 553394
rect 73794 553074 74414 553158
rect 73794 552838 73826 553074
rect 74062 552838 74146 553074
rect 74382 552838 74414 553074
rect 73794 551000 74414 552838
rect 82794 552454 83414 554000
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 551000 83414 551898
rect 91794 553394 92414 554000
rect 91794 553158 91826 553394
rect 92062 553158 92146 553394
rect 92382 553158 92414 553394
rect 91794 553074 92414 553158
rect 91794 552838 91826 553074
rect 92062 552838 92146 553074
rect 92382 552838 92414 553074
rect 91794 551000 92414 552838
rect 100794 552454 101414 554000
rect 100794 552218 100826 552454
rect 101062 552218 101146 552454
rect 101382 552218 101414 552454
rect 100794 552134 101414 552218
rect 100794 551898 100826 552134
rect 101062 551898 101146 552134
rect 101382 551898 101414 552134
rect 100794 551000 101414 551898
rect 109794 553394 110414 554000
rect 109794 553158 109826 553394
rect 110062 553158 110146 553394
rect 110382 553158 110414 553394
rect 109794 553074 110414 553158
rect 109794 552838 109826 553074
rect 110062 552838 110146 553074
rect 110382 552838 110414 553074
rect 109794 551000 110414 552838
rect 118794 552454 119414 554000
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 551000 119414 551898
rect 127794 553394 128414 554000
rect 127794 553158 127826 553394
rect 128062 553158 128146 553394
rect 128382 553158 128414 553394
rect 127794 553074 128414 553158
rect 127794 552838 127826 553074
rect 128062 552838 128146 553074
rect 128382 552838 128414 553074
rect 127794 551000 128414 552838
rect 136794 552454 137414 554000
rect 136794 552218 136826 552454
rect 137062 552218 137146 552454
rect 137382 552218 137414 552454
rect 136794 552134 137414 552218
rect 136794 551898 136826 552134
rect 137062 551898 137146 552134
rect 137382 551898 137414 552134
rect 136794 551000 137414 551898
rect 145794 553394 146414 554000
rect 145794 553158 145826 553394
rect 146062 553158 146146 553394
rect 146382 553158 146414 553394
rect 145794 553074 146414 553158
rect 145794 552838 145826 553074
rect 146062 552838 146146 553074
rect 146382 552838 146414 553074
rect 145794 551000 146414 552838
rect 154794 552454 155414 554000
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 551000 155414 551898
rect 163794 553394 164414 554000
rect 163794 553158 163826 553394
rect 164062 553158 164146 553394
rect 164382 553158 164414 553394
rect 163794 553074 164414 553158
rect 163794 552838 163826 553074
rect 164062 552838 164146 553074
rect 164382 552838 164414 553074
rect 163794 551000 164414 552838
rect 172794 552454 173414 554000
rect 172794 552218 172826 552454
rect 173062 552218 173146 552454
rect 173382 552218 173414 552454
rect 172794 552134 173414 552218
rect 172794 551898 172826 552134
rect 173062 551898 173146 552134
rect 173382 551898 173414 552134
rect 172794 551000 173414 551898
rect 181794 553394 182414 554000
rect 181794 553158 181826 553394
rect 182062 553158 182146 553394
rect 182382 553158 182414 553394
rect 181794 553074 182414 553158
rect 181794 552838 181826 553074
rect 182062 552838 182146 553074
rect 182382 552838 182414 553074
rect 181794 551000 182414 552838
rect 190794 552454 191414 554000
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 551000 191414 551898
rect 199794 553394 200414 554000
rect 199794 553158 199826 553394
rect 200062 553158 200146 553394
rect 200382 553158 200414 553394
rect 199794 553074 200414 553158
rect 199794 552838 199826 553074
rect 200062 552838 200146 553074
rect 200382 552838 200414 553074
rect 199794 551000 200414 552838
rect 208794 552454 209414 554000
rect 208794 552218 208826 552454
rect 209062 552218 209146 552454
rect 209382 552218 209414 552454
rect 208794 552134 209414 552218
rect 208794 551898 208826 552134
rect 209062 551898 209146 552134
rect 209382 551898 209414 552134
rect 208794 551000 209414 551898
rect 217794 553394 218414 554000
rect 217794 553158 217826 553394
rect 218062 553158 218146 553394
rect 218382 553158 218414 553394
rect 217794 553074 218414 553158
rect 217794 552838 217826 553074
rect 218062 552838 218146 553074
rect 218382 552838 218414 553074
rect 217794 551000 218414 552838
rect 226794 552454 227414 554000
rect 226794 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 227414 552454
rect 226794 552134 227414 552218
rect 226794 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 227414 552134
rect 226794 551000 227414 551898
rect 235794 553394 236414 554000
rect 235794 553158 235826 553394
rect 236062 553158 236146 553394
rect 236382 553158 236414 553394
rect 235794 553074 236414 553158
rect 235794 552838 235826 553074
rect 236062 552838 236146 553074
rect 236382 552838 236414 553074
rect 235794 551000 236414 552838
rect 244794 552454 245414 554000
rect 244794 552218 244826 552454
rect 245062 552218 245146 552454
rect 245382 552218 245414 552454
rect 244794 552134 245414 552218
rect 244794 551898 244826 552134
rect 245062 551898 245146 552134
rect 245382 551898 245414 552134
rect 244794 551000 245414 551898
rect 253794 553394 254414 554000
rect 253794 553158 253826 553394
rect 254062 553158 254146 553394
rect 254382 553158 254414 553394
rect 253794 553074 254414 553158
rect 253794 552838 253826 553074
rect 254062 552838 254146 553074
rect 254382 552838 254414 553074
rect 253794 551000 254414 552838
rect 262794 552454 263414 554000
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 551000 263414 551898
rect 271794 553394 272414 554000
rect 271794 553158 271826 553394
rect 272062 553158 272146 553394
rect 272382 553158 272414 553394
rect 271794 553074 272414 553158
rect 271794 552838 271826 553074
rect 272062 552838 272146 553074
rect 272382 552838 272414 553074
rect 271794 551000 272414 552838
rect 280794 552454 281414 554000
rect 280794 552218 280826 552454
rect 281062 552218 281146 552454
rect 281382 552218 281414 552454
rect 280794 552134 281414 552218
rect 280794 551898 280826 552134
rect 281062 551898 281146 552134
rect 281382 551898 281414 552134
rect 280794 551000 281414 551898
rect 289794 553394 290414 554000
rect 289794 553158 289826 553394
rect 290062 553158 290146 553394
rect 290382 553158 290414 553394
rect 289794 553074 290414 553158
rect 289794 552838 289826 553074
rect 290062 552838 290146 553074
rect 290382 552838 290414 553074
rect 289794 551000 290414 552838
rect 298794 552454 299414 554000
rect 298794 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 299414 552454
rect 298794 552134 299414 552218
rect 298794 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 299414 552134
rect 298794 551000 299414 551898
rect 307794 553394 308414 554000
rect 307794 553158 307826 553394
rect 308062 553158 308146 553394
rect 308382 553158 308414 553394
rect 307794 553074 308414 553158
rect 307794 552838 307826 553074
rect 308062 552838 308146 553074
rect 308382 552838 308414 553074
rect 307794 551000 308414 552838
rect 316794 552454 317414 554000
rect 316794 552218 316826 552454
rect 317062 552218 317146 552454
rect 317382 552218 317414 552454
rect 316794 552134 317414 552218
rect 316794 551898 316826 552134
rect 317062 551898 317146 552134
rect 317382 551898 317414 552134
rect 316794 551000 317414 551898
rect 325794 553394 326414 554000
rect 325794 553158 325826 553394
rect 326062 553158 326146 553394
rect 326382 553158 326414 553394
rect 325794 553074 326414 553158
rect 325794 552838 325826 553074
rect 326062 552838 326146 553074
rect 326382 552838 326414 553074
rect 325794 551000 326414 552838
rect 334794 552454 335414 554000
rect 334794 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 335414 552454
rect 334794 552134 335414 552218
rect 334794 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 335414 552134
rect 334794 551000 335414 551898
rect 343794 553394 344414 554000
rect 343794 553158 343826 553394
rect 344062 553158 344146 553394
rect 344382 553158 344414 553394
rect 343794 553074 344414 553158
rect 343794 552838 343826 553074
rect 344062 552838 344146 553074
rect 344382 552838 344414 553074
rect 343794 551000 344414 552838
rect 352794 552454 353414 554000
rect 352794 552218 352826 552454
rect 353062 552218 353146 552454
rect 353382 552218 353414 552454
rect 352794 552134 353414 552218
rect 352794 551898 352826 552134
rect 353062 551898 353146 552134
rect 353382 551898 353414 552134
rect 352794 551000 353414 551898
rect 361794 553394 362414 554000
rect 361794 553158 361826 553394
rect 362062 553158 362146 553394
rect 362382 553158 362414 553394
rect 361794 553074 362414 553158
rect 361794 552838 361826 553074
rect 362062 552838 362146 553074
rect 362382 552838 362414 553074
rect 361794 551000 362414 552838
rect 370794 552454 371414 554000
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 551000 371414 551898
rect 379794 553394 380414 554000
rect 379794 553158 379826 553394
rect 380062 553158 380146 553394
rect 380382 553158 380414 553394
rect 379794 553074 380414 553158
rect 379794 552838 379826 553074
rect 380062 552838 380146 553074
rect 380382 552838 380414 553074
rect 379794 551000 380414 552838
rect 388794 552454 389414 554000
rect 388794 552218 388826 552454
rect 389062 552218 389146 552454
rect 389382 552218 389414 552454
rect 388794 552134 389414 552218
rect 388794 551898 388826 552134
rect 389062 551898 389146 552134
rect 389382 551898 389414 552134
rect 388794 551000 389414 551898
rect 397794 553394 398414 554000
rect 397794 553158 397826 553394
rect 398062 553158 398146 553394
rect 398382 553158 398414 553394
rect 397794 553074 398414 553158
rect 397794 552838 397826 553074
rect 398062 552838 398146 553074
rect 398382 552838 398414 553074
rect 397794 551000 398414 552838
rect 406794 552454 407414 554000
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 551000 407414 551898
rect 415794 553394 416414 554000
rect 415794 553158 415826 553394
rect 416062 553158 416146 553394
rect 416382 553158 416414 553394
rect 415794 553074 416414 553158
rect 415794 552838 415826 553074
rect 416062 552838 416146 553074
rect 416382 552838 416414 553074
rect 415794 551000 416414 552838
rect 424794 552454 425414 554000
rect 424794 552218 424826 552454
rect 425062 552218 425146 552454
rect 425382 552218 425414 552454
rect 424794 552134 425414 552218
rect 424794 551898 424826 552134
rect 425062 551898 425146 552134
rect 425382 551898 425414 552134
rect 424794 551000 425414 551898
rect 433794 553394 434414 554000
rect 433794 553158 433826 553394
rect 434062 553158 434146 553394
rect 434382 553158 434414 553394
rect 433794 553074 434414 553158
rect 433794 552838 433826 553074
rect 434062 552838 434146 553074
rect 434382 552838 434414 553074
rect 433794 551000 434414 552838
rect 442794 552454 443414 554000
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 551000 443414 551898
rect 451794 553394 452414 554000
rect 451794 553158 451826 553394
rect 452062 553158 452146 553394
rect 452382 553158 452414 553394
rect 451794 553074 452414 553158
rect 451794 552838 451826 553074
rect 452062 552838 452146 553074
rect 452382 552838 452414 553074
rect 451794 551000 452414 552838
rect 460794 552454 461414 554000
rect 460794 552218 460826 552454
rect 461062 552218 461146 552454
rect 461382 552218 461414 552454
rect 460794 552134 461414 552218
rect 460794 551898 460826 552134
rect 461062 551898 461146 552134
rect 461382 551898 461414 552134
rect 460794 551000 461414 551898
rect 469794 553394 470414 554000
rect 469794 553158 469826 553394
rect 470062 553158 470146 553394
rect 470382 553158 470414 553394
rect 469794 553074 470414 553158
rect 469794 552838 469826 553074
rect 470062 552838 470146 553074
rect 470382 552838 470414 553074
rect 469794 551000 470414 552838
rect 478794 552454 479414 554000
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 551000 479414 551898
rect 487794 553394 488414 554000
rect 487794 553158 487826 553394
rect 488062 553158 488146 553394
rect 488382 553158 488414 553394
rect 487794 553074 488414 553158
rect 487794 552838 487826 553074
rect 488062 552838 488146 553074
rect 488382 552838 488414 553074
rect 487794 551000 488414 552838
rect 496794 552454 497414 554000
rect 496794 552218 496826 552454
rect 497062 552218 497146 552454
rect 497382 552218 497414 552454
rect 496794 552134 497414 552218
rect 496794 551898 496826 552134
rect 497062 551898 497146 552134
rect 497382 551898 497414 552134
rect 496794 551000 497414 551898
rect 505794 553394 506414 554000
rect 505794 553158 505826 553394
rect 506062 553158 506146 553394
rect 506382 553158 506414 553394
rect 505794 553074 506414 553158
rect 505794 552838 505826 553074
rect 506062 552838 506146 553074
rect 506382 552838 506414 553074
rect 505794 551000 506414 552838
rect 514794 552454 515414 554000
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 551000 515414 551898
rect 523794 553394 524414 554000
rect 523794 553158 523826 553394
rect 524062 553158 524146 553394
rect 524382 553158 524414 553394
rect 523794 553074 524414 553158
rect 523794 552838 523826 553074
rect 524062 552838 524146 553074
rect 524382 552838 524414 553074
rect 523794 551000 524414 552838
rect 532794 552454 533414 554000
rect 532794 552218 532826 552454
rect 533062 552218 533146 552454
rect 533382 552218 533414 552454
rect 532794 552134 533414 552218
rect 532794 551898 532826 552134
rect 533062 551898 533146 552134
rect 533382 551898 533414 552134
rect 532794 551000 533414 551898
rect 541794 553394 542414 554000
rect 541794 553158 541826 553394
rect 542062 553158 542146 553394
rect 542382 553158 542414 553394
rect 541794 553074 542414 553158
rect 541794 552838 541826 553074
rect 542062 552838 542146 553074
rect 542382 552838 542414 553074
rect 541794 551000 542414 552838
rect 550794 552454 551414 554000
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 551000 551414 551898
rect 19910 543454 20230 543486
rect 19910 543218 19952 543454
rect 20188 543218 20230 543454
rect 19910 543134 20230 543218
rect 19910 542898 19952 543134
rect 20188 542898 20230 543134
rect 19910 542866 20230 542898
rect 25840 543454 26160 543486
rect 25840 543218 25882 543454
rect 26118 543218 26160 543454
rect 25840 543134 26160 543218
rect 25840 542898 25882 543134
rect 26118 542898 26160 543134
rect 25840 542866 26160 542898
rect 31771 543454 32091 543486
rect 31771 543218 31813 543454
rect 32049 543218 32091 543454
rect 31771 543134 32091 543218
rect 31771 542898 31813 543134
rect 32049 542898 32091 543134
rect 31771 542866 32091 542898
rect 46910 543454 47230 543486
rect 46910 543218 46952 543454
rect 47188 543218 47230 543454
rect 46910 543134 47230 543218
rect 46910 542898 46952 543134
rect 47188 542898 47230 543134
rect 46910 542866 47230 542898
rect 52840 543454 53160 543486
rect 52840 543218 52882 543454
rect 53118 543218 53160 543454
rect 52840 543134 53160 543218
rect 52840 542898 52882 543134
rect 53118 542898 53160 543134
rect 52840 542866 53160 542898
rect 58771 543454 59091 543486
rect 58771 543218 58813 543454
rect 59049 543218 59091 543454
rect 58771 543134 59091 543218
rect 58771 542898 58813 543134
rect 59049 542898 59091 543134
rect 58771 542866 59091 542898
rect 73910 543454 74230 543486
rect 73910 543218 73952 543454
rect 74188 543218 74230 543454
rect 73910 543134 74230 543218
rect 73910 542898 73952 543134
rect 74188 542898 74230 543134
rect 73910 542866 74230 542898
rect 79840 543454 80160 543486
rect 79840 543218 79882 543454
rect 80118 543218 80160 543454
rect 79840 543134 80160 543218
rect 79840 542898 79882 543134
rect 80118 542898 80160 543134
rect 79840 542866 80160 542898
rect 85771 543454 86091 543486
rect 85771 543218 85813 543454
rect 86049 543218 86091 543454
rect 85771 543134 86091 543218
rect 85771 542898 85813 543134
rect 86049 542898 86091 543134
rect 85771 542866 86091 542898
rect 100910 543454 101230 543486
rect 100910 543218 100952 543454
rect 101188 543218 101230 543454
rect 100910 543134 101230 543218
rect 100910 542898 100952 543134
rect 101188 542898 101230 543134
rect 100910 542866 101230 542898
rect 106840 543454 107160 543486
rect 106840 543218 106882 543454
rect 107118 543218 107160 543454
rect 106840 543134 107160 543218
rect 106840 542898 106882 543134
rect 107118 542898 107160 543134
rect 106840 542866 107160 542898
rect 112771 543454 113091 543486
rect 112771 543218 112813 543454
rect 113049 543218 113091 543454
rect 112771 543134 113091 543218
rect 112771 542898 112813 543134
rect 113049 542898 113091 543134
rect 112771 542866 113091 542898
rect 127910 543454 128230 543486
rect 127910 543218 127952 543454
rect 128188 543218 128230 543454
rect 127910 543134 128230 543218
rect 127910 542898 127952 543134
rect 128188 542898 128230 543134
rect 127910 542866 128230 542898
rect 133840 543454 134160 543486
rect 133840 543218 133882 543454
rect 134118 543218 134160 543454
rect 133840 543134 134160 543218
rect 133840 542898 133882 543134
rect 134118 542898 134160 543134
rect 133840 542866 134160 542898
rect 139771 543454 140091 543486
rect 139771 543218 139813 543454
rect 140049 543218 140091 543454
rect 139771 543134 140091 543218
rect 139771 542898 139813 543134
rect 140049 542898 140091 543134
rect 139771 542866 140091 542898
rect 154910 543454 155230 543486
rect 154910 543218 154952 543454
rect 155188 543218 155230 543454
rect 154910 543134 155230 543218
rect 154910 542898 154952 543134
rect 155188 542898 155230 543134
rect 154910 542866 155230 542898
rect 160840 543454 161160 543486
rect 160840 543218 160882 543454
rect 161118 543218 161160 543454
rect 160840 543134 161160 543218
rect 160840 542898 160882 543134
rect 161118 542898 161160 543134
rect 160840 542866 161160 542898
rect 166771 543454 167091 543486
rect 166771 543218 166813 543454
rect 167049 543218 167091 543454
rect 166771 543134 167091 543218
rect 166771 542898 166813 543134
rect 167049 542898 167091 543134
rect 166771 542866 167091 542898
rect 181910 543454 182230 543486
rect 181910 543218 181952 543454
rect 182188 543218 182230 543454
rect 181910 543134 182230 543218
rect 181910 542898 181952 543134
rect 182188 542898 182230 543134
rect 181910 542866 182230 542898
rect 187840 543454 188160 543486
rect 187840 543218 187882 543454
rect 188118 543218 188160 543454
rect 187840 543134 188160 543218
rect 187840 542898 187882 543134
rect 188118 542898 188160 543134
rect 187840 542866 188160 542898
rect 193771 543454 194091 543486
rect 193771 543218 193813 543454
rect 194049 543218 194091 543454
rect 193771 543134 194091 543218
rect 193771 542898 193813 543134
rect 194049 542898 194091 543134
rect 193771 542866 194091 542898
rect 208910 543454 209230 543486
rect 208910 543218 208952 543454
rect 209188 543218 209230 543454
rect 208910 543134 209230 543218
rect 208910 542898 208952 543134
rect 209188 542898 209230 543134
rect 208910 542866 209230 542898
rect 214840 543454 215160 543486
rect 214840 543218 214882 543454
rect 215118 543218 215160 543454
rect 214840 543134 215160 543218
rect 214840 542898 214882 543134
rect 215118 542898 215160 543134
rect 214840 542866 215160 542898
rect 220771 543454 221091 543486
rect 220771 543218 220813 543454
rect 221049 543218 221091 543454
rect 220771 543134 221091 543218
rect 220771 542898 220813 543134
rect 221049 542898 221091 543134
rect 220771 542866 221091 542898
rect 235910 543454 236230 543486
rect 235910 543218 235952 543454
rect 236188 543218 236230 543454
rect 235910 543134 236230 543218
rect 235910 542898 235952 543134
rect 236188 542898 236230 543134
rect 235910 542866 236230 542898
rect 241840 543454 242160 543486
rect 241840 543218 241882 543454
rect 242118 543218 242160 543454
rect 241840 543134 242160 543218
rect 241840 542898 241882 543134
rect 242118 542898 242160 543134
rect 241840 542866 242160 542898
rect 247771 543454 248091 543486
rect 247771 543218 247813 543454
rect 248049 543218 248091 543454
rect 247771 543134 248091 543218
rect 247771 542898 247813 543134
rect 248049 542898 248091 543134
rect 247771 542866 248091 542898
rect 262910 543454 263230 543486
rect 262910 543218 262952 543454
rect 263188 543218 263230 543454
rect 262910 543134 263230 543218
rect 262910 542898 262952 543134
rect 263188 542898 263230 543134
rect 262910 542866 263230 542898
rect 268840 543454 269160 543486
rect 268840 543218 268882 543454
rect 269118 543218 269160 543454
rect 268840 543134 269160 543218
rect 268840 542898 268882 543134
rect 269118 542898 269160 543134
rect 268840 542866 269160 542898
rect 274771 543454 275091 543486
rect 274771 543218 274813 543454
rect 275049 543218 275091 543454
rect 274771 543134 275091 543218
rect 274771 542898 274813 543134
rect 275049 542898 275091 543134
rect 274771 542866 275091 542898
rect 289910 543454 290230 543486
rect 289910 543218 289952 543454
rect 290188 543218 290230 543454
rect 289910 543134 290230 543218
rect 289910 542898 289952 543134
rect 290188 542898 290230 543134
rect 289910 542866 290230 542898
rect 295840 543454 296160 543486
rect 295840 543218 295882 543454
rect 296118 543218 296160 543454
rect 295840 543134 296160 543218
rect 295840 542898 295882 543134
rect 296118 542898 296160 543134
rect 295840 542866 296160 542898
rect 301771 543454 302091 543486
rect 301771 543218 301813 543454
rect 302049 543218 302091 543454
rect 301771 543134 302091 543218
rect 301771 542898 301813 543134
rect 302049 542898 302091 543134
rect 301771 542866 302091 542898
rect 316910 543454 317230 543486
rect 316910 543218 316952 543454
rect 317188 543218 317230 543454
rect 316910 543134 317230 543218
rect 316910 542898 316952 543134
rect 317188 542898 317230 543134
rect 316910 542866 317230 542898
rect 322840 543454 323160 543486
rect 322840 543218 322882 543454
rect 323118 543218 323160 543454
rect 322840 543134 323160 543218
rect 322840 542898 322882 543134
rect 323118 542898 323160 543134
rect 322840 542866 323160 542898
rect 328771 543454 329091 543486
rect 328771 543218 328813 543454
rect 329049 543218 329091 543454
rect 328771 543134 329091 543218
rect 328771 542898 328813 543134
rect 329049 542898 329091 543134
rect 328771 542866 329091 542898
rect 343910 543454 344230 543486
rect 343910 543218 343952 543454
rect 344188 543218 344230 543454
rect 343910 543134 344230 543218
rect 343910 542898 343952 543134
rect 344188 542898 344230 543134
rect 343910 542866 344230 542898
rect 349840 543454 350160 543486
rect 349840 543218 349882 543454
rect 350118 543218 350160 543454
rect 349840 543134 350160 543218
rect 349840 542898 349882 543134
rect 350118 542898 350160 543134
rect 349840 542866 350160 542898
rect 355771 543454 356091 543486
rect 355771 543218 355813 543454
rect 356049 543218 356091 543454
rect 355771 543134 356091 543218
rect 355771 542898 355813 543134
rect 356049 542898 356091 543134
rect 355771 542866 356091 542898
rect 370910 543454 371230 543486
rect 370910 543218 370952 543454
rect 371188 543218 371230 543454
rect 370910 543134 371230 543218
rect 370910 542898 370952 543134
rect 371188 542898 371230 543134
rect 370910 542866 371230 542898
rect 376840 543454 377160 543486
rect 376840 543218 376882 543454
rect 377118 543218 377160 543454
rect 376840 543134 377160 543218
rect 376840 542898 376882 543134
rect 377118 542898 377160 543134
rect 376840 542866 377160 542898
rect 382771 543454 383091 543486
rect 382771 543218 382813 543454
rect 383049 543218 383091 543454
rect 382771 543134 383091 543218
rect 382771 542898 382813 543134
rect 383049 542898 383091 543134
rect 382771 542866 383091 542898
rect 397910 543454 398230 543486
rect 397910 543218 397952 543454
rect 398188 543218 398230 543454
rect 397910 543134 398230 543218
rect 397910 542898 397952 543134
rect 398188 542898 398230 543134
rect 397910 542866 398230 542898
rect 403840 543454 404160 543486
rect 403840 543218 403882 543454
rect 404118 543218 404160 543454
rect 403840 543134 404160 543218
rect 403840 542898 403882 543134
rect 404118 542898 404160 543134
rect 403840 542866 404160 542898
rect 409771 543454 410091 543486
rect 409771 543218 409813 543454
rect 410049 543218 410091 543454
rect 409771 543134 410091 543218
rect 409771 542898 409813 543134
rect 410049 542898 410091 543134
rect 409771 542866 410091 542898
rect 424910 543454 425230 543486
rect 424910 543218 424952 543454
rect 425188 543218 425230 543454
rect 424910 543134 425230 543218
rect 424910 542898 424952 543134
rect 425188 542898 425230 543134
rect 424910 542866 425230 542898
rect 430840 543454 431160 543486
rect 430840 543218 430882 543454
rect 431118 543218 431160 543454
rect 430840 543134 431160 543218
rect 430840 542898 430882 543134
rect 431118 542898 431160 543134
rect 430840 542866 431160 542898
rect 436771 543454 437091 543486
rect 436771 543218 436813 543454
rect 437049 543218 437091 543454
rect 436771 543134 437091 543218
rect 436771 542898 436813 543134
rect 437049 542898 437091 543134
rect 436771 542866 437091 542898
rect 451910 543454 452230 543486
rect 451910 543218 451952 543454
rect 452188 543218 452230 543454
rect 451910 543134 452230 543218
rect 451910 542898 451952 543134
rect 452188 542898 452230 543134
rect 451910 542866 452230 542898
rect 457840 543454 458160 543486
rect 457840 543218 457882 543454
rect 458118 543218 458160 543454
rect 457840 543134 458160 543218
rect 457840 542898 457882 543134
rect 458118 542898 458160 543134
rect 457840 542866 458160 542898
rect 463771 543454 464091 543486
rect 463771 543218 463813 543454
rect 464049 543218 464091 543454
rect 463771 543134 464091 543218
rect 463771 542898 463813 543134
rect 464049 542898 464091 543134
rect 463771 542866 464091 542898
rect 478910 543454 479230 543486
rect 478910 543218 478952 543454
rect 479188 543218 479230 543454
rect 478910 543134 479230 543218
rect 478910 542898 478952 543134
rect 479188 542898 479230 543134
rect 478910 542866 479230 542898
rect 484840 543454 485160 543486
rect 484840 543218 484882 543454
rect 485118 543218 485160 543454
rect 484840 543134 485160 543218
rect 484840 542898 484882 543134
rect 485118 542898 485160 543134
rect 484840 542866 485160 542898
rect 490771 543454 491091 543486
rect 490771 543218 490813 543454
rect 491049 543218 491091 543454
rect 490771 543134 491091 543218
rect 490771 542898 490813 543134
rect 491049 542898 491091 543134
rect 490771 542866 491091 542898
rect 505910 543454 506230 543486
rect 505910 543218 505952 543454
rect 506188 543218 506230 543454
rect 505910 543134 506230 543218
rect 505910 542898 505952 543134
rect 506188 542898 506230 543134
rect 505910 542866 506230 542898
rect 511840 543454 512160 543486
rect 511840 543218 511882 543454
rect 512118 543218 512160 543454
rect 511840 543134 512160 543218
rect 511840 542898 511882 543134
rect 512118 542898 512160 543134
rect 511840 542866 512160 542898
rect 517771 543454 518091 543486
rect 517771 543218 517813 543454
rect 518049 543218 518091 543454
rect 517771 543134 518091 543218
rect 517771 542898 517813 543134
rect 518049 542898 518091 543134
rect 517771 542866 518091 542898
rect 532910 543454 533230 543486
rect 532910 543218 532952 543454
rect 533188 543218 533230 543454
rect 532910 543134 533230 543218
rect 532910 542898 532952 543134
rect 533188 542898 533230 543134
rect 532910 542866 533230 542898
rect 538840 543454 539160 543486
rect 538840 543218 538882 543454
rect 539118 543218 539160 543454
rect 538840 543134 539160 543218
rect 538840 542898 538882 543134
rect 539118 542898 539160 543134
rect 538840 542866 539160 542898
rect 544771 543454 545091 543486
rect 544771 543218 544813 543454
rect 545049 543218 545091 543454
rect 544771 543134 545091 543218
rect 544771 542898 544813 543134
rect 545049 542898 545091 543134
rect 544771 542866 545091 542898
rect 559794 543454 560414 560898
rect 559794 543218 559826 543454
rect 560062 543218 560146 543454
rect 560382 543218 560414 543454
rect 559794 543134 560414 543218
rect 559794 542898 559826 543134
rect 560062 542898 560146 543134
rect 560382 542898 560414 543134
rect 10794 534218 10826 534454
rect 11062 534218 11146 534454
rect 11382 534218 11414 534454
rect 10794 534134 11414 534218
rect 10794 533898 10826 534134
rect 11062 533898 11146 534134
rect 11382 533898 11414 534134
rect 10794 516454 11414 533898
rect 22874 534454 23194 534486
rect 22874 534218 22916 534454
rect 23152 534218 23194 534454
rect 22874 534134 23194 534218
rect 22874 533898 22916 534134
rect 23152 533898 23194 534134
rect 22874 533866 23194 533898
rect 28805 534454 29125 534486
rect 28805 534218 28847 534454
rect 29083 534218 29125 534454
rect 28805 534134 29125 534218
rect 28805 533898 28847 534134
rect 29083 533898 29125 534134
rect 28805 533866 29125 533898
rect 49874 534454 50194 534486
rect 49874 534218 49916 534454
rect 50152 534218 50194 534454
rect 49874 534134 50194 534218
rect 49874 533898 49916 534134
rect 50152 533898 50194 534134
rect 49874 533866 50194 533898
rect 55805 534454 56125 534486
rect 55805 534218 55847 534454
rect 56083 534218 56125 534454
rect 55805 534134 56125 534218
rect 55805 533898 55847 534134
rect 56083 533898 56125 534134
rect 55805 533866 56125 533898
rect 76874 534454 77194 534486
rect 76874 534218 76916 534454
rect 77152 534218 77194 534454
rect 76874 534134 77194 534218
rect 76874 533898 76916 534134
rect 77152 533898 77194 534134
rect 76874 533866 77194 533898
rect 82805 534454 83125 534486
rect 82805 534218 82847 534454
rect 83083 534218 83125 534454
rect 82805 534134 83125 534218
rect 82805 533898 82847 534134
rect 83083 533898 83125 534134
rect 82805 533866 83125 533898
rect 103874 534454 104194 534486
rect 103874 534218 103916 534454
rect 104152 534218 104194 534454
rect 103874 534134 104194 534218
rect 103874 533898 103916 534134
rect 104152 533898 104194 534134
rect 103874 533866 104194 533898
rect 109805 534454 110125 534486
rect 109805 534218 109847 534454
rect 110083 534218 110125 534454
rect 109805 534134 110125 534218
rect 109805 533898 109847 534134
rect 110083 533898 110125 534134
rect 109805 533866 110125 533898
rect 130874 534454 131194 534486
rect 130874 534218 130916 534454
rect 131152 534218 131194 534454
rect 130874 534134 131194 534218
rect 130874 533898 130916 534134
rect 131152 533898 131194 534134
rect 130874 533866 131194 533898
rect 136805 534454 137125 534486
rect 136805 534218 136847 534454
rect 137083 534218 137125 534454
rect 136805 534134 137125 534218
rect 136805 533898 136847 534134
rect 137083 533898 137125 534134
rect 136805 533866 137125 533898
rect 157874 534454 158194 534486
rect 157874 534218 157916 534454
rect 158152 534218 158194 534454
rect 157874 534134 158194 534218
rect 157874 533898 157916 534134
rect 158152 533898 158194 534134
rect 157874 533866 158194 533898
rect 163805 534454 164125 534486
rect 163805 534218 163847 534454
rect 164083 534218 164125 534454
rect 163805 534134 164125 534218
rect 163805 533898 163847 534134
rect 164083 533898 164125 534134
rect 163805 533866 164125 533898
rect 184874 534454 185194 534486
rect 184874 534218 184916 534454
rect 185152 534218 185194 534454
rect 184874 534134 185194 534218
rect 184874 533898 184916 534134
rect 185152 533898 185194 534134
rect 184874 533866 185194 533898
rect 190805 534454 191125 534486
rect 190805 534218 190847 534454
rect 191083 534218 191125 534454
rect 190805 534134 191125 534218
rect 190805 533898 190847 534134
rect 191083 533898 191125 534134
rect 190805 533866 191125 533898
rect 211874 534454 212194 534486
rect 211874 534218 211916 534454
rect 212152 534218 212194 534454
rect 211874 534134 212194 534218
rect 211874 533898 211916 534134
rect 212152 533898 212194 534134
rect 211874 533866 212194 533898
rect 217805 534454 218125 534486
rect 217805 534218 217847 534454
rect 218083 534218 218125 534454
rect 217805 534134 218125 534218
rect 217805 533898 217847 534134
rect 218083 533898 218125 534134
rect 217805 533866 218125 533898
rect 238874 534454 239194 534486
rect 238874 534218 238916 534454
rect 239152 534218 239194 534454
rect 238874 534134 239194 534218
rect 238874 533898 238916 534134
rect 239152 533898 239194 534134
rect 238874 533866 239194 533898
rect 244805 534454 245125 534486
rect 244805 534218 244847 534454
rect 245083 534218 245125 534454
rect 244805 534134 245125 534218
rect 244805 533898 244847 534134
rect 245083 533898 245125 534134
rect 244805 533866 245125 533898
rect 265874 534454 266194 534486
rect 265874 534218 265916 534454
rect 266152 534218 266194 534454
rect 265874 534134 266194 534218
rect 265874 533898 265916 534134
rect 266152 533898 266194 534134
rect 265874 533866 266194 533898
rect 271805 534454 272125 534486
rect 271805 534218 271847 534454
rect 272083 534218 272125 534454
rect 271805 534134 272125 534218
rect 271805 533898 271847 534134
rect 272083 533898 272125 534134
rect 271805 533866 272125 533898
rect 292874 534454 293194 534486
rect 292874 534218 292916 534454
rect 293152 534218 293194 534454
rect 292874 534134 293194 534218
rect 292874 533898 292916 534134
rect 293152 533898 293194 534134
rect 292874 533866 293194 533898
rect 298805 534454 299125 534486
rect 298805 534218 298847 534454
rect 299083 534218 299125 534454
rect 298805 534134 299125 534218
rect 298805 533898 298847 534134
rect 299083 533898 299125 534134
rect 298805 533866 299125 533898
rect 319874 534454 320194 534486
rect 319874 534218 319916 534454
rect 320152 534218 320194 534454
rect 319874 534134 320194 534218
rect 319874 533898 319916 534134
rect 320152 533898 320194 534134
rect 319874 533866 320194 533898
rect 325805 534454 326125 534486
rect 325805 534218 325847 534454
rect 326083 534218 326125 534454
rect 325805 534134 326125 534218
rect 325805 533898 325847 534134
rect 326083 533898 326125 534134
rect 325805 533866 326125 533898
rect 346874 534454 347194 534486
rect 346874 534218 346916 534454
rect 347152 534218 347194 534454
rect 346874 534134 347194 534218
rect 346874 533898 346916 534134
rect 347152 533898 347194 534134
rect 346874 533866 347194 533898
rect 352805 534454 353125 534486
rect 352805 534218 352847 534454
rect 353083 534218 353125 534454
rect 352805 534134 353125 534218
rect 352805 533898 352847 534134
rect 353083 533898 353125 534134
rect 352805 533866 353125 533898
rect 373874 534454 374194 534486
rect 373874 534218 373916 534454
rect 374152 534218 374194 534454
rect 373874 534134 374194 534218
rect 373874 533898 373916 534134
rect 374152 533898 374194 534134
rect 373874 533866 374194 533898
rect 379805 534454 380125 534486
rect 379805 534218 379847 534454
rect 380083 534218 380125 534454
rect 379805 534134 380125 534218
rect 379805 533898 379847 534134
rect 380083 533898 380125 534134
rect 379805 533866 380125 533898
rect 400874 534454 401194 534486
rect 400874 534218 400916 534454
rect 401152 534218 401194 534454
rect 400874 534134 401194 534218
rect 400874 533898 400916 534134
rect 401152 533898 401194 534134
rect 400874 533866 401194 533898
rect 406805 534454 407125 534486
rect 406805 534218 406847 534454
rect 407083 534218 407125 534454
rect 406805 534134 407125 534218
rect 406805 533898 406847 534134
rect 407083 533898 407125 534134
rect 406805 533866 407125 533898
rect 427874 534454 428194 534486
rect 427874 534218 427916 534454
rect 428152 534218 428194 534454
rect 427874 534134 428194 534218
rect 427874 533898 427916 534134
rect 428152 533898 428194 534134
rect 427874 533866 428194 533898
rect 433805 534454 434125 534486
rect 433805 534218 433847 534454
rect 434083 534218 434125 534454
rect 433805 534134 434125 534218
rect 433805 533898 433847 534134
rect 434083 533898 434125 534134
rect 433805 533866 434125 533898
rect 454874 534454 455194 534486
rect 454874 534218 454916 534454
rect 455152 534218 455194 534454
rect 454874 534134 455194 534218
rect 454874 533898 454916 534134
rect 455152 533898 455194 534134
rect 454874 533866 455194 533898
rect 460805 534454 461125 534486
rect 460805 534218 460847 534454
rect 461083 534218 461125 534454
rect 460805 534134 461125 534218
rect 460805 533898 460847 534134
rect 461083 533898 461125 534134
rect 460805 533866 461125 533898
rect 481874 534454 482194 534486
rect 481874 534218 481916 534454
rect 482152 534218 482194 534454
rect 481874 534134 482194 534218
rect 481874 533898 481916 534134
rect 482152 533898 482194 534134
rect 481874 533866 482194 533898
rect 487805 534454 488125 534486
rect 487805 534218 487847 534454
rect 488083 534218 488125 534454
rect 487805 534134 488125 534218
rect 487805 533898 487847 534134
rect 488083 533898 488125 534134
rect 487805 533866 488125 533898
rect 508874 534454 509194 534486
rect 508874 534218 508916 534454
rect 509152 534218 509194 534454
rect 508874 534134 509194 534218
rect 508874 533898 508916 534134
rect 509152 533898 509194 534134
rect 508874 533866 509194 533898
rect 514805 534454 515125 534486
rect 514805 534218 514847 534454
rect 515083 534218 515125 534454
rect 514805 534134 515125 534218
rect 514805 533898 514847 534134
rect 515083 533898 515125 534134
rect 514805 533866 515125 533898
rect 535874 534454 536194 534486
rect 535874 534218 535916 534454
rect 536152 534218 536194 534454
rect 535874 534134 536194 534218
rect 535874 533898 535916 534134
rect 536152 533898 536194 534134
rect 535874 533866 536194 533898
rect 541805 534454 542125 534486
rect 541805 534218 541847 534454
rect 542083 534218 542125 534454
rect 541805 534134 542125 534218
rect 541805 533898 541847 534134
rect 542083 533898 542125 534134
rect 541805 533866 542125 533898
rect 19794 525454 20414 527000
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 524000 20414 524898
rect 28794 526394 29414 527000
rect 28794 526158 28826 526394
rect 29062 526158 29146 526394
rect 29382 526158 29414 526394
rect 28794 526074 29414 526158
rect 28794 525838 28826 526074
rect 29062 525838 29146 526074
rect 29382 525838 29414 526074
rect 28794 524000 29414 525838
rect 37794 525454 38414 527000
rect 37794 525218 37826 525454
rect 38062 525218 38146 525454
rect 38382 525218 38414 525454
rect 37794 525134 38414 525218
rect 37794 524898 37826 525134
rect 38062 524898 38146 525134
rect 38382 524898 38414 525134
rect 37794 524000 38414 524898
rect 46794 526394 47414 527000
rect 46794 526158 46826 526394
rect 47062 526158 47146 526394
rect 47382 526158 47414 526394
rect 46794 526074 47414 526158
rect 46794 525838 46826 526074
rect 47062 525838 47146 526074
rect 47382 525838 47414 526074
rect 46794 524000 47414 525838
rect 55794 525454 56414 527000
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 524000 56414 524898
rect 64794 526394 65414 527000
rect 64794 526158 64826 526394
rect 65062 526158 65146 526394
rect 65382 526158 65414 526394
rect 64794 526074 65414 526158
rect 64794 525838 64826 526074
rect 65062 525838 65146 526074
rect 65382 525838 65414 526074
rect 64794 524000 65414 525838
rect 73794 525454 74414 527000
rect 73794 525218 73826 525454
rect 74062 525218 74146 525454
rect 74382 525218 74414 525454
rect 73794 525134 74414 525218
rect 73794 524898 73826 525134
rect 74062 524898 74146 525134
rect 74382 524898 74414 525134
rect 73794 524000 74414 524898
rect 82794 526394 83414 527000
rect 82794 526158 82826 526394
rect 83062 526158 83146 526394
rect 83382 526158 83414 526394
rect 82794 526074 83414 526158
rect 82794 525838 82826 526074
rect 83062 525838 83146 526074
rect 83382 525838 83414 526074
rect 82794 524000 83414 525838
rect 91794 525454 92414 527000
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 524000 92414 524898
rect 100794 526394 101414 527000
rect 100794 526158 100826 526394
rect 101062 526158 101146 526394
rect 101382 526158 101414 526394
rect 100794 526074 101414 526158
rect 100794 525838 100826 526074
rect 101062 525838 101146 526074
rect 101382 525838 101414 526074
rect 100794 524000 101414 525838
rect 109794 525454 110414 527000
rect 109794 525218 109826 525454
rect 110062 525218 110146 525454
rect 110382 525218 110414 525454
rect 109794 525134 110414 525218
rect 109794 524898 109826 525134
rect 110062 524898 110146 525134
rect 110382 524898 110414 525134
rect 109794 524000 110414 524898
rect 118794 526394 119414 527000
rect 118794 526158 118826 526394
rect 119062 526158 119146 526394
rect 119382 526158 119414 526394
rect 118794 526074 119414 526158
rect 118794 525838 118826 526074
rect 119062 525838 119146 526074
rect 119382 525838 119414 526074
rect 118794 524000 119414 525838
rect 127794 525454 128414 527000
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 524000 128414 524898
rect 136794 526394 137414 527000
rect 136794 526158 136826 526394
rect 137062 526158 137146 526394
rect 137382 526158 137414 526394
rect 136794 526074 137414 526158
rect 136794 525838 136826 526074
rect 137062 525838 137146 526074
rect 137382 525838 137414 526074
rect 136794 524000 137414 525838
rect 145794 525454 146414 527000
rect 145794 525218 145826 525454
rect 146062 525218 146146 525454
rect 146382 525218 146414 525454
rect 145794 525134 146414 525218
rect 145794 524898 145826 525134
rect 146062 524898 146146 525134
rect 146382 524898 146414 525134
rect 145794 524000 146414 524898
rect 154794 526394 155414 527000
rect 154794 526158 154826 526394
rect 155062 526158 155146 526394
rect 155382 526158 155414 526394
rect 154794 526074 155414 526158
rect 154794 525838 154826 526074
rect 155062 525838 155146 526074
rect 155382 525838 155414 526074
rect 154794 524000 155414 525838
rect 163794 525454 164414 527000
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 524000 164414 524898
rect 172794 526394 173414 527000
rect 172794 526158 172826 526394
rect 173062 526158 173146 526394
rect 173382 526158 173414 526394
rect 172794 526074 173414 526158
rect 172794 525838 172826 526074
rect 173062 525838 173146 526074
rect 173382 525838 173414 526074
rect 172794 524000 173414 525838
rect 181794 525454 182414 527000
rect 181794 525218 181826 525454
rect 182062 525218 182146 525454
rect 182382 525218 182414 525454
rect 181794 525134 182414 525218
rect 181794 524898 181826 525134
rect 182062 524898 182146 525134
rect 182382 524898 182414 525134
rect 181794 524000 182414 524898
rect 190794 526394 191414 527000
rect 190794 526158 190826 526394
rect 191062 526158 191146 526394
rect 191382 526158 191414 526394
rect 190794 526074 191414 526158
rect 190794 525838 190826 526074
rect 191062 525838 191146 526074
rect 191382 525838 191414 526074
rect 190794 524000 191414 525838
rect 199794 525454 200414 527000
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 524000 200414 524898
rect 208794 526394 209414 527000
rect 208794 526158 208826 526394
rect 209062 526158 209146 526394
rect 209382 526158 209414 526394
rect 208794 526074 209414 526158
rect 208794 525838 208826 526074
rect 209062 525838 209146 526074
rect 209382 525838 209414 526074
rect 208794 524000 209414 525838
rect 217794 525454 218414 527000
rect 217794 525218 217826 525454
rect 218062 525218 218146 525454
rect 218382 525218 218414 525454
rect 217794 525134 218414 525218
rect 217794 524898 217826 525134
rect 218062 524898 218146 525134
rect 218382 524898 218414 525134
rect 217794 524000 218414 524898
rect 226794 526394 227414 527000
rect 226794 526158 226826 526394
rect 227062 526158 227146 526394
rect 227382 526158 227414 526394
rect 226794 526074 227414 526158
rect 226794 525838 226826 526074
rect 227062 525838 227146 526074
rect 227382 525838 227414 526074
rect 226794 524000 227414 525838
rect 235794 525454 236414 527000
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 524000 236414 524898
rect 244794 526394 245414 527000
rect 244794 526158 244826 526394
rect 245062 526158 245146 526394
rect 245382 526158 245414 526394
rect 244794 526074 245414 526158
rect 244794 525838 244826 526074
rect 245062 525838 245146 526074
rect 245382 525838 245414 526074
rect 244794 524000 245414 525838
rect 253794 525454 254414 527000
rect 253794 525218 253826 525454
rect 254062 525218 254146 525454
rect 254382 525218 254414 525454
rect 253794 525134 254414 525218
rect 253794 524898 253826 525134
rect 254062 524898 254146 525134
rect 254382 524898 254414 525134
rect 253794 524000 254414 524898
rect 262794 526394 263414 527000
rect 262794 526158 262826 526394
rect 263062 526158 263146 526394
rect 263382 526158 263414 526394
rect 262794 526074 263414 526158
rect 262794 525838 262826 526074
rect 263062 525838 263146 526074
rect 263382 525838 263414 526074
rect 262794 524000 263414 525838
rect 271794 525454 272414 527000
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 524000 272414 524898
rect 280794 526394 281414 527000
rect 280794 526158 280826 526394
rect 281062 526158 281146 526394
rect 281382 526158 281414 526394
rect 280794 526074 281414 526158
rect 280794 525838 280826 526074
rect 281062 525838 281146 526074
rect 281382 525838 281414 526074
rect 280794 524000 281414 525838
rect 289794 525454 290414 527000
rect 289794 525218 289826 525454
rect 290062 525218 290146 525454
rect 290382 525218 290414 525454
rect 289794 525134 290414 525218
rect 289794 524898 289826 525134
rect 290062 524898 290146 525134
rect 290382 524898 290414 525134
rect 289794 524000 290414 524898
rect 298794 526394 299414 527000
rect 298794 526158 298826 526394
rect 299062 526158 299146 526394
rect 299382 526158 299414 526394
rect 298794 526074 299414 526158
rect 298794 525838 298826 526074
rect 299062 525838 299146 526074
rect 299382 525838 299414 526074
rect 298794 524000 299414 525838
rect 307794 525454 308414 527000
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 524000 308414 524898
rect 316794 526394 317414 527000
rect 316794 526158 316826 526394
rect 317062 526158 317146 526394
rect 317382 526158 317414 526394
rect 316794 526074 317414 526158
rect 316794 525838 316826 526074
rect 317062 525838 317146 526074
rect 317382 525838 317414 526074
rect 316794 524000 317414 525838
rect 325794 525454 326414 527000
rect 325794 525218 325826 525454
rect 326062 525218 326146 525454
rect 326382 525218 326414 525454
rect 325794 525134 326414 525218
rect 325794 524898 325826 525134
rect 326062 524898 326146 525134
rect 326382 524898 326414 525134
rect 325794 524000 326414 524898
rect 334794 526394 335414 527000
rect 334794 526158 334826 526394
rect 335062 526158 335146 526394
rect 335382 526158 335414 526394
rect 334794 526074 335414 526158
rect 334794 525838 334826 526074
rect 335062 525838 335146 526074
rect 335382 525838 335414 526074
rect 334794 524000 335414 525838
rect 343794 525454 344414 527000
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 524000 344414 524898
rect 352794 526394 353414 527000
rect 352794 526158 352826 526394
rect 353062 526158 353146 526394
rect 353382 526158 353414 526394
rect 352794 526074 353414 526158
rect 352794 525838 352826 526074
rect 353062 525838 353146 526074
rect 353382 525838 353414 526074
rect 352794 524000 353414 525838
rect 361794 525454 362414 527000
rect 361794 525218 361826 525454
rect 362062 525218 362146 525454
rect 362382 525218 362414 525454
rect 361794 525134 362414 525218
rect 361794 524898 361826 525134
rect 362062 524898 362146 525134
rect 362382 524898 362414 525134
rect 361794 524000 362414 524898
rect 370794 526394 371414 527000
rect 370794 526158 370826 526394
rect 371062 526158 371146 526394
rect 371382 526158 371414 526394
rect 370794 526074 371414 526158
rect 370794 525838 370826 526074
rect 371062 525838 371146 526074
rect 371382 525838 371414 526074
rect 370794 524000 371414 525838
rect 379794 525454 380414 527000
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 524000 380414 524898
rect 388794 526394 389414 527000
rect 388794 526158 388826 526394
rect 389062 526158 389146 526394
rect 389382 526158 389414 526394
rect 388794 526074 389414 526158
rect 388794 525838 388826 526074
rect 389062 525838 389146 526074
rect 389382 525838 389414 526074
rect 388794 524000 389414 525838
rect 397794 525454 398414 527000
rect 397794 525218 397826 525454
rect 398062 525218 398146 525454
rect 398382 525218 398414 525454
rect 397794 525134 398414 525218
rect 397794 524898 397826 525134
rect 398062 524898 398146 525134
rect 398382 524898 398414 525134
rect 397794 524000 398414 524898
rect 406794 526394 407414 527000
rect 406794 526158 406826 526394
rect 407062 526158 407146 526394
rect 407382 526158 407414 526394
rect 406794 526074 407414 526158
rect 406794 525838 406826 526074
rect 407062 525838 407146 526074
rect 407382 525838 407414 526074
rect 406794 524000 407414 525838
rect 415794 525454 416414 527000
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 524000 416414 524898
rect 424794 526394 425414 527000
rect 424794 526158 424826 526394
rect 425062 526158 425146 526394
rect 425382 526158 425414 526394
rect 424794 526074 425414 526158
rect 424794 525838 424826 526074
rect 425062 525838 425146 526074
rect 425382 525838 425414 526074
rect 424794 524000 425414 525838
rect 433794 525454 434414 527000
rect 433794 525218 433826 525454
rect 434062 525218 434146 525454
rect 434382 525218 434414 525454
rect 433794 525134 434414 525218
rect 433794 524898 433826 525134
rect 434062 524898 434146 525134
rect 434382 524898 434414 525134
rect 433794 524000 434414 524898
rect 442794 526394 443414 527000
rect 442794 526158 442826 526394
rect 443062 526158 443146 526394
rect 443382 526158 443414 526394
rect 442794 526074 443414 526158
rect 442794 525838 442826 526074
rect 443062 525838 443146 526074
rect 443382 525838 443414 526074
rect 442794 524000 443414 525838
rect 451794 525454 452414 527000
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 524000 452414 524898
rect 460794 526394 461414 527000
rect 460794 526158 460826 526394
rect 461062 526158 461146 526394
rect 461382 526158 461414 526394
rect 460794 526074 461414 526158
rect 460794 525838 460826 526074
rect 461062 525838 461146 526074
rect 461382 525838 461414 526074
rect 460794 524000 461414 525838
rect 469794 525454 470414 527000
rect 469794 525218 469826 525454
rect 470062 525218 470146 525454
rect 470382 525218 470414 525454
rect 469794 525134 470414 525218
rect 469794 524898 469826 525134
rect 470062 524898 470146 525134
rect 470382 524898 470414 525134
rect 469794 524000 470414 524898
rect 478794 526394 479414 527000
rect 478794 526158 478826 526394
rect 479062 526158 479146 526394
rect 479382 526158 479414 526394
rect 478794 526074 479414 526158
rect 478794 525838 478826 526074
rect 479062 525838 479146 526074
rect 479382 525838 479414 526074
rect 478794 524000 479414 525838
rect 487794 525454 488414 527000
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 524000 488414 524898
rect 496794 526394 497414 527000
rect 496794 526158 496826 526394
rect 497062 526158 497146 526394
rect 497382 526158 497414 526394
rect 496794 526074 497414 526158
rect 496794 525838 496826 526074
rect 497062 525838 497146 526074
rect 497382 525838 497414 526074
rect 496794 524000 497414 525838
rect 505794 525454 506414 527000
rect 505794 525218 505826 525454
rect 506062 525218 506146 525454
rect 506382 525218 506414 525454
rect 505794 525134 506414 525218
rect 505794 524898 505826 525134
rect 506062 524898 506146 525134
rect 506382 524898 506414 525134
rect 505794 524000 506414 524898
rect 514794 526394 515414 527000
rect 514794 526158 514826 526394
rect 515062 526158 515146 526394
rect 515382 526158 515414 526394
rect 514794 526074 515414 526158
rect 514794 525838 514826 526074
rect 515062 525838 515146 526074
rect 515382 525838 515414 526074
rect 514794 524000 515414 525838
rect 523794 525454 524414 527000
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 524000 524414 524898
rect 532794 526394 533414 527000
rect 532794 526158 532826 526394
rect 533062 526158 533146 526394
rect 533382 526158 533414 526394
rect 532794 526074 533414 526158
rect 532794 525838 532826 526074
rect 533062 525838 533146 526074
rect 533382 525838 533414 526074
rect 532794 524000 533414 525838
rect 541794 525454 542414 527000
rect 541794 525218 541826 525454
rect 542062 525218 542146 525454
rect 542382 525218 542414 525454
rect 541794 525134 542414 525218
rect 541794 524898 541826 525134
rect 542062 524898 542146 525134
rect 542382 524898 542414 525134
rect 541794 524000 542414 524898
rect 550794 526394 551414 527000
rect 550794 526158 550826 526394
rect 551062 526158 551146 526394
rect 551382 526158 551414 526394
rect 550794 526074 551414 526158
rect 550794 525838 550826 526074
rect 551062 525838 551146 526074
rect 551382 525838 551414 526074
rect 550794 524000 551414 525838
rect 559794 525454 560414 542898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 498454 11414 515898
rect 22874 516454 23194 516486
rect 22874 516218 22916 516454
rect 23152 516218 23194 516454
rect 22874 516134 23194 516218
rect 22874 515898 22916 516134
rect 23152 515898 23194 516134
rect 22874 515866 23194 515898
rect 28805 516454 29125 516486
rect 28805 516218 28847 516454
rect 29083 516218 29125 516454
rect 28805 516134 29125 516218
rect 28805 515898 28847 516134
rect 29083 515898 29125 516134
rect 28805 515866 29125 515898
rect 49874 516454 50194 516486
rect 49874 516218 49916 516454
rect 50152 516218 50194 516454
rect 49874 516134 50194 516218
rect 49874 515898 49916 516134
rect 50152 515898 50194 516134
rect 49874 515866 50194 515898
rect 55805 516454 56125 516486
rect 55805 516218 55847 516454
rect 56083 516218 56125 516454
rect 55805 516134 56125 516218
rect 55805 515898 55847 516134
rect 56083 515898 56125 516134
rect 55805 515866 56125 515898
rect 76874 516454 77194 516486
rect 76874 516218 76916 516454
rect 77152 516218 77194 516454
rect 76874 516134 77194 516218
rect 76874 515898 76916 516134
rect 77152 515898 77194 516134
rect 76874 515866 77194 515898
rect 82805 516454 83125 516486
rect 82805 516218 82847 516454
rect 83083 516218 83125 516454
rect 82805 516134 83125 516218
rect 82805 515898 82847 516134
rect 83083 515898 83125 516134
rect 82805 515866 83125 515898
rect 103874 516454 104194 516486
rect 103874 516218 103916 516454
rect 104152 516218 104194 516454
rect 103874 516134 104194 516218
rect 103874 515898 103916 516134
rect 104152 515898 104194 516134
rect 103874 515866 104194 515898
rect 109805 516454 110125 516486
rect 109805 516218 109847 516454
rect 110083 516218 110125 516454
rect 109805 516134 110125 516218
rect 109805 515898 109847 516134
rect 110083 515898 110125 516134
rect 109805 515866 110125 515898
rect 130874 516454 131194 516486
rect 130874 516218 130916 516454
rect 131152 516218 131194 516454
rect 130874 516134 131194 516218
rect 130874 515898 130916 516134
rect 131152 515898 131194 516134
rect 130874 515866 131194 515898
rect 136805 516454 137125 516486
rect 136805 516218 136847 516454
rect 137083 516218 137125 516454
rect 136805 516134 137125 516218
rect 136805 515898 136847 516134
rect 137083 515898 137125 516134
rect 136805 515866 137125 515898
rect 157874 516454 158194 516486
rect 157874 516218 157916 516454
rect 158152 516218 158194 516454
rect 157874 516134 158194 516218
rect 157874 515898 157916 516134
rect 158152 515898 158194 516134
rect 157874 515866 158194 515898
rect 163805 516454 164125 516486
rect 163805 516218 163847 516454
rect 164083 516218 164125 516454
rect 163805 516134 164125 516218
rect 163805 515898 163847 516134
rect 164083 515898 164125 516134
rect 163805 515866 164125 515898
rect 184874 516454 185194 516486
rect 184874 516218 184916 516454
rect 185152 516218 185194 516454
rect 184874 516134 185194 516218
rect 184874 515898 184916 516134
rect 185152 515898 185194 516134
rect 184874 515866 185194 515898
rect 190805 516454 191125 516486
rect 190805 516218 190847 516454
rect 191083 516218 191125 516454
rect 190805 516134 191125 516218
rect 190805 515898 190847 516134
rect 191083 515898 191125 516134
rect 190805 515866 191125 515898
rect 211874 516454 212194 516486
rect 211874 516218 211916 516454
rect 212152 516218 212194 516454
rect 211874 516134 212194 516218
rect 211874 515898 211916 516134
rect 212152 515898 212194 516134
rect 211874 515866 212194 515898
rect 217805 516454 218125 516486
rect 217805 516218 217847 516454
rect 218083 516218 218125 516454
rect 217805 516134 218125 516218
rect 217805 515898 217847 516134
rect 218083 515898 218125 516134
rect 217805 515866 218125 515898
rect 238874 516454 239194 516486
rect 238874 516218 238916 516454
rect 239152 516218 239194 516454
rect 238874 516134 239194 516218
rect 238874 515898 238916 516134
rect 239152 515898 239194 516134
rect 238874 515866 239194 515898
rect 244805 516454 245125 516486
rect 244805 516218 244847 516454
rect 245083 516218 245125 516454
rect 244805 516134 245125 516218
rect 244805 515898 244847 516134
rect 245083 515898 245125 516134
rect 244805 515866 245125 515898
rect 265874 516454 266194 516486
rect 265874 516218 265916 516454
rect 266152 516218 266194 516454
rect 265874 516134 266194 516218
rect 265874 515898 265916 516134
rect 266152 515898 266194 516134
rect 265874 515866 266194 515898
rect 271805 516454 272125 516486
rect 271805 516218 271847 516454
rect 272083 516218 272125 516454
rect 271805 516134 272125 516218
rect 271805 515898 271847 516134
rect 272083 515898 272125 516134
rect 271805 515866 272125 515898
rect 292874 516454 293194 516486
rect 292874 516218 292916 516454
rect 293152 516218 293194 516454
rect 292874 516134 293194 516218
rect 292874 515898 292916 516134
rect 293152 515898 293194 516134
rect 292874 515866 293194 515898
rect 298805 516454 299125 516486
rect 298805 516218 298847 516454
rect 299083 516218 299125 516454
rect 298805 516134 299125 516218
rect 298805 515898 298847 516134
rect 299083 515898 299125 516134
rect 298805 515866 299125 515898
rect 319874 516454 320194 516486
rect 319874 516218 319916 516454
rect 320152 516218 320194 516454
rect 319874 516134 320194 516218
rect 319874 515898 319916 516134
rect 320152 515898 320194 516134
rect 319874 515866 320194 515898
rect 325805 516454 326125 516486
rect 325805 516218 325847 516454
rect 326083 516218 326125 516454
rect 325805 516134 326125 516218
rect 325805 515898 325847 516134
rect 326083 515898 326125 516134
rect 325805 515866 326125 515898
rect 346874 516454 347194 516486
rect 346874 516218 346916 516454
rect 347152 516218 347194 516454
rect 346874 516134 347194 516218
rect 346874 515898 346916 516134
rect 347152 515898 347194 516134
rect 346874 515866 347194 515898
rect 352805 516454 353125 516486
rect 352805 516218 352847 516454
rect 353083 516218 353125 516454
rect 352805 516134 353125 516218
rect 352805 515898 352847 516134
rect 353083 515898 353125 516134
rect 352805 515866 353125 515898
rect 373874 516454 374194 516486
rect 373874 516218 373916 516454
rect 374152 516218 374194 516454
rect 373874 516134 374194 516218
rect 373874 515898 373916 516134
rect 374152 515898 374194 516134
rect 373874 515866 374194 515898
rect 379805 516454 380125 516486
rect 379805 516218 379847 516454
rect 380083 516218 380125 516454
rect 379805 516134 380125 516218
rect 379805 515898 379847 516134
rect 380083 515898 380125 516134
rect 379805 515866 380125 515898
rect 400874 516454 401194 516486
rect 400874 516218 400916 516454
rect 401152 516218 401194 516454
rect 400874 516134 401194 516218
rect 400874 515898 400916 516134
rect 401152 515898 401194 516134
rect 400874 515866 401194 515898
rect 406805 516454 407125 516486
rect 406805 516218 406847 516454
rect 407083 516218 407125 516454
rect 406805 516134 407125 516218
rect 406805 515898 406847 516134
rect 407083 515898 407125 516134
rect 406805 515866 407125 515898
rect 427874 516454 428194 516486
rect 427874 516218 427916 516454
rect 428152 516218 428194 516454
rect 427874 516134 428194 516218
rect 427874 515898 427916 516134
rect 428152 515898 428194 516134
rect 427874 515866 428194 515898
rect 433805 516454 434125 516486
rect 433805 516218 433847 516454
rect 434083 516218 434125 516454
rect 433805 516134 434125 516218
rect 433805 515898 433847 516134
rect 434083 515898 434125 516134
rect 433805 515866 434125 515898
rect 454874 516454 455194 516486
rect 454874 516218 454916 516454
rect 455152 516218 455194 516454
rect 454874 516134 455194 516218
rect 454874 515898 454916 516134
rect 455152 515898 455194 516134
rect 454874 515866 455194 515898
rect 460805 516454 461125 516486
rect 460805 516218 460847 516454
rect 461083 516218 461125 516454
rect 460805 516134 461125 516218
rect 460805 515898 460847 516134
rect 461083 515898 461125 516134
rect 460805 515866 461125 515898
rect 481874 516454 482194 516486
rect 481874 516218 481916 516454
rect 482152 516218 482194 516454
rect 481874 516134 482194 516218
rect 481874 515898 481916 516134
rect 482152 515898 482194 516134
rect 481874 515866 482194 515898
rect 487805 516454 488125 516486
rect 487805 516218 487847 516454
rect 488083 516218 488125 516454
rect 487805 516134 488125 516218
rect 487805 515898 487847 516134
rect 488083 515898 488125 516134
rect 487805 515866 488125 515898
rect 508874 516454 509194 516486
rect 508874 516218 508916 516454
rect 509152 516218 509194 516454
rect 508874 516134 509194 516218
rect 508874 515898 508916 516134
rect 509152 515898 509194 516134
rect 508874 515866 509194 515898
rect 514805 516454 515125 516486
rect 514805 516218 514847 516454
rect 515083 516218 515125 516454
rect 514805 516134 515125 516218
rect 514805 515898 514847 516134
rect 515083 515898 515125 516134
rect 514805 515866 515125 515898
rect 535874 516454 536194 516486
rect 535874 516218 535916 516454
rect 536152 516218 536194 516454
rect 535874 516134 536194 516218
rect 535874 515898 535916 516134
rect 536152 515898 536194 516134
rect 535874 515866 536194 515898
rect 541805 516454 542125 516486
rect 541805 516218 541847 516454
rect 542083 516218 542125 516454
rect 541805 516134 542125 516218
rect 541805 515898 541847 516134
rect 542083 515898 542125 516134
rect 541805 515866 542125 515898
rect 19910 507454 20230 507486
rect 19910 507218 19952 507454
rect 20188 507218 20230 507454
rect 19910 507134 20230 507218
rect 19910 506898 19952 507134
rect 20188 506898 20230 507134
rect 19910 506866 20230 506898
rect 25840 507454 26160 507486
rect 25840 507218 25882 507454
rect 26118 507218 26160 507454
rect 25840 507134 26160 507218
rect 25840 506898 25882 507134
rect 26118 506898 26160 507134
rect 25840 506866 26160 506898
rect 31771 507454 32091 507486
rect 31771 507218 31813 507454
rect 32049 507218 32091 507454
rect 31771 507134 32091 507218
rect 31771 506898 31813 507134
rect 32049 506898 32091 507134
rect 31771 506866 32091 506898
rect 46910 507454 47230 507486
rect 46910 507218 46952 507454
rect 47188 507218 47230 507454
rect 46910 507134 47230 507218
rect 46910 506898 46952 507134
rect 47188 506898 47230 507134
rect 46910 506866 47230 506898
rect 52840 507454 53160 507486
rect 52840 507218 52882 507454
rect 53118 507218 53160 507454
rect 52840 507134 53160 507218
rect 52840 506898 52882 507134
rect 53118 506898 53160 507134
rect 52840 506866 53160 506898
rect 58771 507454 59091 507486
rect 58771 507218 58813 507454
rect 59049 507218 59091 507454
rect 58771 507134 59091 507218
rect 58771 506898 58813 507134
rect 59049 506898 59091 507134
rect 58771 506866 59091 506898
rect 73910 507454 74230 507486
rect 73910 507218 73952 507454
rect 74188 507218 74230 507454
rect 73910 507134 74230 507218
rect 73910 506898 73952 507134
rect 74188 506898 74230 507134
rect 73910 506866 74230 506898
rect 79840 507454 80160 507486
rect 79840 507218 79882 507454
rect 80118 507218 80160 507454
rect 79840 507134 80160 507218
rect 79840 506898 79882 507134
rect 80118 506898 80160 507134
rect 79840 506866 80160 506898
rect 85771 507454 86091 507486
rect 85771 507218 85813 507454
rect 86049 507218 86091 507454
rect 85771 507134 86091 507218
rect 85771 506898 85813 507134
rect 86049 506898 86091 507134
rect 85771 506866 86091 506898
rect 100910 507454 101230 507486
rect 100910 507218 100952 507454
rect 101188 507218 101230 507454
rect 100910 507134 101230 507218
rect 100910 506898 100952 507134
rect 101188 506898 101230 507134
rect 100910 506866 101230 506898
rect 106840 507454 107160 507486
rect 106840 507218 106882 507454
rect 107118 507218 107160 507454
rect 106840 507134 107160 507218
rect 106840 506898 106882 507134
rect 107118 506898 107160 507134
rect 106840 506866 107160 506898
rect 112771 507454 113091 507486
rect 112771 507218 112813 507454
rect 113049 507218 113091 507454
rect 112771 507134 113091 507218
rect 112771 506898 112813 507134
rect 113049 506898 113091 507134
rect 112771 506866 113091 506898
rect 127910 507454 128230 507486
rect 127910 507218 127952 507454
rect 128188 507218 128230 507454
rect 127910 507134 128230 507218
rect 127910 506898 127952 507134
rect 128188 506898 128230 507134
rect 127910 506866 128230 506898
rect 133840 507454 134160 507486
rect 133840 507218 133882 507454
rect 134118 507218 134160 507454
rect 133840 507134 134160 507218
rect 133840 506898 133882 507134
rect 134118 506898 134160 507134
rect 133840 506866 134160 506898
rect 139771 507454 140091 507486
rect 139771 507218 139813 507454
rect 140049 507218 140091 507454
rect 139771 507134 140091 507218
rect 139771 506898 139813 507134
rect 140049 506898 140091 507134
rect 139771 506866 140091 506898
rect 154910 507454 155230 507486
rect 154910 507218 154952 507454
rect 155188 507218 155230 507454
rect 154910 507134 155230 507218
rect 154910 506898 154952 507134
rect 155188 506898 155230 507134
rect 154910 506866 155230 506898
rect 160840 507454 161160 507486
rect 160840 507218 160882 507454
rect 161118 507218 161160 507454
rect 160840 507134 161160 507218
rect 160840 506898 160882 507134
rect 161118 506898 161160 507134
rect 160840 506866 161160 506898
rect 166771 507454 167091 507486
rect 166771 507218 166813 507454
rect 167049 507218 167091 507454
rect 166771 507134 167091 507218
rect 166771 506898 166813 507134
rect 167049 506898 167091 507134
rect 166771 506866 167091 506898
rect 181910 507454 182230 507486
rect 181910 507218 181952 507454
rect 182188 507218 182230 507454
rect 181910 507134 182230 507218
rect 181910 506898 181952 507134
rect 182188 506898 182230 507134
rect 181910 506866 182230 506898
rect 187840 507454 188160 507486
rect 187840 507218 187882 507454
rect 188118 507218 188160 507454
rect 187840 507134 188160 507218
rect 187840 506898 187882 507134
rect 188118 506898 188160 507134
rect 187840 506866 188160 506898
rect 193771 507454 194091 507486
rect 193771 507218 193813 507454
rect 194049 507218 194091 507454
rect 193771 507134 194091 507218
rect 193771 506898 193813 507134
rect 194049 506898 194091 507134
rect 193771 506866 194091 506898
rect 208910 507454 209230 507486
rect 208910 507218 208952 507454
rect 209188 507218 209230 507454
rect 208910 507134 209230 507218
rect 208910 506898 208952 507134
rect 209188 506898 209230 507134
rect 208910 506866 209230 506898
rect 214840 507454 215160 507486
rect 214840 507218 214882 507454
rect 215118 507218 215160 507454
rect 214840 507134 215160 507218
rect 214840 506898 214882 507134
rect 215118 506898 215160 507134
rect 214840 506866 215160 506898
rect 220771 507454 221091 507486
rect 220771 507218 220813 507454
rect 221049 507218 221091 507454
rect 220771 507134 221091 507218
rect 220771 506898 220813 507134
rect 221049 506898 221091 507134
rect 220771 506866 221091 506898
rect 235910 507454 236230 507486
rect 235910 507218 235952 507454
rect 236188 507218 236230 507454
rect 235910 507134 236230 507218
rect 235910 506898 235952 507134
rect 236188 506898 236230 507134
rect 235910 506866 236230 506898
rect 241840 507454 242160 507486
rect 241840 507218 241882 507454
rect 242118 507218 242160 507454
rect 241840 507134 242160 507218
rect 241840 506898 241882 507134
rect 242118 506898 242160 507134
rect 241840 506866 242160 506898
rect 247771 507454 248091 507486
rect 247771 507218 247813 507454
rect 248049 507218 248091 507454
rect 247771 507134 248091 507218
rect 247771 506898 247813 507134
rect 248049 506898 248091 507134
rect 247771 506866 248091 506898
rect 262910 507454 263230 507486
rect 262910 507218 262952 507454
rect 263188 507218 263230 507454
rect 262910 507134 263230 507218
rect 262910 506898 262952 507134
rect 263188 506898 263230 507134
rect 262910 506866 263230 506898
rect 268840 507454 269160 507486
rect 268840 507218 268882 507454
rect 269118 507218 269160 507454
rect 268840 507134 269160 507218
rect 268840 506898 268882 507134
rect 269118 506898 269160 507134
rect 268840 506866 269160 506898
rect 274771 507454 275091 507486
rect 274771 507218 274813 507454
rect 275049 507218 275091 507454
rect 274771 507134 275091 507218
rect 274771 506898 274813 507134
rect 275049 506898 275091 507134
rect 274771 506866 275091 506898
rect 289910 507454 290230 507486
rect 289910 507218 289952 507454
rect 290188 507218 290230 507454
rect 289910 507134 290230 507218
rect 289910 506898 289952 507134
rect 290188 506898 290230 507134
rect 289910 506866 290230 506898
rect 295840 507454 296160 507486
rect 295840 507218 295882 507454
rect 296118 507218 296160 507454
rect 295840 507134 296160 507218
rect 295840 506898 295882 507134
rect 296118 506898 296160 507134
rect 295840 506866 296160 506898
rect 301771 507454 302091 507486
rect 301771 507218 301813 507454
rect 302049 507218 302091 507454
rect 301771 507134 302091 507218
rect 301771 506898 301813 507134
rect 302049 506898 302091 507134
rect 301771 506866 302091 506898
rect 316910 507454 317230 507486
rect 316910 507218 316952 507454
rect 317188 507218 317230 507454
rect 316910 507134 317230 507218
rect 316910 506898 316952 507134
rect 317188 506898 317230 507134
rect 316910 506866 317230 506898
rect 322840 507454 323160 507486
rect 322840 507218 322882 507454
rect 323118 507218 323160 507454
rect 322840 507134 323160 507218
rect 322840 506898 322882 507134
rect 323118 506898 323160 507134
rect 322840 506866 323160 506898
rect 328771 507454 329091 507486
rect 328771 507218 328813 507454
rect 329049 507218 329091 507454
rect 328771 507134 329091 507218
rect 328771 506898 328813 507134
rect 329049 506898 329091 507134
rect 328771 506866 329091 506898
rect 343910 507454 344230 507486
rect 343910 507218 343952 507454
rect 344188 507218 344230 507454
rect 343910 507134 344230 507218
rect 343910 506898 343952 507134
rect 344188 506898 344230 507134
rect 343910 506866 344230 506898
rect 349840 507454 350160 507486
rect 349840 507218 349882 507454
rect 350118 507218 350160 507454
rect 349840 507134 350160 507218
rect 349840 506898 349882 507134
rect 350118 506898 350160 507134
rect 349840 506866 350160 506898
rect 355771 507454 356091 507486
rect 355771 507218 355813 507454
rect 356049 507218 356091 507454
rect 355771 507134 356091 507218
rect 355771 506898 355813 507134
rect 356049 506898 356091 507134
rect 355771 506866 356091 506898
rect 370910 507454 371230 507486
rect 370910 507218 370952 507454
rect 371188 507218 371230 507454
rect 370910 507134 371230 507218
rect 370910 506898 370952 507134
rect 371188 506898 371230 507134
rect 370910 506866 371230 506898
rect 376840 507454 377160 507486
rect 376840 507218 376882 507454
rect 377118 507218 377160 507454
rect 376840 507134 377160 507218
rect 376840 506898 376882 507134
rect 377118 506898 377160 507134
rect 376840 506866 377160 506898
rect 382771 507454 383091 507486
rect 382771 507218 382813 507454
rect 383049 507218 383091 507454
rect 382771 507134 383091 507218
rect 382771 506898 382813 507134
rect 383049 506898 383091 507134
rect 382771 506866 383091 506898
rect 397910 507454 398230 507486
rect 397910 507218 397952 507454
rect 398188 507218 398230 507454
rect 397910 507134 398230 507218
rect 397910 506898 397952 507134
rect 398188 506898 398230 507134
rect 397910 506866 398230 506898
rect 403840 507454 404160 507486
rect 403840 507218 403882 507454
rect 404118 507218 404160 507454
rect 403840 507134 404160 507218
rect 403840 506898 403882 507134
rect 404118 506898 404160 507134
rect 403840 506866 404160 506898
rect 409771 507454 410091 507486
rect 409771 507218 409813 507454
rect 410049 507218 410091 507454
rect 409771 507134 410091 507218
rect 409771 506898 409813 507134
rect 410049 506898 410091 507134
rect 409771 506866 410091 506898
rect 424910 507454 425230 507486
rect 424910 507218 424952 507454
rect 425188 507218 425230 507454
rect 424910 507134 425230 507218
rect 424910 506898 424952 507134
rect 425188 506898 425230 507134
rect 424910 506866 425230 506898
rect 430840 507454 431160 507486
rect 430840 507218 430882 507454
rect 431118 507218 431160 507454
rect 430840 507134 431160 507218
rect 430840 506898 430882 507134
rect 431118 506898 431160 507134
rect 430840 506866 431160 506898
rect 436771 507454 437091 507486
rect 436771 507218 436813 507454
rect 437049 507218 437091 507454
rect 436771 507134 437091 507218
rect 436771 506898 436813 507134
rect 437049 506898 437091 507134
rect 436771 506866 437091 506898
rect 451910 507454 452230 507486
rect 451910 507218 451952 507454
rect 452188 507218 452230 507454
rect 451910 507134 452230 507218
rect 451910 506898 451952 507134
rect 452188 506898 452230 507134
rect 451910 506866 452230 506898
rect 457840 507454 458160 507486
rect 457840 507218 457882 507454
rect 458118 507218 458160 507454
rect 457840 507134 458160 507218
rect 457840 506898 457882 507134
rect 458118 506898 458160 507134
rect 457840 506866 458160 506898
rect 463771 507454 464091 507486
rect 463771 507218 463813 507454
rect 464049 507218 464091 507454
rect 463771 507134 464091 507218
rect 463771 506898 463813 507134
rect 464049 506898 464091 507134
rect 463771 506866 464091 506898
rect 478910 507454 479230 507486
rect 478910 507218 478952 507454
rect 479188 507218 479230 507454
rect 478910 507134 479230 507218
rect 478910 506898 478952 507134
rect 479188 506898 479230 507134
rect 478910 506866 479230 506898
rect 484840 507454 485160 507486
rect 484840 507218 484882 507454
rect 485118 507218 485160 507454
rect 484840 507134 485160 507218
rect 484840 506898 484882 507134
rect 485118 506898 485160 507134
rect 484840 506866 485160 506898
rect 490771 507454 491091 507486
rect 490771 507218 490813 507454
rect 491049 507218 491091 507454
rect 490771 507134 491091 507218
rect 490771 506898 490813 507134
rect 491049 506898 491091 507134
rect 490771 506866 491091 506898
rect 505910 507454 506230 507486
rect 505910 507218 505952 507454
rect 506188 507218 506230 507454
rect 505910 507134 506230 507218
rect 505910 506898 505952 507134
rect 506188 506898 506230 507134
rect 505910 506866 506230 506898
rect 511840 507454 512160 507486
rect 511840 507218 511882 507454
rect 512118 507218 512160 507454
rect 511840 507134 512160 507218
rect 511840 506898 511882 507134
rect 512118 506898 512160 507134
rect 511840 506866 512160 506898
rect 517771 507454 518091 507486
rect 517771 507218 517813 507454
rect 518049 507218 518091 507454
rect 517771 507134 518091 507218
rect 517771 506898 517813 507134
rect 518049 506898 518091 507134
rect 517771 506866 518091 506898
rect 532910 507454 533230 507486
rect 532910 507218 532952 507454
rect 533188 507218 533230 507454
rect 532910 507134 533230 507218
rect 532910 506898 532952 507134
rect 533188 506898 533230 507134
rect 532910 506866 533230 506898
rect 538840 507454 539160 507486
rect 538840 507218 538882 507454
rect 539118 507218 539160 507454
rect 538840 507134 539160 507218
rect 538840 506898 538882 507134
rect 539118 506898 539160 507134
rect 538840 506866 539160 506898
rect 544771 507454 545091 507486
rect 544771 507218 544813 507454
rect 545049 507218 545091 507454
rect 544771 507134 545091 507218
rect 544771 506898 544813 507134
rect 545049 506898 545091 507134
rect 544771 506866 545091 506898
rect 559794 507454 560414 524898
rect 559794 507218 559826 507454
rect 560062 507218 560146 507454
rect 560382 507218 560414 507454
rect 559794 507134 560414 507218
rect 559794 506898 559826 507134
rect 560062 506898 560146 507134
rect 560382 506898 560414 507134
rect 10794 498218 10826 498454
rect 11062 498218 11146 498454
rect 11382 498218 11414 498454
rect 10794 498134 11414 498218
rect 10794 497898 10826 498134
rect 11062 497898 11146 498134
rect 11382 497898 11414 498134
rect 10794 480454 11414 497898
rect 19794 499394 20414 500000
rect 19794 499158 19826 499394
rect 20062 499158 20146 499394
rect 20382 499158 20414 499394
rect 19794 499074 20414 499158
rect 19794 498838 19826 499074
rect 20062 498838 20146 499074
rect 20382 498838 20414 499074
rect 19794 497000 20414 498838
rect 28794 498454 29414 500000
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 497000 29414 497898
rect 37794 499394 38414 500000
rect 37794 499158 37826 499394
rect 38062 499158 38146 499394
rect 38382 499158 38414 499394
rect 37794 499074 38414 499158
rect 37794 498838 37826 499074
rect 38062 498838 38146 499074
rect 38382 498838 38414 499074
rect 37794 497000 38414 498838
rect 46794 498454 47414 500000
rect 46794 498218 46826 498454
rect 47062 498218 47146 498454
rect 47382 498218 47414 498454
rect 46794 498134 47414 498218
rect 46794 497898 46826 498134
rect 47062 497898 47146 498134
rect 47382 497898 47414 498134
rect 46794 497000 47414 497898
rect 55794 499394 56414 500000
rect 55794 499158 55826 499394
rect 56062 499158 56146 499394
rect 56382 499158 56414 499394
rect 55794 499074 56414 499158
rect 55794 498838 55826 499074
rect 56062 498838 56146 499074
rect 56382 498838 56414 499074
rect 55794 497000 56414 498838
rect 64794 498454 65414 500000
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 497000 65414 497898
rect 73794 499394 74414 500000
rect 73794 499158 73826 499394
rect 74062 499158 74146 499394
rect 74382 499158 74414 499394
rect 73794 499074 74414 499158
rect 73794 498838 73826 499074
rect 74062 498838 74146 499074
rect 74382 498838 74414 499074
rect 73794 497000 74414 498838
rect 82794 498454 83414 500000
rect 82794 498218 82826 498454
rect 83062 498218 83146 498454
rect 83382 498218 83414 498454
rect 82794 498134 83414 498218
rect 82794 497898 82826 498134
rect 83062 497898 83146 498134
rect 83382 497898 83414 498134
rect 82794 497000 83414 497898
rect 91794 499394 92414 500000
rect 91794 499158 91826 499394
rect 92062 499158 92146 499394
rect 92382 499158 92414 499394
rect 91794 499074 92414 499158
rect 91794 498838 91826 499074
rect 92062 498838 92146 499074
rect 92382 498838 92414 499074
rect 91794 497000 92414 498838
rect 100794 498454 101414 500000
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 497000 101414 497898
rect 109794 499394 110414 500000
rect 109794 499158 109826 499394
rect 110062 499158 110146 499394
rect 110382 499158 110414 499394
rect 109794 499074 110414 499158
rect 109794 498838 109826 499074
rect 110062 498838 110146 499074
rect 110382 498838 110414 499074
rect 109794 497000 110414 498838
rect 118794 498454 119414 500000
rect 118794 498218 118826 498454
rect 119062 498218 119146 498454
rect 119382 498218 119414 498454
rect 118794 498134 119414 498218
rect 118794 497898 118826 498134
rect 119062 497898 119146 498134
rect 119382 497898 119414 498134
rect 118794 497000 119414 497898
rect 127794 499394 128414 500000
rect 127794 499158 127826 499394
rect 128062 499158 128146 499394
rect 128382 499158 128414 499394
rect 127794 499074 128414 499158
rect 127794 498838 127826 499074
rect 128062 498838 128146 499074
rect 128382 498838 128414 499074
rect 127794 497000 128414 498838
rect 136794 498454 137414 500000
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 497000 137414 497898
rect 145794 499394 146414 500000
rect 145794 499158 145826 499394
rect 146062 499158 146146 499394
rect 146382 499158 146414 499394
rect 145794 499074 146414 499158
rect 145794 498838 145826 499074
rect 146062 498838 146146 499074
rect 146382 498838 146414 499074
rect 145794 497000 146414 498838
rect 154794 498454 155414 500000
rect 154794 498218 154826 498454
rect 155062 498218 155146 498454
rect 155382 498218 155414 498454
rect 154794 498134 155414 498218
rect 154794 497898 154826 498134
rect 155062 497898 155146 498134
rect 155382 497898 155414 498134
rect 154794 497000 155414 497898
rect 163794 499394 164414 500000
rect 163794 499158 163826 499394
rect 164062 499158 164146 499394
rect 164382 499158 164414 499394
rect 163794 499074 164414 499158
rect 163794 498838 163826 499074
rect 164062 498838 164146 499074
rect 164382 498838 164414 499074
rect 163794 497000 164414 498838
rect 172794 498454 173414 500000
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 497000 173414 497898
rect 181794 499394 182414 500000
rect 181794 499158 181826 499394
rect 182062 499158 182146 499394
rect 182382 499158 182414 499394
rect 181794 499074 182414 499158
rect 181794 498838 181826 499074
rect 182062 498838 182146 499074
rect 182382 498838 182414 499074
rect 181794 497000 182414 498838
rect 190794 498454 191414 500000
rect 190794 498218 190826 498454
rect 191062 498218 191146 498454
rect 191382 498218 191414 498454
rect 190794 498134 191414 498218
rect 190794 497898 190826 498134
rect 191062 497898 191146 498134
rect 191382 497898 191414 498134
rect 190794 497000 191414 497898
rect 199794 499394 200414 500000
rect 199794 499158 199826 499394
rect 200062 499158 200146 499394
rect 200382 499158 200414 499394
rect 199794 499074 200414 499158
rect 199794 498838 199826 499074
rect 200062 498838 200146 499074
rect 200382 498838 200414 499074
rect 199794 497000 200414 498838
rect 208794 498454 209414 500000
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 497000 209414 497898
rect 217794 499394 218414 500000
rect 217794 499158 217826 499394
rect 218062 499158 218146 499394
rect 218382 499158 218414 499394
rect 217794 499074 218414 499158
rect 217794 498838 217826 499074
rect 218062 498838 218146 499074
rect 218382 498838 218414 499074
rect 217794 497000 218414 498838
rect 226794 498454 227414 500000
rect 226794 498218 226826 498454
rect 227062 498218 227146 498454
rect 227382 498218 227414 498454
rect 226794 498134 227414 498218
rect 226794 497898 226826 498134
rect 227062 497898 227146 498134
rect 227382 497898 227414 498134
rect 226794 497000 227414 497898
rect 235794 499394 236414 500000
rect 235794 499158 235826 499394
rect 236062 499158 236146 499394
rect 236382 499158 236414 499394
rect 235794 499074 236414 499158
rect 235794 498838 235826 499074
rect 236062 498838 236146 499074
rect 236382 498838 236414 499074
rect 235794 497000 236414 498838
rect 244794 498454 245414 500000
rect 244794 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 245414 498454
rect 244794 498134 245414 498218
rect 244794 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 245414 498134
rect 244794 497000 245414 497898
rect 253794 499394 254414 500000
rect 253794 499158 253826 499394
rect 254062 499158 254146 499394
rect 254382 499158 254414 499394
rect 253794 499074 254414 499158
rect 253794 498838 253826 499074
rect 254062 498838 254146 499074
rect 254382 498838 254414 499074
rect 253794 497000 254414 498838
rect 262794 498454 263414 500000
rect 262794 498218 262826 498454
rect 263062 498218 263146 498454
rect 263382 498218 263414 498454
rect 262794 498134 263414 498218
rect 262794 497898 262826 498134
rect 263062 497898 263146 498134
rect 263382 497898 263414 498134
rect 262794 497000 263414 497898
rect 271794 499394 272414 500000
rect 271794 499158 271826 499394
rect 272062 499158 272146 499394
rect 272382 499158 272414 499394
rect 271794 499074 272414 499158
rect 271794 498838 271826 499074
rect 272062 498838 272146 499074
rect 272382 498838 272414 499074
rect 271794 497000 272414 498838
rect 280794 498454 281414 500000
rect 280794 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 281414 498454
rect 280794 498134 281414 498218
rect 280794 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 281414 498134
rect 280794 497000 281414 497898
rect 289794 499394 290414 500000
rect 289794 499158 289826 499394
rect 290062 499158 290146 499394
rect 290382 499158 290414 499394
rect 289794 499074 290414 499158
rect 289794 498838 289826 499074
rect 290062 498838 290146 499074
rect 290382 498838 290414 499074
rect 289794 497000 290414 498838
rect 298794 498454 299414 500000
rect 298794 498218 298826 498454
rect 299062 498218 299146 498454
rect 299382 498218 299414 498454
rect 298794 498134 299414 498218
rect 298794 497898 298826 498134
rect 299062 497898 299146 498134
rect 299382 497898 299414 498134
rect 298794 497000 299414 497898
rect 307794 499394 308414 500000
rect 307794 499158 307826 499394
rect 308062 499158 308146 499394
rect 308382 499158 308414 499394
rect 307794 499074 308414 499158
rect 307794 498838 307826 499074
rect 308062 498838 308146 499074
rect 308382 498838 308414 499074
rect 307794 497000 308414 498838
rect 316794 498454 317414 500000
rect 316794 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 317414 498454
rect 316794 498134 317414 498218
rect 316794 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 317414 498134
rect 316794 497000 317414 497898
rect 325794 499394 326414 500000
rect 325794 499158 325826 499394
rect 326062 499158 326146 499394
rect 326382 499158 326414 499394
rect 325794 499074 326414 499158
rect 325794 498838 325826 499074
rect 326062 498838 326146 499074
rect 326382 498838 326414 499074
rect 325794 497000 326414 498838
rect 334794 498454 335414 500000
rect 334794 498218 334826 498454
rect 335062 498218 335146 498454
rect 335382 498218 335414 498454
rect 334794 498134 335414 498218
rect 334794 497898 334826 498134
rect 335062 497898 335146 498134
rect 335382 497898 335414 498134
rect 334794 497000 335414 497898
rect 343794 499394 344414 500000
rect 343794 499158 343826 499394
rect 344062 499158 344146 499394
rect 344382 499158 344414 499394
rect 343794 499074 344414 499158
rect 343794 498838 343826 499074
rect 344062 498838 344146 499074
rect 344382 498838 344414 499074
rect 343794 497000 344414 498838
rect 352794 498454 353414 500000
rect 352794 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 353414 498454
rect 352794 498134 353414 498218
rect 352794 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 353414 498134
rect 352794 497000 353414 497898
rect 361794 499394 362414 500000
rect 361794 499158 361826 499394
rect 362062 499158 362146 499394
rect 362382 499158 362414 499394
rect 361794 499074 362414 499158
rect 361794 498838 361826 499074
rect 362062 498838 362146 499074
rect 362382 498838 362414 499074
rect 361794 497000 362414 498838
rect 370794 498454 371414 500000
rect 370794 498218 370826 498454
rect 371062 498218 371146 498454
rect 371382 498218 371414 498454
rect 370794 498134 371414 498218
rect 370794 497898 370826 498134
rect 371062 497898 371146 498134
rect 371382 497898 371414 498134
rect 370794 497000 371414 497898
rect 379794 499394 380414 500000
rect 379794 499158 379826 499394
rect 380062 499158 380146 499394
rect 380382 499158 380414 499394
rect 379794 499074 380414 499158
rect 379794 498838 379826 499074
rect 380062 498838 380146 499074
rect 380382 498838 380414 499074
rect 379794 497000 380414 498838
rect 388794 498454 389414 500000
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 497000 389414 497898
rect 397794 499394 398414 500000
rect 397794 499158 397826 499394
rect 398062 499158 398146 499394
rect 398382 499158 398414 499394
rect 397794 499074 398414 499158
rect 397794 498838 397826 499074
rect 398062 498838 398146 499074
rect 398382 498838 398414 499074
rect 397794 497000 398414 498838
rect 406794 498454 407414 500000
rect 406794 498218 406826 498454
rect 407062 498218 407146 498454
rect 407382 498218 407414 498454
rect 406794 498134 407414 498218
rect 406794 497898 406826 498134
rect 407062 497898 407146 498134
rect 407382 497898 407414 498134
rect 406794 497000 407414 497898
rect 415794 499394 416414 500000
rect 415794 499158 415826 499394
rect 416062 499158 416146 499394
rect 416382 499158 416414 499394
rect 415794 499074 416414 499158
rect 415794 498838 415826 499074
rect 416062 498838 416146 499074
rect 416382 498838 416414 499074
rect 415794 497000 416414 498838
rect 424794 498454 425414 500000
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 497000 425414 497898
rect 433794 499394 434414 500000
rect 433794 499158 433826 499394
rect 434062 499158 434146 499394
rect 434382 499158 434414 499394
rect 433794 499074 434414 499158
rect 433794 498838 433826 499074
rect 434062 498838 434146 499074
rect 434382 498838 434414 499074
rect 433794 497000 434414 498838
rect 442794 498454 443414 500000
rect 442794 498218 442826 498454
rect 443062 498218 443146 498454
rect 443382 498218 443414 498454
rect 442794 498134 443414 498218
rect 442794 497898 442826 498134
rect 443062 497898 443146 498134
rect 443382 497898 443414 498134
rect 442794 497000 443414 497898
rect 451794 499394 452414 500000
rect 451794 499158 451826 499394
rect 452062 499158 452146 499394
rect 452382 499158 452414 499394
rect 451794 499074 452414 499158
rect 451794 498838 451826 499074
rect 452062 498838 452146 499074
rect 452382 498838 452414 499074
rect 451794 497000 452414 498838
rect 460794 498454 461414 500000
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 497000 461414 497898
rect 469794 499394 470414 500000
rect 469794 499158 469826 499394
rect 470062 499158 470146 499394
rect 470382 499158 470414 499394
rect 469794 499074 470414 499158
rect 469794 498838 469826 499074
rect 470062 498838 470146 499074
rect 470382 498838 470414 499074
rect 469794 497000 470414 498838
rect 478794 498454 479414 500000
rect 478794 498218 478826 498454
rect 479062 498218 479146 498454
rect 479382 498218 479414 498454
rect 478794 498134 479414 498218
rect 478794 497898 478826 498134
rect 479062 497898 479146 498134
rect 479382 497898 479414 498134
rect 478794 497000 479414 497898
rect 487794 499394 488414 500000
rect 487794 499158 487826 499394
rect 488062 499158 488146 499394
rect 488382 499158 488414 499394
rect 487794 499074 488414 499158
rect 487794 498838 487826 499074
rect 488062 498838 488146 499074
rect 488382 498838 488414 499074
rect 487794 497000 488414 498838
rect 496794 498454 497414 500000
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 497000 497414 497898
rect 505794 499394 506414 500000
rect 505794 499158 505826 499394
rect 506062 499158 506146 499394
rect 506382 499158 506414 499394
rect 505794 499074 506414 499158
rect 505794 498838 505826 499074
rect 506062 498838 506146 499074
rect 506382 498838 506414 499074
rect 505794 497000 506414 498838
rect 514794 498454 515414 500000
rect 514794 498218 514826 498454
rect 515062 498218 515146 498454
rect 515382 498218 515414 498454
rect 514794 498134 515414 498218
rect 514794 497898 514826 498134
rect 515062 497898 515146 498134
rect 515382 497898 515414 498134
rect 514794 497000 515414 497898
rect 523794 499394 524414 500000
rect 523794 499158 523826 499394
rect 524062 499158 524146 499394
rect 524382 499158 524414 499394
rect 523794 499074 524414 499158
rect 523794 498838 523826 499074
rect 524062 498838 524146 499074
rect 524382 498838 524414 499074
rect 523794 497000 524414 498838
rect 532794 498454 533414 500000
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 497000 533414 497898
rect 541794 499394 542414 500000
rect 541794 499158 541826 499394
rect 542062 499158 542146 499394
rect 542382 499158 542414 499394
rect 541794 499074 542414 499158
rect 541794 498838 541826 499074
rect 542062 498838 542146 499074
rect 542382 498838 542414 499074
rect 541794 497000 542414 498838
rect 550794 498454 551414 500000
rect 550794 498218 550826 498454
rect 551062 498218 551146 498454
rect 551382 498218 551414 498454
rect 550794 498134 551414 498218
rect 550794 497898 550826 498134
rect 551062 497898 551146 498134
rect 551382 497898 551414 498134
rect 550794 497000 551414 497898
rect 19910 489454 20230 489486
rect 19910 489218 19952 489454
rect 20188 489218 20230 489454
rect 19910 489134 20230 489218
rect 19910 488898 19952 489134
rect 20188 488898 20230 489134
rect 19910 488866 20230 488898
rect 25840 489454 26160 489486
rect 25840 489218 25882 489454
rect 26118 489218 26160 489454
rect 25840 489134 26160 489218
rect 25840 488898 25882 489134
rect 26118 488898 26160 489134
rect 25840 488866 26160 488898
rect 31771 489454 32091 489486
rect 31771 489218 31813 489454
rect 32049 489218 32091 489454
rect 31771 489134 32091 489218
rect 31771 488898 31813 489134
rect 32049 488898 32091 489134
rect 31771 488866 32091 488898
rect 46910 489454 47230 489486
rect 46910 489218 46952 489454
rect 47188 489218 47230 489454
rect 46910 489134 47230 489218
rect 46910 488898 46952 489134
rect 47188 488898 47230 489134
rect 46910 488866 47230 488898
rect 52840 489454 53160 489486
rect 52840 489218 52882 489454
rect 53118 489218 53160 489454
rect 52840 489134 53160 489218
rect 52840 488898 52882 489134
rect 53118 488898 53160 489134
rect 52840 488866 53160 488898
rect 58771 489454 59091 489486
rect 58771 489218 58813 489454
rect 59049 489218 59091 489454
rect 58771 489134 59091 489218
rect 58771 488898 58813 489134
rect 59049 488898 59091 489134
rect 58771 488866 59091 488898
rect 73910 489454 74230 489486
rect 73910 489218 73952 489454
rect 74188 489218 74230 489454
rect 73910 489134 74230 489218
rect 73910 488898 73952 489134
rect 74188 488898 74230 489134
rect 73910 488866 74230 488898
rect 79840 489454 80160 489486
rect 79840 489218 79882 489454
rect 80118 489218 80160 489454
rect 79840 489134 80160 489218
rect 79840 488898 79882 489134
rect 80118 488898 80160 489134
rect 79840 488866 80160 488898
rect 85771 489454 86091 489486
rect 85771 489218 85813 489454
rect 86049 489218 86091 489454
rect 85771 489134 86091 489218
rect 85771 488898 85813 489134
rect 86049 488898 86091 489134
rect 85771 488866 86091 488898
rect 100910 489454 101230 489486
rect 100910 489218 100952 489454
rect 101188 489218 101230 489454
rect 100910 489134 101230 489218
rect 100910 488898 100952 489134
rect 101188 488898 101230 489134
rect 100910 488866 101230 488898
rect 106840 489454 107160 489486
rect 106840 489218 106882 489454
rect 107118 489218 107160 489454
rect 106840 489134 107160 489218
rect 106840 488898 106882 489134
rect 107118 488898 107160 489134
rect 106840 488866 107160 488898
rect 112771 489454 113091 489486
rect 112771 489218 112813 489454
rect 113049 489218 113091 489454
rect 112771 489134 113091 489218
rect 112771 488898 112813 489134
rect 113049 488898 113091 489134
rect 112771 488866 113091 488898
rect 127910 489454 128230 489486
rect 127910 489218 127952 489454
rect 128188 489218 128230 489454
rect 127910 489134 128230 489218
rect 127910 488898 127952 489134
rect 128188 488898 128230 489134
rect 127910 488866 128230 488898
rect 133840 489454 134160 489486
rect 133840 489218 133882 489454
rect 134118 489218 134160 489454
rect 133840 489134 134160 489218
rect 133840 488898 133882 489134
rect 134118 488898 134160 489134
rect 133840 488866 134160 488898
rect 139771 489454 140091 489486
rect 139771 489218 139813 489454
rect 140049 489218 140091 489454
rect 139771 489134 140091 489218
rect 139771 488898 139813 489134
rect 140049 488898 140091 489134
rect 139771 488866 140091 488898
rect 154910 489454 155230 489486
rect 154910 489218 154952 489454
rect 155188 489218 155230 489454
rect 154910 489134 155230 489218
rect 154910 488898 154952 489134
rect 155188 488898 155230 489134
rect 154910 488866 155230 488898
rect 160840 489454 161160 489486
rect 160840 489218 160882 489454
rect 161118 489218 161160 489454
rect 160840 489134 161160 489218
rect 160840 488898 160882 489134
rect 161118 488898 161160 489134
rect 160840 488866 161160 488898
rect 166771 489454 167091 489486
rect 166771 489218 166813 489454
rect 167049 489218 167091 489454
rect 166771 489134 167091 489218
rect 166771 488898 166813 489134
rect 167049 488898 167091 489134
rect 166771 488866 167091 488898
rect 181910 489454 182230 489486
rect 181910 489218 181952 489454
rect 182188 489218 182230 489454
rect 181910 489134 182230 489218
rect 181910 488898 181952 489134
rect 182188 488898 182230 489134
rect 181910 488866 182230 488898
rect 187840 489454 188160 489486
rect 187840 489218 187882 489454
rect 188118 489218 188160 489454
rect 187840 489134 188160 489218
rect 187840 488898 187882 489134
rect 188118 488898 188160 489134
rect 187840 488866 188160 488898
rect 193771 489454 194091 489486
rect 193771 489218 193813 489454
rect 194049 489218 194091 489454
rect 193771 489134 194091 489218
rect 193771 488898 193813 489134
rect 194049 488898 194091 489134
rect 193771 488866 194091 488898
rect 208910 489454 209230 489486
rect 208910 489218 208952 489454
rect 209188 489218 209230 489454
rect 208910 489134 209230 489218
rect 208910 488898 208952 489134
rect 209188 488898 209230 489134
rect 208910 488866 209230 488898
rect 214840 489454 215160 489486
rect 214840 489218 214882 489454
rect 215118 489218 215160 489454
rect 214840 489134 215160 489218
rect 214840 488898 214882 489134
rect 215118 488898 215160 489134
rect 214840 488866 215160 488898
rect 220771 489454 221091 489486
rect 220771 489218 220813 489454
rect 221049 489218 221091 489454
rect 220771 489134 221091 489218
rect 220771 488898 220813 489134
rect 221049 488898 221091 489134
rect 220771 488866 221091 488898
rect 235910 489454 236230 489486
rect 235910 489218 235952 489454
rect 236188 489218 236230 489454
rect 235910 489134 236230 489218
rect 235910 488898 235952 489134
rect 236188 488898 236230 489134
rect 235910 488866 236230 488898
rect 241840 489454 242160 489486
rect 241840 489218 241882 489454
rect 242118 489218 242160 489454
rect 241840 489134 242160 489218
rect 241840 488898 241882 489134
rect 242118 488898 242160 489134
rect 241840 488866 242160 488898
rect 247771 489454 248091 489486
rect 247771 489218 247813 489454
rect 248049 489218 248091 489454
rect 247771 489134 248091 489218
rect 247771 488898 247813 489134
rect 248049 488898 248091 489134
rect 247771 488866 248091 488898
rect 262910 489454 263230 489486
rect 262910 489218 262952 489454
rect 263188 489218 263230 489454
rect 262910 489134 263230 489218
rect 262910 488898 262952 489134
rect 263188 488898 263230 489134
rect 262910 488866 263230 488898
rect 268840 489454 269160 489486
rect 268840 489218 268882 489454
rect 269118 489218 269160 489454
rect 268840 489134 269160 489218
rect 268840 488898 268882 489134
rect 269118 488898 269160 489134
rect 268840 488866 269160 488898
rect 274771 489454 275091 489486
rect 274771 489218 274813 489454
rect 275049 489218 275091 489454
rect 274771 489134 275091 489218
rect 274771 488898 274813 489134
rect 275049 488898 275091 489134
rect 274771 488866 275091 488898
rect 289910 489454 290230 489486
rect 289910 489218 289952 489454
rect 290188 489218 290230 489454
rect 289910 489134 290230 489218
rect 289910 488898 289952 489134
rect 290188 488898 290230 489134
rect 289910 488866 290230 488898
rect 295840 489454 296160 489486
rect 295840 489218 295882 489454
rect 296118 489218 296160 489454
rect 295840 489134 296160 489218
rect 295840 488898 295882 489134
rect 296118 488898 296160 489134
rect 295840 488866 296160 488898
rect 301771 489454 302091 489486
rect 301771 489218 301813 489454
rect 302049 489218 302091 489454
rect 301771 489134 302091 489218
rect 301771 488898 301813 489134
rect 302049 488898 302091 489134
rect 301771 488866 302091 488898
rect 316910 489454 317230 489486
rect 316910 489218 316952 489454
rect 317188 489218 317230 489454
rect 316910 489134 317230 489218
rect 316910 488898 316952 489134
rect 317188 488898 317230 489134
rect 316910 488866 317230 488898
rect 322840 489454 323160 489486
rect 322840 489218 322882 489454
rect 323118 489218 323160 489454
rect 322840 489134 323160 489218
rect 322840 488898 322882 489134
rect 323118 488898 323160 489134
rect 322840 488866 323160 488898
rect 328771 489454 329091 489486
rect 328771 489218 328813 489454
rect 329049 489218 329091 489454
rect 328771 489134 329091 489218
rect 328771 488898 328813 489134
rect 329049 488898 329091 489134
rect 328771 488866 329091 488898
rect 343910 489454 344230 489486
rect 343910 489218 343952 489454
rect 344188 489218 344230 489454
rect 343910 489134 344230 489218
rect 343910 488898 343952 489134
rect 344188 488898 344230 489134
rect 343910 488866 344230 488898
rect 349840 489454 350160 489486
rect 349840 489218 349882 489454
rect 350118 489218 350160 489454
rect 349840 489134 350160 489218
rect 349840 488898 349882 489134
rect 350118 488898 350160 489134
rect 349840 488866 350160 488898
rect 355771 489454 356091 489486
rect 355771 489218 355813 489454
rect 356049 489218 356091 489454
rect 355771 489134 356091 489218
rect 355771 488898 355813 489134
rect 356049 488898 356091 489134
rect 355771 488866 356091 488898
rect 370910 489454 371230 489486
rect 370910 489218 370952 489454
rect 371188 489218 371230 489454
rect 370910 489134 371230 489218
rect 370910 488898 370952 489134
rect 371188 488898 371230 489134
rect 370910 488866 371230 488898
rect 376840 489454 377160 489486
rect 376840 489218 376882 489454
rect 377118 489218 377160 489454
rect 376840 489134 377160 489218
rect 376840 488898 376882 489134
rect 377118 488898 377160 489134
rect 376840 488866 377160 488898
rect 382771 489454 383091 489486
rect 382771 489218 382813 489454
rect 383049 489218 383091 489454
rect 382771 489134 383091 489218
rect 382771 488898 382813 489134
rect 383049 488898 383091 489134
rect 382771 488866 383091 488898
rect 397910 489454 398230 489486
rect 397910 489218 397952 489454
rect 398188 489218 398230 489454
rect 397910 489134 398230 489218
rect 397910 488898 397952 489134
rect 398188 488898 398230 489134
rect 397910 488866 398230 488898
rect 403840 489454 404160 489486
rect 403840 489218 403882 489454
rect 404118 489218 404160 489454
rect 403840 489134 404160 489218
rect 403840 488898 403882 489134
rect 404118 488898 404160 489134
rect 403840 488866 404160 488898
rect 409771 489454 410091 489486
rect 409771 489218 409813 489454
rect 410049 489218 410091 489454
rect 409771 489134 410091 489218
rect 409771 488898 409813 489134
rect 410049 488898 410091 489134
rect 409771 488866 410091 488898
rect 424910 489454 425230 489486
rect 424910 489218 424952 489454
rect 425188 489218 425230 489454
rect 424910 489134 425230 489218
rect 424910 488898 424952 489134
rect 425188 488898 425230 489134
rect 424910 488866 425230 488898
rect 430840 489454 431160 489486
rect 430840 489218 430882 489454
rect 431118 489218 431160 489454
rect 430840 489134 431160 489218
rect 430840 488898 430882 489134
rect 431118 488898 431160 489134
rect 430840 488866 431160 488898
rect 436771 489454 437091 489486
rect 436771 489218 436813 489454
rect 437049 489218 437091 489454
rect 436771 489134 437091 489218
rect 436771 488898 436813 489134
rect 437049 488898 437091 489134
rect 436771 488866 437091 488898
rect 451910 489454 452230 489486
rect 451910 489218 451952 489454
rect 452188 489218 452230 489454
rect 451910 489134 452230 489218
rect 451910 488898 451952 489134
rect 452188 488898 452230 489134
rect 451910 488866 452230 488898
rect 457840 489454 458160 489486
rect 457840 489218 457882 489454
rect 458118 489218 458160 489454
rect 457840 489134 458160 489218
rect 457840 488898 457882 489134
rect 458118 488898 458160 489134
rect 457840 488866 458160 488898
rect 463771 489454 464091 489486
rect 463771 489218 463813 489454
rect 464049 489218 464091 489454
rect 463771 489134 464091 489218
rect 463771 488898 463813 489134
rect 464049 488898 464091 489134
rect 463771 488866 464091 488898
rect 478910 489454 479230 489486
rect 478910 489218 478952 489454
rect 479188 489218 479230 489454
rect 478910 489134 479230 489218
rect 478910 488898 478952 489134
rect 479188 488898 479230 489134
rect 478910 488866 479230 488898
rect 484840 489454 485160 489486
rect 484840 489218 484882 489454
rect 485118 489218 485160 489454
rect 484840 489134 485160 489218
rect 484840 488898 484882 489134
rect 485118 488898 485160 489134
rect 484840 488866 485160 488898
rect 490771 489454 491091 489486
rect 490771 489218 490813 489454
rect 491049 489218 491091 489454
rect 490771 489134 491091 489218
rect 490771 488898 490813 489134
rect 491049 488898 491091 489134
rect 490771 488866 491091 488898
rect 505910 489454 506230 489486
rect 505910 489218 505952 489454
rect 506188 489218 506230 489454
rect 505910 489134 506230 489218
rect 505910 488898 505952 489134
rect 506188 488898 506230 489134
rect 505910 488866 506230 488898
rect 511840 489454 512160 489486
rect 511840 489218 511882 489454
rect 512118 489218 512160 489454
rect 511840 489134 512160 489218
rect 511840 488898 511882 489134
rect 512118 488898 512160 489134
rect 511840 488866 512160 488898
rect 517771 489454 518091 489486
rect 517771 489218 517813 489454
rect 518049 489218 518091 489454
rect 517771 489134 518091 489218
rect 517771 488898 517813 489134
rect 518049 488898 518091 489134
rect 517771 488866 518091 488898
rect 532910 489454 533230 489486
rect 532910 489218 532952 489454
rect 533188 489218 533230 489454
rect 532910 489134 533230 489218
rect 532910 488898 532952 489134
rect 533188 488898 533230 489134
rect 532910 488866 533230 488898
rect 538840 489454 539160 489486
rect 538840 489218 538882 489454
rect 539118 489218 539160 489454
rect 538840 489134 539160 489218
rect 538840 488898 538882 489134
rect 539118 488898 539160 489134
rect 538840 488866 539160 488898
rect 544771 489454 545091 489486
rect 544771 489218 544813 489454
rect 545049 489218 545091 489454
rect 544771 489134 545091 489218
rect 544771 488898 544813 489134
rect 545049 488898 545091 489134
rect 544771 488866 545091 488898
rect 559794 489454 560414 506898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 462454 11414 479898
rect 22874 480454 23194 480486
rect 22874 480218 22916 480454
rect 23152 480218 23194 480454
rect 22874 480134 23194 480218
rect 22874 479898 22916 480134
rect 23152 479898 23194 480134
rect 22874 479866 23194 479898
rect 28805 480454 29125 480486
rect 28805 480218 28847 480454
rect 29083 480218 29125 480454
rect 28805 480134 29125 480218
rect 28805 479898 28847 480134
rect 29083 479898 29125 480134
rect 28805 479866 29125 479898
rect 49874 480454 50194 480486
rect 49874 480218 49916 480454
rect 50152 480218 50194 480454
rect 49874 480134 50194 480218
rect 49874 479898 49916 480134
rect 50152 479898 50194 480134
rect 49874 479866 50194 479898
rect 55805 480454 56125 480486
rect 55805 480218 55847 480454
rect 56083 480218 56125 480454
rect 55805 480134 56125 480218
rect 55805 479898 55847 480134
rect 56083 479898 56125 480134
rect 55805 479866 56125 479898
rect 76874 480454 77194 480486
rect 76874 480218 76916 480454
rect 77152 480218 77194 480454
rect 76874 480134 77194 480218
rect 76874 479898 76916 480134
rect 77152 479898 77194 480134
rect 76874 479866 77194 479898
rect 82805 480454 83125 480486
rect 82805 480218 82847 480454
rect 83083 480218 83125 480454
rect 82805 480134 83125 480218
rect 82805 479898 82847 480134
rect 83083 479898 83125 480134
rect 82805 479866 83125 479898
rect 103874 480454 104194 480486
rect 103874 480218 103916 480454
rect 104152 480218 104194 480454
rect 103874 480134 104194 480218
rect 103874 479898 103916 480134
rect 104152 479898 104194 480134
rect 103874 479866 104194 479898
rect 109805 480454 110125 480486
rect 109805 480218 109847 480454
rect 110083 480218 110125 480454
rect 109805 480134 110125 480218
rect 109805 479898 109847 480134
rect 110083 479898 110125 480134
rect 109805 479866 110125 479898
rect 130874 480454 131194 480486
rect 130874 480218 130916 480454
rect 131152 480218 131194 480454
rect 130874 480134 131194 480218
rect 130874 479898 130916 480134
rect 131152 479898 131194 480134
rect 130874 479866 131194 479898
rect 136805 480454 137125 480486
rect 136805 480218 136847 480454
rect 137083 480218 137125 480454
rect 136805 480134 137125 480218
rect 136805 479898 136847 480134
rect 137083 479898 137125 480134
rect 136805 479866 137125 479898
rect 157874 480454 158194 480486
rect 157874 480218 157916 480454
rect 158152 480218 158194 480454
rect 157874 480134 158194 480218
rect 157874 479898 157916 480134
rect 158152 479898 158194 480134
rect 157874 479866 158194 479898
rect 163805 480454 164125 480486
rect 163805 480218 163847 480454
rect 164083 480218 164125 480454
rect 163805 480134 164125 480218
rect 163805 479898 163847 480134
rect 164083 479898 164125 480134
rect 163805 479866 164125 479898
rect 184874 480454 185194 480486
rect 184874 480218 184916 480454
rect 185152 480218 185194 480454
rect 184874 480134 185194 480218
rect 184874 479898 184916 480134
rect 185152 479898 185194 480134
rect 184874 479866 185194 479898
rect 190805 480454 191125 480486
rect 190805 480218 190847 480454
rect 191083 480218 191125 480454
rect 190805 480134 191125 480218
rect 190805 479898 190847 480134
rect 191083 479898 191125 480134
rect 190805 479866 191125 479898
rect 211874 480454 212194 480486
rect 211874 480218 211916 480454
rect 212152 480218 212194 480454
rect 211874 480134 212194 480218
rect 211874 479898 211916 480134
rect 212152 479898 212194 480134
rect 211874 479866 212194 479898
rect 217805 480454 218125 480486
rect 217805 480218 217847 480454
rect 218083 480218 218125 480454
rect 217805 480134 218125 480218
rect 217805 479898 217847 480134
rect 218083 479898 218125 480134
rect 217805 479866 218125 479898
rect 238874 480454 239194 480486
rect 238874 480218 238916 480454
rect 239152 480218 239194 480454
rect 238874 480134 239194 480218
rect 238874 479898 238916 480134
rect 239152 479898 239194 480134
rect 238874 479866 239194 479898
rect 244805 480454 245125 480486
rect 244805 480218 244847 480454
rect 245083 480218 245125 480454
rect 244805 480134 245125 480218
rect 244805 479898 244847 480134
rect 245083 479898 245125 480134
rect 244805 479866 245125 479898
rect 265874 480454 266194 480486
rect 265874 480218 265916 480454
rect 266152 480218 266194 480454
rect 265874 480134 266194 480218
rect 265874 479898 265916 480134
rect 266152 479898 266194 480134
rect 265874 479866 266194 479898
rect 271805 480454 272125 480486
rect 271805 480218 271847 480454
rect 272083 480218 272125 480454
rect 271805 480134 272125 480218
rect 271805 479898 271847 480134
rect 272083 479898 272125 480134
rect 271805 479866 272125 479898
rect 292874 480454 293194 480486
rect 292874 480218 292916 480454
rect 293152 480218 293194 480454
rect 292874 480134 293194 480218
rect 292874 479898 292916 480134
rect 293152 479898 293194 480134
rect 292874 479866 293194 479898
rect 298805 480454 299125 480486
rect 298805 480218 298847 480454
rect 299083 480218 299125 480454
rect 298805 480134 299125 480218
rect 298805 479898 298847 480134
rect 299083 479898 299125 480134
rect 298805 479866 299125 479898
rect 319874 480454 320194 480486
rect 319874 480218 319916 480454
rect 320152 480218 320194 480454
rect 319874 480134 320194 480218
rect 319874 479898 319916 480134
rect 320152 479898 320194 480134
rect 319874 479866 320194 479898
rect 325805 480454 326125 480486
rect 325805 480218 325847 480454
rect 326083 480218 326125 480454
rect 325805 480134 326125 480218
rect 325805 479898 325847 480134
rect 326083 479898 326125 480134
rect 325805 479866 326125 479898
rect 346874 480454 347194 480486
rect 346874 480218 346916 480454
rect 347152 480218 347194 480454
rect 346874 480134 347194 480218
rect 346874 479898 346916 480134
rect 347152 479898 347194 480134
rect 346874 479866 347194 479898
rect 352805 480454 353125 480486
rect 352805 480218 352847 480454
rect 353083 480218 353125 480454
rect 352805 480134 353125 480218
rect 352805 479898 352847 480134
rect 353083 479898 353125 480134
rect 352805 479866 353125 479898
rect 373874 480454 374194 480486
rect 373874 480218 373916 480454
rect 374152 480218 374194 480454
rect 373874 480134 374194 480218
rect 373874 479898 373916 480134
rect 374152 479898 374194 480134
rect 373874 479866 374194 479898
rect 379805 480454 380125 480486
rect 379805 480218 379847 480454
rect 380083 480218 380125 480454
rect 379805 480134 380125 480218
rect 379805 479898 379847 480134
rect 380083 479898 380125 480134
rect 379805 479866 380125 479898
rect 400874 480454 401194 480486
rect 400874 480218 400916 480454
rect 401152 480218 401194 480454
rect 400874 480134 401194 480218
rect 400874 479898 400916 480134
rect 401152 479898 401194 480134
rect 400874 479866 401194 479898
rect 406805 480454 407125 480486
rect 406805 480218 406847 480454
rect 407083 480218 407125 480454
rect 406805 480134 407125 480218
rect 406805 479898 406847 480134
rect 407083 479898 407125 480134
rect 406805 479866 407125 479898
rect 427874 480454 428194 480486
rect 427874 480218 427916 480454
rect 428152 480218 428194 480454
rect 427874 480134 428194 480218
rect 427874 479898 427916 480134
rect 428152 479898 428194 480134
rect 427874 479866 428194 479898
rect 433805 480454 434125 480486
rect 433805 480218 433847 480454
rect 434083 480218 434125 480454
rect 433805 480134 434125 480218
rect 433805 479898 433847 480134
rect 434083 479898 434125 480134
rect 433805 479866 434125 479898
rect 454874 480454 455194 480486
rect 454874 480218 454916 480454
rect 455152 480218 455194 480454
rect 454874 480134 455194 480218
rect 454874 479898 454916 480134
rect 455152 479898 455194 480134
rect 454874 479866 455194 479898
rect 460805 480454 461125 480486
rect 460805 480218 460847 480454
rect 461083 480218 461125 480454
rect 460805 480134 461125 480218
rect 460805 479898 460847 480134
rect 461083 479898 461125 480134
rect 460805 479866 461125 479898
rect 481874 480454 482194 480486
rect 481874 480218 481916 480454
rect 482152 480218 482194 480454
rect 481874 480134 482194 480218
rect 481874 479898 481916 480134
rect 482152 479898 482194 480134
rect 481874 479866 482194 479898
rect 487805 480454 488125 480486
rect 487805 480218 487847 480454
rect 488083 480218 488125 480454
rect 487805 480134 488125 480218
rect 487805 479898 487847 480134
rect 488083 479898 488125 480134
rect 487805 479866 488125 479898
rect 508874 480454 509194 480486
rect 508874 480218 508916 480454
rect 509152 480218 509194 480454
rect 508874 480134 509194 480218
rect 508874 479898 508916 480134
rect 509152 479898 509194 480134
rect 508874 479866 509194 479898
rect 514805 480454 515125 480486
rect 514805 480218 514847 480454
rect 515083 480218 515125 480454
rect 514805 480134 515125 480218
rect 514805 479898 514847 480134
rect 515083 479898 515125 480134
rect 514805 479866 515125 479898
rect 535874 480454 536194 480486
rect 535874 480218 535916 480454
rect 536152 480218 536194 480454
rect 535874 480134 536194 480218
rect 535874 479898 535916 480134
rect 536152 479898 536194 480134
rect 535874 479866 536194 479898
rect 541805 480454 542125 480486
rect 541805 480218 541847 480454
rect 542083 480218 542125 480454
rect 541805 480134 542125 480218
rect 541805 479898 541847 480134
rect 542083 479898 542125 480134
rect 541805 479866 542125 479898
rect 19794 471454 20414 473000
rect 19794 471218 19826 471454
rect 20062 471218 20146 471454
rect 20382 471218 20414 471454
rect 19794 471134 20414 471218
rect 19794 470898 19826 471134
rect 20062 470898 20146 471134
rect 20382 470898 20414 471134
rect 19794 470000 20414 470898
rect 28794 472394 29414 473000
rect 28794 472158 28826 472394
rect 29062 472158 29146 472394
rect 29382 472158 29414 472394
rect 28794 472074 29414 472158
rect 28794 471838 28826 472074
rect 29062 471838 29146 472074
rect 29382 471838 29414 472074
rect 28794 470000 29414 471838
rect 37794 471454 38414 473000
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 470000 38414 470898
rect 46794 472394 47414 473000
rect 46794 472158 46826 472394
rect 47062 472158 47146 472394
rect 47382 472158 47414 472394
rect 46794 472074 47414 472158
rect 46794 471838 46826 472074
rect 47062 471838 47146 472074
rect 47382 471838 47414 472074
rect 46794 470000 47414 471838
rect 55794 471454 56414 473000
rect 55794 471218 55826 471454
rect 56062 471218 56146 471454
rect 56382 471218 56414 471454
rect 55794 471134 56414 471218
rect 55794 470898 55826 471134
rect 56062 470898 56146 471134
rect 56382 470898 56414 471134
rect 55794 470000 56414 470898
rect 64794 472394 65414 473000
rect 64794 472158 64826 472394
rect 65062 472158 65146 472394
rect 65382 472158 65414 472394
rect 64794 472074 65414 472158
rect 64794 471838 64826 472074
rect 65062 471838 65146 472074
rect 65382 471838 65414 472074
rect 64794 470000 65414 471838
rect 73794 471454 74414 473000
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 470000 74414 470898
rect 82794 472394 83414 473000
rect 82794 472158 82826 472394
rect 83062 472158 83146 472394
rect 83382 472158 83414 472394
rect 82794 472074 83414 472158
rect 82794 471838 82826 472074
rect 83062 471838 83146 472074
rect 83382 471838 83414 472074
rect 82794 470000 83414 471838
rect 91794 471454 92414 473000
rect 91794 471218 91826 471454
rect 92062 471218 92146 471454
rect 92382 471218 92414 471454
rect 91794 471134 92414 471218
rect 91794 470898 91826 471134
rect 92062 470898 92146 471134
rect 92382 470898 92414 471134
rect 91794 470000 92414 470898
rect 100794 472394 101414 473000
rect 100794 472158 100826 472394
rect 101062 472158 101146 472394
rect 101382 472158 101414 472394
rect 100794 472074 101414 472158
rect 100794 471838 100826 472074
rect 101062 471838 101146 472074
rect 101382 471838 101414 472074
rect 100794 470000 101414 471838
rect 109794 471454 110414 473000
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 470000 110414 470898
rect 118794 472394 119414 473000
rect 118794 472158 118826 472394
rect 119062 472158 119146 472394
rect 119382 472158 119414 472394
rect 118794 472074 119414 472158
rect 118794 471838 118826 472074
rect 119062 471838 119146 472074
rect 119382 471838 119414 472074
rect 118794 470000 119414 471838
rect 127794 471454 128414 473000
rect 127794 471218 127826 471454
rect 128062 471218 128146 471454
rect 128382 471218 128414 471454
rect 127794 471134 128414 471218
rect 127794 470898 127826 471134
rect 128062 470898 128146 471134
rect 128382 470898 128414 471134
rect 127794 470000 128414 470898
rect 136794 472394 137414 473000
rect 136794 472158 136826 472394
rect 137062 472158 137146 472394
rect 137382 472158 137414 472394
rect 136794 472074 137414 472158
rect 136794 471838 136826 472074
rect 137062 471838 137146 472074
rect 137382 471838 137414 472074
rect 136794 470000 137414 471838
rect 145794 471454 146414 473000
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 470000 146414 470898
rect 154794 472394 155414 473000
rect 154794 472158 154826 472394
rect 155062 472158 155146 472394
rect 155382 472158 155414 472394
rect 154794 472074 155414 472158
rect 154794 471838 154826 472074
rect 155062 471838 155146 472074
rect 155382 471838 155414 472074
rect 154794 470000 155414 471838
rect 163794 471454 164414 473000
rect 163794 471218 163826 471454
rect 164062 471218 164146 471454
rect 164382 471218 164414 471454
rect 163794 471134 164414 471218
rect 163794 470898 163826 471134
rect 164062 470898 164146 471134
rect 164382 470898 164414 471134
rect 163794 470000 164414 470898
rect 172794 472394 173414 473000
rect 172794 472158 172826 472394
rect 173062 472158 173146 472394
rect 173382 472158 173414 472394
rect 172794 472074 173414 472158
rect 172794 471838 172826 472074
rect 173062 471838 173146 472074
rect 173382 471838 173414 472074
rect 172794 470000 173414 471838
rect 181794 471454 182414 473000
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 470000 182414 470898
rect 190794 472394 191414 473000
rect 190794 472158 190826 472394
rect 191062 472158 191146 472394
rect 191382 472158 191414 472394
rect 190794 472074 191414 472158
rect 190794 471838 190826 472074
rect 191062 471838 191146 472074
rect 191382 471838 191414 472074
rect 190794 470000 191414 471838
rect 199794 471454 200414 473000
rect 199794 471218 199826 471454
rect 200062 471218 200146 471454
rect 200382 471218 200414 471454
rect 199794 471134 200414 471218
rect 199794 470898 199826 471134
rect 200062 470898 200146 471134
rect 200382 470898 200414 471134
rect 199794 470000 200414 470898
rect 208794 472394 209414 473000
rect 208794 472158 208826 472394
rect 209062 472158 209146 472394
rect 209382 472158 209414 472394
rect 208794 472074 209414 472158
rect 208794 471838 208826 472074
rect 209062 471838 209146 472074
rect 209382 471838 209414 472074
rect 208794 470000 209414 471838
rect 217794 471454 218414 473000
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 470000 218414 470898
rect 226794 472394 227414 473000
rect 226794 472158 226826 472394
rect 227062 472158 227146 472394
rect 227382 472158 227414 472394
rect 226794 472074 227414 472158
rect 226794 471838 226826 472074
rect 227062 471838 227146 472074
rect 227382 471838 227414 472074
rect 226794 470000 227414 471838
rect 235794 471454 236414 473000
rect 235794 471218 235826 471454
rect 236062 471218 236146 471454
rect 236382 471218 236414 471454
rect 235794 471134 236414 471218
rect 235794 470898 235826 471134
rect 236062 470898 236146 471134
rect 236382 470898 236414 471134
rect 235794 470000 236414 470898
rect 244794 472394 245414 473000
rect 244794 472158 244826 472394
rect 245062 472158 245146 472394
rect 245382 472158 245414 472394
rect 244794 472074 245414 472158
rect 244794 471838 244826 472074
rect 245062 471838 245146 472074
rect 245382 471838 245414 472074
rect 244794 470000 245414 471838
rect 253794 471454 254414 473000
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 470000 254414 470898
rect 262794 472394 263414 473000
rect 262794 472158 262826 472394
rect 263062 472158 263146 472394
rect 263382 472158 263414 472394
rect 262794 472074 263414 472158
rect 262794 471838 262826 472074
rect 263062 471838 263146 472074
rect 263382 471838 263414 472074
rect 262794 470000 263414 471838
rect 271794 471454 272414 473000
rect 271794 471218 271826 471454
rect 272062 471218 272146 471454
rect 272382 471218 272414 471454
rect 271794 471134 272414 471218
rect 271794 470898 271826 471134
rect 272062 470898 272146 471134
rect 272382 470898 272414 471134
rect 271794 470000 272414 470898
rect 280794 472394 281414 473000
rect 280794 472158 280826 472394
rect 281062 472158 281146 472394
rect 281382 472158 281414 472394
rect 280794 472074 281414 472158
rect 280794 471838 280826 472074
rect 281062 471838 281146 472074
rect 281382 471838 281414 472074
rect 280794 470000 281414 471838
rect 289794 471454 290414 473000
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 470000 290414 470898
rect 298794 472394 299414 473000
rect 298794 472158 298826 472394
rect 299062 472158 299146 472394
rect 299382 472158 299414 472394
rect 298794 472074 299414 472158
rect 298794 471838 298826 472074
rect 299062 471838 299146 472074
rect 299382 471838 299414 472074
rect 298794 470000 299414 471838
rect 307794 471454 308414 473000
rect 307794 471218 307826 471454
rect 308062 471218 308146 471454
rect 308382 471218 308414 471454
rect 307794 471134 308414 471218
rect 307794 470898 307826 471134
rect 308062 470898 308146 471134
rect 308382 470898 308414 471134
rect 307794 470000 308414 470898
rect 316794 472394 317414 473000
rect 316794 472158 316826 472394
rect 317062 472158 317146 472394
rect 317382 472158 317414 472394
rect 316794 472074 317414 472158
rect 316794 471838 316826 472074
rect 317062 471838 317146 472074
rect 317382 471838 317414 472074
rect 316794 470000 317414 471838
rect 325794 471454 326414 473000
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 470000 326414 470898
rect 334794 472394 335414 473000
rect 334794 472158 334826 472394
rect 335062 472158 335146 472394
rect 335382 472158 335414 472394
rect 334794 472074 335414 472158
rect 334794 471838 334826 472074
rect 335062 471838 335146 472074
rect 335382 471838 335414 472074
rect 334794 470000 335414 471838
rect 343794 471454 344414 473000
rect 343794 471218 343826 471454
rect 344062 471218 344146 471454
rect 344382 471218 344414 471454
rect 343794 471134 344414 471218
rect 343794 470898 343826 471134
rect 344062 470898 344146 471134
rect 344382 470898 344414 471134
rect 343794 470000 344414 470898
rect 352794 472394 353414 473000
rect 352794 472158 352826 472394
rect 353062 472158 353146 472394
rect 353382 472158 353414 472394
rect 352794 472074 353414 472158
rect 352794 471838 352826 472074
rect 353062 471838 353146 472074
rect 353382 471838 353414 472074
rect 352794 470000 353414 471838
rect 361794 471454 362414 473000
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 470000 362414 470898
rect 370794 472394 371414 473000
rect 370794 472158 370826 472394
rect 371062 472158 371146 472394
rect 371382 472158 371414 472394
rect 370794 472074 371414 472158
rect 370794 471838 370826 472074
rect 371062 471838 371146 472074
rect 371382 471838 371414 472074
rect 370794 470000 371414 471838
rect 379794 471454 380414 473000
rect 379794 471218 379826 471454
rect 380062 471218 380146 471454
rect 380382 471218 380414 471454
rect 379794 471134 380414 471218
rect 379794 470898 379826 471134
rect 380062 470898 380146 471134
rect 380382 470898 380414 471134
rect 379794 470000 380414 470898
rect 388794 472394 389414 473000
rect 388794 472158 388826 472394
rect 389062 472158 389146 472394
rect 389382 472158 389414 472394
rect 388794 472074 389414 472158
rect 388794 471838 388826 472074
rect 389062 471838 389146 472074
rect 389382 471838 389414 472074
rect 388794 470000 389414 471838
rect 397794 471454 398414 473000
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 470000 398414 470898
rect 406794 472394 407414 473000
rect 406794 472158 406826 472394
rect 407062 472158 407146 472394
rect 407382 472158 407414 472394
rect 406794 472074 407414 472158
rect 406794 471838 406826 472074
rect 407062 471838 407146 472074
rect 407382 471838 407414 472074
rect 406794 470000 407414 471838
rect 415794 471454 416414 473000
rect 415794 471218 415826 471454
rect 416062 471218 416146 471454
rect 416382 471218 416414 471454
rect 415794 471134 416414 471218
rect 415794 470898 415826 471134
rect 416062 470898 416146 471134
rect 416382 470898 416414 471134
rect 415794 470000 416414 470898
rect 424794 472394 425414 473000
rect 424794 472158 424826 472394
rect 425062 472158 425146 472394
rect 425382 472158 425414 472394
rect 424794 472074 425414 472158
rect 424794 471838 424826 472074
rect 425062 471838 425146 472074
rect 425382 471838 425414 472074
rect 424794 470000 425414 471838
rect 433794 471454 434414 473000
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 470000 434414 470898
rect 442794 472394 443414 473000
rect 442794 472158 442826 472394
rect 443062 472158 443146 472394
rect 443382 472158 443414 472394
rect 442794 472074 443414 472158
rect 442794 471838 442826 472074
rect 443062 471838 443146 472074
rect 443382 471838 443414 472074
rect 442794 470000 443414 471838
rect 451794 471454 452414 473000
rect 451794 471218 451826 471454
rect 452062 471218 452146 471454
rect 452382 471218 452414 471454
rect 451794 471134 452414 471218
rect 451794 470898 451826 471134
rect 452062 470898 452146 471134
rect 452382 470898 452414 471134
rect 451794 470000 452414 470898
rect 460794 472394 461414 473000
rect 460794 472158 460826 472394
rect 461062 472158 461146 472394
rect 461382 472158 461414 472394
rect 460794 472074 461414 472158
rect 460794 471838 460826 472074
rect 461062 471838 461146 472074
rect 461382 471838 461414 472074
rect 460794 470000 461414 471838
rect 469794 471454 470414 473000
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 470000 470414 470898
rect 478794 472394 479414 473000
rect 478794 472158 478826 472394
rect 479062 472158 479146 472394
rect 479382 472158 479414 472394
rect 478794 472074 479414 472158
rect 478794 471838 478826 472074
rect 479062 471838 479146 472074
rect 479382 471838 479414 472074
rect 478794 470000 479414 471838
rect 487794 471454 488414 473000
rect 487794 471218 487826 471454
rect 488062 471218 488146 471454
rect 488382 471218 488414 471454
rect 487794 471134 488414 471218
rect 487794 470898 487826 471134
rect 488062 470898 488146 471134
rect 488382 470898 488414 471134
rect 487794 470000 488414 470898
rect 496794 472394 497414 473000
rect 496794 472158 496826 472394
rect 497062 472158 497146 472394
rect 497382 472158 497414 472394
rect 496794 472074 497414 472158
rect 496794 471838 496826 472074
rect 497062 471838 497146 472074
rect 497382 471838 497414 472074
rect 496794 470000 497414 471838
rect 505794 471454 506414 473000
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 470000 506414 470898
rect 514794 472394 515414 473000
rect 514794 472158 514826 472394
rect 515062 472158 515146 472394
rect 515382 472158 515414 472394
rect 514794 472074 515414 472158
rect 514794 471838 514826 472074
rect 515062 471838 515146 472074
rect 515382 471838 515414 472074
rect 514794 470000 515414 471838
rect 523794 471454 524414 473000
rect 523794 471218 523826 471454
rect 524062 471218 524146 471454
rect 524382 471218 524414 471454
rect 523794 471134 524414 471218
rect 523794 470898 523826 471134
rect 524062 470898 524146 471134
rect 524382 470898 524414 471134
rect 523794 470000 524414 470898
rect 532794 472394 533414 473000
rect 532794 472158 532826 472394
rect 533062 472158 533146 472394
rect 533382 472158 533414 472394
rect 532794 472074 533414 472158
rect 532794 471838 532826 472074
rect 533062 471838 533146 472074
rect 533382 471838 533414 472074
rect 532794 470000 533414 471838
rect 541794 471454 542414 473000
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 470000 542414 470898
rect 550794 472394 551414 473000
rect 550794 472158 550826 472394
rect 551062 472158 551146 472394
rect 551382 472158 551414 472394
rect 550794 472074 551414 472158
rect 550794 471838 550826 472074
rect 551062 471838 551146 472074
rect 551382 471838 551414 472074
rect 550794 470000 551414 471838
rect 559794 471454 560414 488898
rect 559794 471218 559826 471454
rect 560062 471218 560146 471454
rect 560382 471218 560414 471454
rect 559794 471134 560414 471218
rect 559794 470898 559826 471134
rect 560062 470898 560146 471134
rect 560382 470898 560414 471134
rect 10794 462218 10826 462454
rect 11062 462218 11146 462454
rect 11382 462218 11414 462454
rect 10794 462134 11414 462218
rect 10794 461898 10826 462134
rect 11062 461898 11146 462134
rect 11382 461898 11414 462134
rect 10794 444454 11414 461898
rect 22874 462454 23194 462486
rect 22874 462218 22916 462454
rect 23152 462218 23194 462454
rect 22874 462134 23194 462218
rect 22874 461898 22916 462134
rect 23152 461898 23194 462134
rect 22874 461866 23194 461898
rect 28805 462454 29125 462486
rect 28805 462218 28847 462454
rect 29083 462218 29125 462454
rect 28805 462134 29125 462218
rect 28805 461898 28847 462134
rect 29083 461898 29125 462134
rect 28805 461866 29125 461898
rect 49874 462454 50194 462486
rect 49874 462218 49916 462454
rect 50152 462218 50194 462454
rect 49874 462134 50194 462218
rect 49874 461898 49916 462134
rect 50152 461898 50194 462134
rect 49874 461866 50194 461898
rect 55805 462454 56125 462486
rect 55805 462218 55847 462454
rect 56083 462218 56125 462454
rect 55805 462134 56125 462218
rect 55805 461898 55847 462134
rect 56083 461898 56125 462134
rect 55805 461866 56125 461898
rect 76874 462454 77194 462486
rect 76874 462218 76916 462454
rect 77152 462218 77194 462454
rect 76874 462134 77194 462218
rect 76874 461898 76916 462134
rect 77152 461898 77194 462134
rect 76874 461866 77194 461898
rect 82805 462454 83125 462486
rect 82805 462218 82847 462454
rect 83083 462218 83125 462454
rect 82805 462134 83125 462218
rect 82805 461898 82847 462134
rect 83083 461898 83125 462134
rect 82805 461866 83125 461898
rect 103874 462454 104194 462486
rect 103874 462218 103916 462454
rect 104152 462218 104194 462454
rect 103874 462134 104194 462218
rect 103874 461898 103916 462134
rect 104152 461898 104194 462134
rect 103874 461866 104194 461898
rect 109805 462454 110125 462486
rect 109805 462218 109847 462454
rect 110083 462218 110125 462454
rect 109805 462134 110125 462218
rect 109805 461898 109847 462134
rect 110083 461898 110125 462134
rect 109805 461866 110125 461898
rect 130874 462454 131194 462486
rect 130874 462218 130916 462454
rect 131152 462218 131194 462454
rect 130874 462134 131194 462218
rect 130874 461898 130916 462134
rect 131152 461898 131194 462134
rect 130874 461866 131194 461898
rect 136805 462454 137125 462486
rect 136805 462218 136847 462454
rect 137083 462218 137125 462454
rect 136805 462134 137125 462218
rect 136805 461898 136847 462134
rect 137083 461898 137125 462134
rect 136805 461866 137125 461898
rect 157874 462454 158194 462486
rect 157874 462218 157916 462454
rect 158152 462218 158194 462454
rect 157874 462134 158194 462218
rect 157874 461898 157916 462134
rect 158152 461898 158194 462134
rect 157874 461866 158194 461898
rect 163805 462454 164125 462486
rect 163805 462218 163847 462454
rect 164083 462218 164125 462454
rect 163805 462134 164125 462218
rect 163805 461898 163847 462134
rect 164083 461898 164125 462134
rect 163805 461866 164125 461898
rect 184874 462454 185194 462486
rect 184874 462218 184916 462454
rect 185152 462218 185194 462454
rect 184874 462134 185194 462218
rect 184874 461898 184916 462134
rect 185152 461898 185194 462134
rect 184874 461866 185194 461898
rect 190805 462454 191125 462486
rect 190805 462218 190847 462454
rect 191083 462218 191125 462454
rect 190805 462134 191125 462218
rect 190805 461898 190847 462134
rect 191083 461898 191125 462134
rect 190805 461866 191125 461898
rect 211874 462454 212194 462486
rect 211874 462218 211916 462454
rect 212152 462218 212194 462454
rect 211874 462134 212194 462218
rect 211874 461898 211916 462134
rect 212152 461898 212194 462134
rect 211874 461866 212194 461898
rect 217805 462454 218125 462486
rect 217805 462218 217847 462454
rect 218083 462218 218125 462454
rect 217805 462134 218125 462218
rect 217805 461898 217847 462134
rect 218083 461898 218125 462134
rect 217805 461866 218125 461898
rect 238874 462454 239194 462486
rect 238874 462218 238916 462454
rect 239152 462218 239194 462454
rect 238874 462134 239194 462218
rect 238874 461898 238916 462134
rect 239152 461898 239194 462134
rect 238874 461866 239194 461898
rect 244805 462454 245125 462486
rect 244805 462218 244847 462454
rect 245083 462218 245125 462454
rect 244805 462134 245125 462218
rect 244805 461898 244847 462134
rect 245083 461898 245125 462134
rect 244805 461866 245125 461898
rect 265874 462454 266194 462486
rect 265874 462218 265916 462454
rect 266152 462218 266194 462454
rect 265874 462134 266194 462218
rect 265874 461898 265916 462134
rect 266152 461898 266194 462134
rect 265874 461866 266194 461898
rect 271805 462454 272125 462486
rect 271805 462218 271847 462454
rect 272083 462218 272125 462454
rect 271805 462134 272125 462218
rect 271805 461898 271847 462134
rect 272083 461898 272125 462134
rect 271805 461866 272125 461898
rect 292874 462454 293194 462486
rect 292874 462218 292916 462454
rect 293152 462218 293194 462454
rect 292874 462134 293194 462218
rect 292874 461898 292916 462134
rect 293152 461898 293194 462134
rect 292874 461866 293194 461898
rect 298805 462454 299125 462486
rect 298805 462218 298847 462454
rect 299083 462218 299125 462454
rect 298805 462134 299125 462218
rect 298805 461898 298847 462134
rect 299083 461898 299125 462134
rect 298805 461866 299125 461898
rect 319874 462454 320194 462486
rect 319874 462218 319916 462454
rect 320152 462218 320194 462454
rect 319874 462134 320194 462218
rect 319874 461898 319916 462134
rect 320152 461898 320194 462134
rect 319874 461866 320194 461898
rect 325805 462454 326125 462486
rect 325805 462218 325847 462454
rect 326083 462218 326125 462454
rect 325805 462134 326125 462218
rect 325805 461898 325847 462134
rect 326083 461898 326125 462134
rect 325805 461866 326125 461898
rect 346874 462454 347194 462486
rect 346874 462218 346916 462454
rect 347152 462218 347194 462454
rect 346874 462134 347194 462218
rect 346874 461898 346916 462134
rect 347152 461898 347194 462134
rect 346874 461866 347194 461898
rect 352805 462454 353125 462486
rect 352805 462218 352847 462454
rect 353083 462218 353125 462454
rect 352805 462134 353125 462218
rect 352805 461898 352847 462134
rect 353083 461898 353125 462134
rect 352805 461866 353125 461898
rect 373874 462454 374194 462486
rect 373874 462218 373916 462454
rect 374152 462218 374194 462454
rect 373874 462134 374194 462218
rect 373874 461898 373916 462134
rect 374152 461898 374194 462134
rect 373874 461866 374194 461898
rect 379805 462454 380125 462486
rect 379805 462218 379847 462454
rect 380083 462218 380125 462454
rect 379805 462134 380125 462218
rect 379805 461898 379847 462134
rect 380083 461898 380125 462134
rect 379805 461866 380125 461898
rect 400874 462454 401194 462486
rect 400874 462218 400916 462454
rect 401152 462218 401194 462454
rect 400874 462134 401194 462218
rect 400874 461898 400916 462134
rect 401152 461898 401194 462134
rect 400874 461866 401194 461898
rect 406805 462454 407125 462486
rect 406805 462218 406847 462454
rect 407083 462218 407125 462454
rect 406805 462134 407125 462218
rect 406805 461898 406847 462134
rect 407083 461898 407125 462134
rect 406805 461866 407125 461898
rect 427874 462454 428194 462486
rect 427874 462218 427916 462454
rect 428152 462218 428194 462454
rect 427874 462134 428194 462218
rect 427874 461898 427916 462134
rect 428152 461898 428194 462134
rect 427874 461866 428194 461898
rect 433805 462454 434125 462486
rect 433805 462218 433847 462454
rect 434083 462218 434125 462454
rect 433805 462134 434125 462218
rect 433805 461898 433847 462134
rect 434083 461898 434125 462134
rect 433805 461866 434125 461898
rect 454874 462454 455194 462486
rect 454874 462218 454916 462454
rect 455152 462218 455194 462454
rect 454874 462134 455194 462218
rect 454874 461898 454916 462134
rect 455152 461898 455194 462134
rect 454874 461866 455194 461898
rect 460805 462454 461125 462486
rect 460805 462218 460847 462454
rect 461083 462218 461125 462454
rect 460805 462134 461125 462218
rect 460805 461898 460847 462134
rect 461083 461898 461125 462134
rect 460805 461866 461125 461898
rect 481874 462454 482194 462486
rect 481874 462218 481916 462454
rect 482152 462218 482194 462454
rect 481874 462134 482194 462218
rect 481874 461898 481916 462134
rect 482152 461898 482194 462134
rect 481874 461866 482194 461898
rect 487805 462454 488125 462486
rect 487805 462218 487847 462454
rect 488083 462218 488125 462454
rect 487805 462134 488125 462218
rect 487805 461898 487847 462134
rect 488083 461898 488125 462134
rect 487805 461866 488125 461898
rect 508874 462454 509194 462486
rect 508874 462218 508916 462454
rect 509152 462218 509194 462454
rect 508874 462134 509194 462218
rect 508874 461898 508916 462134
rect 509152 461898 509194 462134
rect 508874 461866 509194 461898
rect 514805 462454 515125 462486
rect 514805 462218 514847 462454
rect 515083 462218 515125 462454
rect 514805 462134 515125 462218
rect 514805 461898 514847 462134
rect 515083 461898 515125 462134
rect 514805 461866 515125 461898
rect 535874 462454 536194 462486
rect 535874 462218 535916 462454
rect 536152 462218 536194 462454
rect 535874 462134 536194 462218
rect 535874 461898 535916 462134
rect 536152 461898 536194 462134
rect 535874 461866 536194 461898
rect 541805 462454 542125 462486
rect 541805 462218 541847 462454
rect 542083 462218 542125 462454
rect 541805 462134 542125 462218
rect 541805 461898 541847 462134
rect 542083 461898 542125 462134
rect 541805 461866 542125 461898
rect 19910 453454 20230 453486
rect 19910 453218 19952 453454
rect 20188 453218 20230 453454
rect 19910 453134 20230 453218
rect 19910 452898 19952 453134
rect 20188 452898 20230 453134
rect 19910 452866 20230 452898
rect 25840 453454 26160 453486
rect 25840 453218 25882 453454
rect 26118 453218 26160 453454
rect 25840 453134 26160 453218
rect 25840 452898 25882 453134
rect 26118 452898 26160 453134
rect 25840 452866 26160 452898
rect 31771 453454 32091 453486
rect 31771 453218 31813 453454
rect 32049 453218 32091 453454
rect 31771 453134 32091 453218
rect 31771 452898 31813 453134
rect 32049 452898 32091 453134
rect 31771 452866 32091 452898
rect 46910 453454 47230 453486
rect 46910 453218 46952 453454
rect 47188 453218 47230 453454
rect 46910 453134 47230 453218
rect 46910 452898 46952 453134
rect 47188 452898 47230 453134
rect 46910 452866 47230 452898
rect 52840 453454 53160 453486
rect 52840 453218 52882 453454
rect 53118 453218 53160 453454
rect 52840 453134 53160 453218
rect 52840 452898 52882 453134
rect 53118 452898 53160 453134
rect 52840 452866 53160 452898
rect 58771 453454 59091 453486
rect 58771 453218 58813 453454
rect 59049 453218 59091 453454
rect 58771 453134 59091 453218
rect 58771 452898 58813 453134
rect 59049 452898 59091 453134
rect 58771 452866 59091 452898
rect 73910 453454 74230 453486
rect 73910 453218 73952 453454
rect 74188 453218 74230 453454
rect 73910 453134 74230 453218
rect 73910 452898 73952 453134
rect 74188 452898 74230 453134
rect 73910 452866 74230 452898
rect 79840 453454 80160 453486
rect 79840 453218 79882 453454
rect 80118 453218 80160 453454
rect 79840 453134 80160 453218
rect 79840 452898 79882 453134
rect 80118 452898 80160 453134
rect 79840 452866 80160 452898
rect 85771 453454 86091 453486
rect 85771 453218 85813 453454
rect 86049 453218 86091 453454
rect 85771 453134 86091 453218
rect 85771 452898 85813 453134
rect 86049 452898 86091 453134
rect 85771 452866 86091 452898
rect 100910 453454 101230 453486
rect 100910 453218 100952 453454
rect 101188 453218 101230 453454
rect 100910 453134 101230 453218
rect 100910 452898 100952 453134
rect 101188 452898 101230 453134
rect 100910 452866 101230 452898
rect 106840 453454 107160 453486
rect 106840 453218 106882 453454
rect 107118 453218 107160 453454
rect 106840 453134 107160 453218
rect 106840 452898 106882 453134
rect 107118 452898 107160 453134
rect 106840 452866 107160 452898
rect 112771 453454 113091 453486
rect 112771 453218 112813 453454
rect 113049 453218 113091 453454
rect 112771 453134 113091 453218
rect 112771 452898 112813 453134
rect 113049 452898 113091 453134
rect 112771 452866 113091 452898
rect 127910 453454 128230 453486
rect 127910 453218 127952 453454
rect 128188 453218 128230 453454
rect 127910 453134 128230 453218
rect 127910 452898 127952 453134
rect 128188 452898 128230 453134
rect 127910 452866 128230 452898
rect 133840 453454 134160 453486
rect 133840 453218 133882 453454
rect 134118 453218 134160 453454
rect 133840 453134 134160 453218
rect 133840 452898 133882 453134
rect 134118 452898 134160 453134
rect 133840 452866 134160 452898
rect 139771 453454 140091 453486
rect 139771 453218 139813 453454
rect 140049 453218 140091 453454
rect 139771 453134 140091 453218
rect 139771 452898 139813 453134
rect 140049 452898 140091 453134
rect 139771 452866 140091 452898
rect 154910 453454 155230 453486
rect 154910 453218 154952 453454
rect 155188 453218 155230 453454
rect 154910 453134 155230 453218
rect 154910 452898 154952 453134
rect 155188 452898 155230 453134
rect 154910 452866 155230 452898
rect 160840 453454 161160 453486
rect 160840 453218 160882 453454
rect 161118 453218 161160 453454
rect 160840 453134 161160 453218
rect 160840 452898 160882 453134
rect 161118 452898 161160 453134
rect 160840 452866 161160 452898
rect 166771 453454 167091 453486
rect 166771 453218 166813 453454
rect 167049 453218 167091 453454
rect 166771 453134 167091 453218
rect 166771 452898 166813 453134
rect 167049 452898 167091 453134
rect 166771 452866 167091 452898
rect 181910 453454 182230 453486
rect 181910 453218 181952 453454
rect 182188 453218 182230 453454
rect 181910 453134 182230 453218
rect 181910 452898 181952 453134
rect 182188 452898 182230 453134
rect 181910 452866 182230 452898
rect 187840 453454 188160 453486
rect 187840 453218 187882 453454
rect 188118 453218 188160 453454
rect 187840 453134 188160 453218
rect 187840 452898 187882 453134
rect 188118 452898 188160 453134
rect 187840 452866 188160 452898
rect 193771 453454 194091 453486
rect 193771 453218 193813 453454
rect 194049 453218 194091 453454
rect 193771 453134 194091 453218
rect 193771 452898 193813 453134
rect 194049 452898 194091 453134
rect 193771 452866 194091 452898
rect 208910 453454 209230 453486
rect 208910 453218 208952 453454
rect 209188 453218 209230 453454
rect 208910 453134 209230 453218
rect 208910 452898 208952 453134
rect 209188 452898 209230 453134
rect 208910 452866 209230 452898
rect 214840 453454 215160 453486
rect 214840 453218 214882 453454
rect 215118 453218 215160 453454
rect 214840 453134 215160 453218
rect 214840 452898 214882 453134
rect 215118 452898 215160 453134
rect 214840 452866 215160 452898
rect 220771 453454 221091 453486
rect 220771 453218 220813 453454
rect 221049 453218 221091 453454
rect 220771 453134 221091 453218
rect 220771 452898 220813 453134
rect 221049 452898 221091 453134
rect 220771 452866 221091 452898
rect 235910 453454 236230 453486
rect 235910 453218 235952 453454
rect 236188 453218 236230 453454
rect 235910 453134 236230 453218
rect 235910 452898 235952 453134
rect 236188 452898 236230 453134
rect 235910 452866 236230 452898
rect 241840 453454 242160 453486
rect 241840 453218 241882 453454
rect 242118 453218 242160 453454
rect 241840 453134 242160 453218
rect 241840 452898 241882 453134
rect 242118 452898 242160 453134
rect 241840 452866 242160 452898
rect 247771 453454 248091 453486
rect 247771 453218 247813 453454
rect 248049 453218 248091 453454
rect 247771 453134 248091 453218
rect 247771 452898 247813 453134
rect 248049 452898 248091 453134
rect 247771 452866 248091 452898
rect 262910 453454 263230 453486
rect 262910 453218 262952 453454
rect 263188 453218 263230 453454
rect 262910 453134 263230 453218
rect 262910 452898 262952 453134
rect 263188 452898 263230 453134
rect 262910 452866 263230 452898
rect 268840 453454 269160 453486
rect 268840 453218 268882 453454
rect 269118 453218 269160 453454
rect 268840 453134 269160 453218
rect 268840 452898 268882 453134
rect 269118 452898 269160 453134
rect 268840 452866 269160 452898
rect 274771 453454 275091 453486
rect 274771 453218 274813 453454
rect 275049 453218 275091 453454
rect 274771 453134 275091 453218
rect 274771 452898 274813 453134
rect 275049 452898 275091 453134
rect 274771 452866 275091 452898
rect 289910 453454 290230 453486
rect 289910 453218 289952 453454
rect 290188 453218 290230 453454
rect 289910 453134 290230 453218
rect 289910 452898 289952 453134
rect 290188 452898 290230 453134
rect 289910 452866 290230 452898
rect 295840 453454 296160 453486
rect 295840 453218 295882 453454
rect 296118 453218 296160 453454
rect 295840 453134 296160 453218
rect 295840 452898 295882 453134
rect 296118 452898 296160 453134
rect 295840 452866 296160 452898
rect 301771 453454 302091 453486
rect 301771 453218 301813 453454
rect 302049 453218 302091 453454
rect 301771 453134 302091 453218
rect 301771 452898 301813 453134
rect 302049 452898 302091 453134
rect 301771 452866 302091 452898
rect 316910 453454 317230 453486
rect 316910 453218 316952 453454
rect 317188 453218 317230 453454
rect 316910 453134 317230 453218
rect 316910 452898 316952 453134
rect 317188 452898 317230 453134
rect 316910 452866 317230 452898
rect 322840 453454 323160 453486
rect 322840 453218 322882 453454
rect 323118 453218 323160 453454
rect 322840 453134 323160 453218
rect 322840 452898 322882 453134
rect 323118 452898 323160 453134
rect 322840 452866 323160 452898
rect 328771 453454 329091 453486
rect 328771 453218 328813 453454
rect 329049 453218 329091 453454
rect 328771 453134 329091 453218
rect 328771 452898 328813 453134
rect 329049 452898 329091 453134
rect 328771 452866 329091 452898
rect 343910 453454 344230 453486
rect 343910 453218 343952 453454
rect 344188 453218 344230 453454
rect 343910 453134 344230 453218
rect 343910 452898 343952 453134
rect 344188 452898 344230 453134
rect 343910 452866 344230 452898
rect 349840 453454 350160 453486
rect 349840 453218 349882 453454
rect 350118 453218 350160 453454
rect 349840 453134 350160 453218
rect 349840 452898 349882 453134
rect 350118 452898 350160 453134
rect 349840 452866 350160 452898
rect 355771 453454 356091 453486
rect 355771 453218 355813 453454
rect 356049 453218 356091 453454
rect 355771 453134 356091 453218
rect 355771 452898 355813 453134
rect 356049 452898 356091 453134
rect 355771 452866 356091 452898
rect 370910 453454 371230 453486
rect 370910 453218 370952 453454
rect 371188 453218 371230 453454
rect 370910 453134 371230 453218
rect 370910 452898 370952 453134
rect 371188 452898 371230 453134
rect 370910 452866 371230 452898
rect 376840 453454 377160 453486
rect 376840 453218 376882 453454
rect 377118 453218 377160 453454
rect 376840 453134 377160 453218
rect 376840 452898 376882 453134
rect 377118 452898 377160 453134
rect 376840 452866 377160 452898
rect 382771 453454 383091 453486
rect 382771 453218 382813 453454
rect 383049 453218 383091 453454
rect 382771 453134 383091 453218
rect 382771 452898 382813 453134
rect 383049 452898 383091 453134
rect 382771 452866 383091 452898
rect 397910 453454 398230 453486
rect 397910 453218 397952 453454
rect 398188 453218 398230 453454
rect 397910 453134 398230 453218
rect 397910 452898 397952 453134
rect 398188 452898 398230 453134
rect 397910 452866 398230 452898
rect 403840 453454 404160 453486
rect 403840 453218 403882 453454
rect 404118 453218 404160 453454
rect 403840 453134 404160 453218
rect 403840 452898 403882 453134
rect 404118 452898 404160 453134
rect 403840 452866 404160 452898
rect 409771 453454 410091 453486
rect 409771 453218 409813 453454
rect 410049 453218 410091 453454
rect 409771 453134 410091 453218
rect 409771 452898 409813 453134
rect 410049 452898 410091 453134
rect 409771 452866 410091 452898
rect 424910 453454 425230 453486
rect 424910 453218 424952 453454
rect 425188 453218 425230 453454
rect 424910 453134 425230 453218
rect 424910 452898 424952 453134
rect 425188 452898 425230 453134
rect 424910 452866 425230 452898
rect 430840 453454 431160 453486
rect 430840 453218 430882 453454
rect 431118 453218 431160 453454
rect 430840 453134 431160 453218
rect 430840 452898 430882 453134
rect 431118 452898 431160 453134
rect 430840 452866 431160 452898
rect 436771 453454 437091 453486
rect 436771 453218 436813 453454
rect 437049 453218 437091 453454
rect 436771 453134 437091 453218
rect 436771 452898 436813 453134
rect 437049 452898 437091 453134
rect 436771 452866 437091 452898
rect 451910 453454 452230 453486
rect 451910 453218 451952 453454
rect 452188 453218 452230 453454
rect 451910 453134 452230 453218
rect 451910 452898 451952 453134
rect 452188 452898 452230 453134
rect 451910 452866 452230 452898
rect 457840 453454 458160 453486
rect 457840 453218 457882 453454
rect 458118 453218 458160 453454
rect 457840 453134 458160 453218
rect 457840 452898 457882 453134
rect 458118 452898 458160 453134
rect 457840 452866 458160 452898
rect 463771 453454 464091 453486
rect 463771 453218 463813 453454
rect 464049 453218 464091 453454
rect 463771 453134 464091 453218
rect 463771 452898 463813 453134
rect 464049 452898 464091 453134
rect 463771 452866 464091 452898
rect 478910 453454 479230 453486
rect 478910 453218 478952 453454
rect 479188 453218 479230 453454
rect 478910 453134 479230 453218
rect 478910 452898 478952 453134
rect 479188 452898 479230 453134
rect 478910 452866 479230 452898
rect 484840 453454 485160 453486
rect 484840 453218 484882 453454
rect 485118 453218 485160 453454
rect 484840 453134 485160 453218
rect 484840 452898 484882 453134
rect 485118 452898 485160 453134
rect 484840 452866 485160 452898
rect 490771 453454 491091 453486
rect 490771 453218 490813 453454
rect 491049 453218 491091 453454
rect 490771 453134 491091 453218
rect 490771 452898 490813 453134
rect 491049 452898 491091 453134
rect 490771 452866 491091 452898
rect 505910 453454 506230 453486
rect 505910 453218 505952 453454
rect 506188 453218 506230 453454
rect 505910 453134 506230 453218
rect 505910 452898 505952 453134
rect 506188 452898 506230 453134
rect 505910 452866 506230 452898
rect 511840 453454 512160 453486
rect 511840 453218 511882 453454
rect 512118 453218 512160 453454
rect 511840 453134 512160 453218
rect 511840 452898 511882 453134
rect 512118 452898 512160 453134
rect 511840 452866 512160 452898
rect 517771 453454 518091 453486
rect 517771 453218 517813 453454
rect 518049 453218 518091 453454
rect 517771 453134 518091 453218
rect 517771 452898 517813 453134
rect 518049 452898 518091 453134
rect 517771 452866 518091 452898
rect 532910 453454 533230 453486
rect 532910 453218 532952 453454
rect 533188 453218 533230 453454
rect 532910 453134 533230 453218
rect 532910 452898 532952 453134
rect 533188 452898 533230 453134
rect 532910 452866 533230 452898
rect 538840 453454 539160 453486
rect 538840 453218 538882 453454
rect 539118 453218 539160 453454
rect 538840 453134 539160 453218
rect 538840 452898 538882 453134
rect 539118 452898 539160 453134
rect 538840 452866 539160 452898
rect 544771 453454 545091 453486
rect 544771 453218 544813 453454
rect 545049 453218 545091 453454
rect 544771 453134 545091 453218
rect 544771 452898 544813 453134
rect 545049 452898 545091 453134
rect 544771 452866 545091 452898
rect 559794 453454 560414 470898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 426454 11414 443898
rect 19794 445394 20414 446000
rect 19794 445158 19826 445394
rect 20062 445158 20146 445394
rect 20382 445158 20414 445394
rect 19794 445074 20414 445158
rect 19794 444838 19826 445074
rect 20062 444838 20146 445074
rect 20382 444838 20414 445074
rect 19794 443000 20414 444838
rect 28794 444454 29414 446000
rect 28794 444218 28826 444454
rect 29062 444218 29146 444454
rect 29382 444218 29414 444454
rect 28794 444134 29414 444218
rect 28794 443898 28826 444134
rect 29062 443898 29146 444134
rect 29382 443898 29414 444134
rect 28794 443000 29414 443898
rect 37794 445394 38414 446000
rect 37794 445158 37826 445394
rect 38062 445158 38146 445394
rect 38382 445158 38414 445394
rect 37794 445074 38414 445158
rect 37794 444838 37826 445074
rect 38062 444838 38146 445074
rect 38382 444838 38414 445074
rect 37794 443000 38414 444838
rect 46794 444454 47414 446000
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 443000 47414 443898
rect 55794 445394 56414 446000
rect 55794 445158 55826 445394
rect 56062 445158 56146 445394
rect 56382 445158 56414 445394
rect 55794 445074 56414 445158
rect 55794 444838 55826 445074
rect 56062 444838 56146 445074
rect 56382 444838 56414 445074
rect 55794 443000 56414 444838
rect 64794 444454 65414 446000
rect 64794 444218 64826 444454
rect 65062 444218 65146 444454
rect 65382 444218 65414 444454
rect 64794 444134 65414 444218
rect 64794 443898 64826 444134
rect 65062 443898 65146 444134
rect 65382 443898 65414 444134
rect 64794 443000 65414 443898
rect 73794 445394 74414 446000
rect 73794 445158 73826 445394
rect 74062 445158 74146 445394
rect 74382 445158 74414 445394
rect 73794 445074 74414 445158
rect 73794 444838 73826 445074
rect 74062 444838 74146 445074
rect 74382 444838 74414 445074
rect 73794 443000 74414 444838
rect 82794 444454 83414 446000
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 443000 83414 443898
rect 91794 445394 92414 446000
rect 91794 445158 91826 445394
rect 92062 445158 92146 445394
rect 92382 445158 92414 445394
rect 91794 445074 92414 445158
rect 91794 444838 91826 445074
rect 92062 444838 92146 445074
rect 92382 444838 92414 445074
rect 91794 443000 92414 444838
rect 100794 444454 101414 446000
rect 100794 444218 100826 444454
rect 101062 444218 101146 444454
rect 101382 444218 101414 444454
rect 100794 444134 101414 444218
rect 100794 443898 100826 444134
rect 101062 443898 101146 444134
rect 101382 443898 101414 444134
rect 100794 443000 101414 443898
rect 109794 445394 110414 446000
rect 109794 445158 109826 445394
rect 110062 445158 110146 445394
rect 110382 445158 110414 445394
rect 109794 445074 110414 445158
rect 109794 444838 109826 445074
rect 110062 444838 110146 445074
rect 110382 444838 110414 445074
rect 109794 443000 110414 444838
rect 118794 444454 119414 446000
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 443000 119414 443898
rect 127794 445394 128414 446000
rect 127794 445158 127826 445394
rect 128062 445158 128146 445394
rect 128382 445158 128414 445394
rect 127794 445074 128414 445158
rect 127794 444838 127826 445074
rect 128062 444838 128146 445074
rect 128382 444838 128414 445074
rect 127794 443000 128414 444838
rect 136794 444454 137414 446000
rect 136794 444218 136826 444454
rect 137062 444218 137146 444454
rect 137382 444218 137414 444454
rect 136794 444134 137414 444218
rect 136794 443898 136826 444134
rect 137062 443898 137146 444134
rect 137382 443898 137414 444134
rect 136794 443000 137414 443898
rect 145794 445394 146414 446000
rect 145794 445158 145826 445394
rect 146062 445158 146146 445394
rect 146382 445158 146414 445394
rect 145794 445074 146414 445158
rect 145794 444838 145826 445074
rect 146062 444838 146146 445074
rect 146382 444838 146414 445074
rect 145794 443000 146414 444838
rect 154794 444454 155414 446000
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 443000 155414 443898
rect 163794 445394 164414 446000
rect 163794 445158 163826 445394
rect 164062 445158 164146 445394
rect 164382 445158 164414 445394
rect 163794 445074 164414 445158
rect 163794 444838 163826 445074
rect 164062 444838 164146 445074
rect 164382 444838 164414 445074
rect 163794 443000 164414 444838
rect 172794 444454 173414 446000
rect 172794 444218 172826 444454
rect 173062 444218 173146 444454
rect 173382 444218 173414 444454
rect 172794 444134 173414 444218
rect 172794 443898 172826 444134
rect 173062 443898 173146 444134
rect 173382 443898 173414 444134
rect 172794 443000 173414 443898
rect 181794 445394 182414 446000
rect 181794 445158 181826 445394
rect 182062 445158 182146 445394
rect 182382 445158 182414 445394
rect 181794 445074 182414 445158
rect 181794 444838 181826 445074
rect 182062 444838 182146 445074
rect 182382 444838 182414 445074
rect 181794 443000 182414 444838
rect 190794 444454 191414 446000
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 443000 191414 443898
rect 199794 445394 200414 446000
rect 199794 445158 199826 445394
rect 200062 445158 200146 445394
rect 200382 445158 200414 445394
rect 199794 445074 200414 445158
rect 199794 444838 199826 445074
rect 200062 444838 200146 445074
rect 200382 444838 200414 445074
rect 199794 443000 200414 444838
rect 208794 444454 209414 446000
rect 208794 444218 208826 444454
rect 209062 444218 209146 444454
rect 209382 444218 209414 444454
rect 208794 444134 209414 444218
rect 208794 443898 208826 444134
rect 209062 443898 209146 444134
rect 209382 443898 209414 444134
rect 208794 443000 209414 443898
rect 217794 445394 218414 446000
rect 217794 445158 217826 445394
rect 218062 445158 218146 445394
rect 218382 445158 218414 445394
rect 217794 445074 218414 445158
rect 217794 444838 217826 445074
rect 218062 444838 218146 445074
rect 218382 444838 218414 445074
rect 217794 443000 218414 444838
rect 226794 444454 227414 446000
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 443000 227414 443898
rect 235794 445394 236414 446000
rect 235794 445158 235826 445394
rect 236062 445158 236146 445394
rect 236382 445158 236414 445394
rect 235794 445074 236414 445158
rect 235794 444838 235826 445074
rect 236062 444838 236146 445074
rect 236382 444838 236414 445074
rect 235794 443000 236414 444838
rect 244794 444454 245414 446000
rect 244794 444218 244826 444454
rect 245062 444218 245146 444454
rect 245382 444218 245414 444454
rect 244794 444134 245414 444218
rect 244794 443898 244826 444134
rect 245062 443898 245146 444134
rect 245382 443898 245414 444134
rect 244794 443000 245414 443898
rect 253794 445394 254414 446000
rect 253794 445158 253826 445394
rect 254062 445158 254146 445394
rect 254382 445158 254414 445394
rect 253794 445074 254414 445158
rect 253794 444838 253826 445074
rect 254062 444838 254146 445074
rect 254382 444838 254414 445074
rect 253794 443000 254414 444838
rect 262794 444454 263414 446000
rect 262794 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 263414 444454
rect 262794 444134 263414 444218
rect 262794 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 263414 444134
rect 262794 443000 263414 443898
rect 271794 445394 272414 446000
rect 271794 445158 271826 445394
rect 272062 445158 272146 445394
rect 272382 445158 272414 445394
rect 271794 445074 272414 445158
rect 271794 444838 271826 445074
rect 272062 444838 272146 445074
rect 272382 444838 272414 445074
rect 271794 443000 272414 444838
rect 280794 444454 281414 446000
rect 280794 444218 280826 444454
rect 281062 444218 281146 444454
rect 281382 444218 281414 444454
rect 280794 444134 281414 444218
rect 280794 443898 280826 444134
rect 281062 443898 281146 444134
rect 281382 443898 281414 444134
rect 280794 443000 281414 443898
rect 289794 445394 290414 446000
rect 289794 445158 289826 445394
rect 290062 445158 290146 445394
rect 290382 445158 290414 445394
rect 289794 445074 290414 445158
rect 289794 444838 289826 445074
rect 290062 444838 290146 445074
rect 290382 444838 290414 445074
rect 289794 443000 290414 444838
rect 298794 444454 299414 446000
rect 298794 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 299414 444454
rect 298794 444134 299414 444218
rect 298794 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 299414 444134
rect 298794 443000 299414 443898
rect 307794 445394 308414 446000
rect 307794 445158 307826 445394
rect 308062 445158 308146 445394
rect 308382 445158 308414 445394
rect 307794 445074 308414 445158
rect 307794 444838 307826 445074
rect 308062 444838 308146 445074
rect 308382 444838 308414 445074
rect 307794 443000 308414 444838
rect 316794 444454 317414 446000
rect 316794 444218 316826 444454
rect 317062 444218 317146 444454
rect 317382 444218 317414 444454
rect 316794 444134 317414 444218
rect 316794 443898 316826 444134
rect 317062 443898 317146 444134
rect 317382 443898 317414 444134
rect 316794 443000 317414 443898
rect 325794 445394 326414 446000
rect 325794 445158 325826 445394
rect 326062 445158 326146 445394
rect 326382 445158 326414 445394
rect 325794 445074 326414 445158
rect 325794 444838 325826 445074
rect 326062 444838 326146 445074
rect 326382 444838 326414 445074
rect 325794 443000 326414 444838
rect 334794 444454 335414 446000
rect 334794 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 335414 444454
rect 334794 444134 335414 444218
rect 334794 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 335414 444134
rect 334794 443000 335414 443898
rect 343794 445394 344414 446000
rect 343794 445158 343826 445394
rect 344062 445158 344146 445394
rect 344382 445158 344414 445394
rect 343794 445074 344414 445158
rect 343794 444838 343826 445074
rect 344062 444838 344146 445074
rect 344382 444838 344414 445074
rect 343794 443000 344414 444838
rect 352794 444454 353414 446000
rect 352794 444218 352826 444454
rect 353062 444218 353146 444454
rect 353382 444218 353414 444454
rect 352794 444134 353414 444218
rect 352794 443898 352826 444134
rect 353062 443898 353146 444134
rect 353382 443898 353414 444134
rect 352794 443000 353414 443898
rect 361794 445394 362414 446000
rect 361794 445158 361826 445394
rect 362062 445158 362146 445394
rect 362382 445158 362414 445394
rect 361794 445074 362414 445158
rect 361794 444838 361826 445074
rect 362062 444838 362146 445074
rect 362382 444838 362414 445074
rect 361794 443000 362414 444838
rect 370794 444454 371414 446000
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 443000 371414 443898
rect 379794 445394 380414 446000
rect 379794 445158 379826 445394
rect 380062 445158 380146 445394
rect 380382 445158 380414 445394
rect 379794 445074 380414 445158
rect 379794 444838 379826 445074
rect 380062 444838 380146 445074
rect 380382 444838 380414 445074
rect 379794 443000 380414 444838
rect 388794 444454 389414 446000
rect 388794 444218 388826 444454
rect 389062 444218 389146 444454
rect 389382 444218 389414 444454
rect 388794 444134 389414 444218
rect 388794 443898 388826 444134
rect 389062 443898 389146 444134
rect 389382 443898 389414 444134
rect 388794 443000 389414 443898
rect 397794 445394 398414 446000
rect 397794 445158 397826 445394
rect 398062 445158 398146 445394
rect 398382 445158 398414 445394
rect 397794 445074 398414 445158
rect 397794 444838 397826 445074
rect 398062 444838 398146 445074
rect 398382 444838 398414 445074
rect 397794 443000 398414 444838
rect 406794 444454 407414 446000
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 443000 407414 443898
rect 415794 445394 416414 446000
rect 415794 445158 415826 445394
rect 416062 445158 416146 445394
rect 416382 445158 416414 445394
rect 415794 445074 416414 445158
rect 415794 444838 415826 445074
rect 416062 444838 416146 445074
rect 416382 444838 416414 445074
rect 415794 443000 416414 444838
rect 424794 444454 425414 446000
rect 424794 444218 424826 444454
rect 425062 444218 425146 444454
rect 425382 444218 425414 444454
rect 424794 444134 425414 444218
rect 424794 443898 424826 444134
rect 425062 443898 425146 444134
rect 425382 443898 425414 444134
rect 424794 443000 425414 443898
rect 433794 445394 434414 446000
rect 433794 445158 433826 445394
rect 434062 445158 434146 445394
rect 434382 445158 434414 445394
rect 433794 445074 434414 445158
rect 433794 444838 433826 445074
rect 434062 444838 434146 445074
rect 434382 444838 434414 445074
rect 433794 443000 434414 444838
rect 442794 444454 443414 446000
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 443000 443414 443898
rect 451794 445394 452414 446000
rect 451794 445158 451826 445394
rect 452062 445158 452146 445394
rect 452382 445158 452414 445394
rect 451794 445074 452414 445158
rect 451794 444838 451826 445074
rect 452062 444838 452146 445074
rect 452382 444838 452414 445074
rect 451794 443000 452414 444838
rect 460794 444454 461414 446000
rect 460794 444218 460826 444454
rect 461062 444218 461146 444454
rect 461382 444218 461414 444454
rect 460794 444134 461414 444218
rect 460794 443898 460826 444134
rect 461062 443898 461146 444134
rect 461382 443898 461414 444134
rect 460794 443000 461414 443898
rect 469794 445394 470414 446000
rect 469794 445158 469826 445394
rect 470062 445158 470146 445394
rect 470382 445158 470414 445394
rect 469794 445074 470414 445158
rect 469794 444838 469826 445074
rect 470062 444838 470146 445074
rect 470382 444838 470414 445074
rect 469794 443000 470414 444838
rect 478794 444454 479414 446000
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 443000 479414 443898
rect 487794 445394 488414 446000
rect 487794 445158 487826 445394
rect 488062 445158 488146 445394
rect 488382 445158 488414 445394
rect 487794 445074 488414 445158
rect 487794 444838 487826 445074
rect 488062 444838 488146 445074
rect 488382 444838 488414 445074
rect 487794 443000 488414 444838
rect 496794 444454 497414 446000
rect 496794 444218 496826 444454
rect 497062 444218 497146 444454
rect 497382 444218 497414 444454
rect 496794 444134 497414 444218
rect 496794 443898 496826 444134
rect 497062 443898 497146 444134
rect 497382 443898 497414 444134
rect 496794 443000 497414 443898
rect 505794 445394 506414 446000
rect 505794 445158 505826 445394
rect 506062 445158 506146 445394
rect 506382 445158 506414 445394
rect 505794 445074 506414 445158
rect 505794 444838 505826 445074
rect 506062 444838 506146 445074
rect 506382 444838 506414 445074
rect 505794 443000 506414 444838
rect 514794 444454 515414 446000
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 443000 515414 443898
rect 523794 445394 524414 446000
rect 523794 445158 523826 445394
rect 524062 445158 524146 445394
rect 524382 445158 524414 445394
rect 523794 445074 524414 445158
rect 523794 444838 523826 445074
rect 524062 444838 524146 445074
rect 524382 444838 524414 445074
rect 523794 443000 524414 444838
rect 532794 444454 533414 446000
rect 532794 444218 532826 444454
rect 533062 444218 533146 444454
rect 533382 444218 533414 444454
rect 532794 444134 533414 444218
rect 532794 443898 532826 444134
rect 533062 443898 533146 444134
rect 533382 443898 533414 444134
rect 532794 443000 533414 443898
rect 541794 445394 542414 446000
rect 541794 445158 541826 445394
rect 542062 445158 542146 445394
rect 542382 445158 542414 445394
rect 541794 445074 542414 445158
rect 541794 444838 541826 445074
rect 542062 444838 542146 445074
rect 542382 444838 542414 445074
rect 541794 443000 542414 444838
rect 550794 444454 551414 446000
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 443000 551414 443898
rect 19910 435454 20230 435486
rect 19910 435218 19952 435454
rect 20188 435218 20230 435454
rect 19910 435134 20230 435218
rect 19910 434898 19952 435134
rect 20188 434898 20230 435134
rect 19910 434866 20230 434898
rect 25840 435454 26160 435486
rect 25840 435218 25882 435454
rect 26118 435218 26160 435454
rect 25840 435134 26160 435218
rect 25840 434898 25882 435134
rect 26118 434898 26160 435134
rect 25840 434866 26160 434898
rect 31771 435454 32091 435486
rect 31771 435218 31813 435454
rect 32049 435218 32091 435454
rect 31771 435134 32091 435218
rect 31771 434898 31813 435134
rect 32049 434898 32091 435134
rect 31771 434866 32091 434898
rect 46910 435454 47230 435486
rect 46910 435218 46952 435454
rect 47188 435218 47230 435454
rect 46910 435134 47230 435218
rect 46910 434898 46952 435134
rect 47188 434898 47230 435134
rect 46910 434866 47230 434898
rect 52840 435454 53160 435486
rect 52840 435218 52882 435454
rect 53118 435218 53160 435454
rect 52840 435134 53160 435218
rect 52840 434898 52882 435134
rect 53118 434898 53160 435134
rect 52840 434866 53160 434898
rect 58771 435454 59091 435486
rect 58771 435218 58813 435454
rect 59049 435218 59091 435454
rect 58771 435134 59091 435218
rect 58771 434898 58813 435134
rect 59049 434898 59091 435134
rect 58771 434866 59091 434898
rect 73910 435454 74230 435486
rect 73910 435218 73952 435454
rect 74188 435218 74230 435454
rect 73910 435134 74230 435218
rect 73910 434898 73952 435134
rect 74188 434898 74230 435134
rect 73910 434866 74230 434898
rect 79840 435454 80160 435486
rect 79840 435218 79882 435454
rect 80118 435218 80160 435454
rect 79840 435134 80160 435218
rect 79840 434898 79882 435134
rect 80118 434898 80160 435134
rect 79840 434866 80160 434898
rect 85771 435454 86091 435486
rect 85771 435218 85813 435454
rect 86049 435218 86091 435454
rect 85771 435134 86091 435218
rect 85771 434898 85813 435134
rect 86049 434898 86091 435134
rect 85771 434866 86091 434898
rect 100910 435454 101230 435486
rect 100910 435218 100952 435454
rect 101188 435218 101230 435454
rect 100910 435134 101230 435218
rect 100910 434898 100952 435134
rect 101188 434898 101230 435134
rect 100910 434866 101230 434898
rect 106840 435454 107160 435486
rect 106840 435218 106882 435454
rect 107118 435218 107160 435454
rect 106840 435134 107160 435218
rect 106840 434898 106882 435134
rect 107118 434898 107160 435134
rect 106840 434866 107160 434898
rect 112771 435454 113091 435486
rect 112771 435218 112813 435454
rect 113049 435218 113091 435454
rect 112771 435134 113091 435218
rect 112771 434898 112813 435134
rect 113049 434898 113091 435134
rect 112771 434866 113091 434898
rect 127910 435454 128230 435486
rect 127910 435218 127952 435454
rect 128188 435218 128230 435454
rect 127910 435134 128230 435218
rect 127910 434898 127952 435134
rect 128188 434898 128230 435134
rect 127910 434866 128230 434898
rect 133840 435454 134160 435486
rect 133840 435218 133882 435454
rect 134118 435218 134160 435454
rect 133840 435134 134160 435218
rect 133840 434898 133882 435134
rect 134118 434898 134160 435134
rect 133840 434866 134160 434898
rect 139771 435454 140091 435486
rect 139771 435218 139813 435454
rect 140049 435218 140091 435454
rect 139771 435134 140091 435218
rect 139771 434898 139813 435134
rect 140049 434898 140091 435134
rect 139771 434866 140091 434898
rect 154910 435454 155230 435486
rect 154910 435218 154952 435454
rect 155188 435218 155230 435454
rect 154910 435134 155230 435218
rect 154910 434898 154952 435134
rect 155188 434898 155230 435134
rect 154910 434866 155230 434898
rect 160840 435454 161160 435486
rect 160840 435218 160882 435454
rect 161118 435218 161160 435454
rect 160840 435134 161160 435218
rect 160840 434898 160882 435134
rect 161118 434898 161160 435134
rect 160840 434866 161160 434898
rect 166771 435454 167091 435486
rect 166771 435218 166813 435454
rect 167049 435218 167091 435454
rect 166771 435134 167091 435218
rect 166771 434898 166813 435134
rect 167049 434898 167091 435134
rect 166771 434866 167091 434898
rect 181910 435454 182230 435486
rect 181910 435218 181952 435454
rect 182188 435218 182230 435454
rect 181910 435134 182230 435218
rect 181910 434898 181952 435134
rect 182188 434898 182230 435134
rect 181910 434866 182230 434898
rect 187840 435454 188160 435486
rect 187840 435218 187882 435454
rect 188118 435218 188160 435454
rect 187840 435134 188160 435218
rect 187840 434898 187882 435134
rect 188118 434898 188160 435134
rect 187840 434866 188160 434898
rect 193771 435454 194091 435486
rect 193771 435218 193813 435454
rect 194049 435218 194091 435454
rect 193771 435134 194091 435218
rect 193771 434898 193813 435134
rect 194049 434898 194091 435134
rect 193771 434866 194091 434898
rect 208910 435454 209230 435486
rect 208910 435218 208952 435454
rect 209188 435218 209230 435454
rect 208910 435134 209230 435218
rect 208910 434898 208952 435134
rect 209188 434898 209230 435134
rect 208910 434866 209230 434898
rect 214840 435454 215160 435486
rect 214840 435218 214882 435454
rect 215118 435218 215160 435454
rect 214840 435134 215160 435218
rect 214840 434898 214882 435134
rect 215118 434898 215160 435134
rect 214840 434866 215160 434898
rect 220771 435454 221091 435486
rect 220771 435218 220813 435454
rect 221049 435218 221091 435454
rect 220771 435134 221091 435218
rect 220771 434898 220813 435134
rect 221049 434898 221091 435134
rect 220771 434866 221091 434898
rect 235910 435454 236230 435486
rect 235910 435218 235952 435454
rect 236188 435218 236230 435454
rect 235910 435134 236230 435218
rect 235910 434898 235952 435134
rect 236188 434898 236230 435134
rect 235910 434866 236230 434898
rect 241840 435454 242160 435486
rect 241840 435218 241882 435454
rect 242118 435218 242160 435454
rect 241840 435134 242160 435218
rect 241840 434898 241882 435134
rect 242118 434898 242160 435134
rect 241840 434866 242160 434898
rect 247771 435454 248091 435486
rect 247771 435218 247813 435454
rect 248049 435218 248091 435454
rect 247771 435134 248091 435218
rect 247771 434898 247813 435134
rect 248049 434898 248091 435134
rect 247771 434866 248091 434898
rect 262910 435454 263230 435486
rect 262910 435218 262952 435454
rect 263188 435218 263230 435454
rect 262910 435134 263230 435218
rect 262910 434898 262952 435134
rect 263188 434898 263230 435134
rect 262910 434866 263230 434898
rect 268840 435454 269160 435486
rect 268840 435218 268882 435454
rect 269118 435218 269160 435454
rect 268840 435134 269160 435218
rect 268840 434898 268882 435134
rect 269118 434898 269160 435134
rect 268840 434866 269160 434898
rect 274771 435454 275091 435486
rect 274771 435218 274813 435454
rect 275049 435218 275091 435454
rect 274771 435134 275091 435218
rect 274771 434898 274813 435134
rect 275049 434898 275091 435134
rect 274771 434866 275091 434898
rect 289910 435454 290230 435486
rect 289910 435218 289952 435454
rect 290188 435218 290230 435454
rect 289910 435134 290230 435218
rect 289910 434898 289952 435134
rect 290188 434898 290230 435134
rect 289910 434866 290230 434898
rect 295840 435454 296160 435486
rect 295840 435218 295882 435454
rect 296118 435218 296160 435454
rect 295840 435134 296160 435218
rect 295840 434898 295882 435134
rect 296118 434898 296160 435134
rect 295840 434866 296160 434898
rect 301771 435454 302091 435486
rect 301771 435218 301813 435454
rect 302049 435218 302091 435454
rect 301771 435134 302091 435218
rect 301771 434898 301813 435134
rect 302049 434898 302091 435134
rect 301771 434866 302091 434898
rect 316910 435454 317230 435486
rect 316910 435218 316952 435454
rect 317188 435218 317230 435454
rect 316910 435134 317230 435218
rect 316910 434898 316952 435134
rect 317188 434898 317230 435134
rect 316910 434866 317230 434898
rect 322840 435454 323160 435486
rect 322840 435218 322882 435454
rect 323118 435218 323160 435454
rect 322840 435134 323160 435218
rect 322840 434898 322882 435134
rect 323118 434898 323160 435134
rect 322840 434866 323160 434898
rect 328771 435454 329091 435486
rect 328771 435218 328813 435454
rect 329049 435218 329091 435454
rect 328771 435134 329091 435218
rect 328771 434898 328813 435134
rect 329049 434898 329091 435134
rect 328771 434866 329091 434898
rect 343910 435454 344230 435486
rect 343910 435218 343952 435454
rect 344188 435218 344230 435454
rect 343910 435134 344230 435218
rect 343910 434898 343952 435134
rect 344188 434898 344230 435134
rect 343910 434866 344230 434898
rect 349840 435454 350160 435486
rect 349840 435218 349882 435454
rect 350118 435218 350160 435454
rect 349840 435134 350160 435218
rect 349840 434898 349882 435134
rect 350118 434898 350160 435134
rect 349840 434866 350160 434898
rect 355771 435454 356091 435486
rect 355771 435218 355813 435454
rect 356049 435218 356091 435454
rect 355771 435134 356091 435218
rect 355771 434898 355813 435134
rect 356049 434898 356091 435134
rect 355771 434866 356091 434898
rect 370910 435454 371230 435486
rect 370910 435218 370952 435454
rect 371188 435218 371230 435454
rect 370910 435134 371230 435218
rect 370910 434898 370952 435134
rect 371188 434898 371230 435134
rect 370910 434866 371230 434898
rect 376840 435454 377160 435486
rect 376840 435218 376882 435454
rect 377118 435218 377160 435454
rect 376840 435134 377160 435218
rect 376840 434898 376882 435134
rect 377118 434898 377160 435134
rect 376840 434866 377160 434898
rect 382771 435454 383091 435486
rect 382771 435218 382813 435454
rect 383049 435218 383091 435454
rect 382771 435134 383091 435218
rect 382771 434898 382813 435134
rect 383049 434898 383091 435134
rect 382771 434866 383091 434898
rect 397910 435454 398230 435486
rect 397910 435218 397952 435454
rect 398188 435218 398230 435454
rect 397910 435134 398230 435218
rect 397910 434898 397952 435134
rect 398188 434898 398230 435134
rect 397910 434866 398230 434898
rect 403840 435454 404160 435486
rect 403840 435218 403882 435454
rect 404118 435218 404160 435454
rect 403840 435134 404160 435218
rect 403840 434898 403882 435134
rect 404118 434898 404160 435134
rect 403840 434866 404160 434898
rect 409771 435454 410091 435486
rect 409771 435218 409813 435454
rect 410049 435218 410091 435454
rect 409771 435134 410091 435218
rect 409771 434898 409813 435134
rect 410049 434898 410091 435134
rect 409771 434866 410091 434898
rect 424910 435454 425230 435486
rect 424910 435218 424952 435454
rect 425188 435218 425230 435454
rect 424910 435134 425230 435218
rect 424910 434898 424952 435134
rect 425188 434898 425230 435134
rect 424910 434866 425230 434898
rect 430840 435454 431160 435486
rect 430840 435218 430882 435454
rect 431118 435218 431160 435454
rect 430840 435134 431160 435218
rect 430840 434898 430882 435134
rect 431118 434898 431160 435134
rect 430840 434866 431160 434898
rect 436771 435454 437091 435486
rect 436771 435218 436813 435454
rect 437049 435218 437091 435454
rect 436771 435134 437091 435218
rect 436771 434898 436813 435134
rect 437049 434898 437091 435134
rect 436771 434866 437091 434898
rect 451910 435454 452230 435486
rect 451910 435218 451952 435454
rect 452188 435218 452230 435454
rect 451910 435134 452230 435218
rect 451910 434898 451952 435134
rect 452188 434898 452230 435134
rect 451910 434866 452230 434898
rect 457840 435454 458160 435486
rect 457840 435218 457882 435454
rect 458118 435218 458160 435454
rect 457840 435134 458160 435218
rect 457840 434898 457882 435134
rect 458118 434898 458160 435134
rect 457840 434866 458160 434898
rect 463771 435454 464091 435486
rect 463771 435218 463813 435454
rect 464049 435218 464091 435454
rect 463771 435134 464091 435218
rect 463771 434898 463813 435134
rect 464049 434898 464091 435134
rect 463771 434866 464091 434898
rect 478910 435454 479230 435486
rect 478910 435218 478952 435454
rect 479188 435218 479230 435454
rect 478910 435134 479230 435218
rect 478910 434898 478952 435134
rect 479188 434898 479230 435134
rect 478910 434866 479230 434898
rect 484840 435454 485160 435486
rect 484840 435218 484882 435454
rect 485118 435218 485160 435454
rect 484840 435134 485160 435218
rect 484840 434898 484882 435134
rect 485118 434898 485160 435134
rect 484840 434866 485160 434898
rect 490771 435454 491091 435486
rect 490771 435218 490813 435454
rect 491049 435218 491091 435454
rect 490771 435134 491091 435218
rect 490771 434898 490813 435134
rect 491049 434898 491091 435134
rect 490771 434866 491091 434898
rect 505910 435454 506230 435486
rect 505910 435218 505952 435454
rect 506188 435218 506230 435454
rect 505910 435134 506230 435218
rect 505910 434898 505952 435134
rect 506188 434898 506230 435134
rect 505910 434866 506230 434898
rect 511840 435454 512160 435486
rect 511840 435218 511882 435454
rect 512118 435218 512160 435454
rect 511840 435134 512160 435218
rect 511840 434898 511882 435134
rect 512118 434898 512160 435134
rect 511840 434866 512160 434898
rect 517771 435454 518091 435486
rect 517771 435218 517813 435454
rect 518049 435218 518091 435454
rect 517771 435134 518091 435218
rect 517771 434898 517813 435134
rect 518049 434898 518091 435134
rect 517771 434866 518091 434898
rect 532910 435454 533230 435486
rect 532910 435218 532952 435454
rect 533188 435218 533230 435454
rect 532910 435134 533230 435218
rect 532910 434898 532952 435134
rect 533188 434898 533230 435134
rect 532910 434866 533230 434898
rect 538840 435454 539160 435486
rect 538840 435218 538882 435454
rect 539118 435218 539160 435454
rect 538840 435134 539160 435218
rect 538840 434898 538882 435134
rect 539118 434898 539160 435134
rect 538840 434866 539160 434898
rect 544771 435454 545091 435486
rect 544771 435218 544813 435454
rect 545049 435218 545091 435454
rect 544771 435134 545091 435218
rect 544771 434898 544813 435134
rect 545049 434898 545091 435134
rect 544771 434866 545091 434898
rect 559794 435454 560414 452898
rect 559794 435218 559826 435454
rect 560062 435218 560146 435454
rect 560382 435218 560414 435454
rect 559794 435134 560414 435218
rect 559794 434898 559826 435134
rect 560062 434898 560146 435134
rect 560382 434898 560414 435134
rect 10794 426218 10826 426454
rect 11062 426218 11146 426454
rect 11382 426218 11414 426454
rect 10794 426134 11414 426218
rect 10794 425898 10826 426134
rect 11062 425898 11146 426134
rect 11382 425898 11414 426134
rect 10794 408454 11414 425898
rect 22874 426454 23194 426486
rect 22874 426218 22916 426454
rect 23152 426218 23194 426454
rect 22874 426134 23194 426218
rect 22874 425898 22916 426134
rect 23152 425898 23194 426134
rect 22874 425866 23194 425898
rect 28805 426454 29125 426486
rect 28805 426218 28847 426454
rect 29083 426218 29125 426454
rect 28805 426134 29125 426218
rect 28805 425898 28847 426134
rect 29083 425898 29125 426134
rect 28805 425866 29125 425898
rect 49874 426454 50194 426486
rect 49874 426218 49916 426454
rect 50152 426218 50194 426454
rect 49874 426134 50194 426218
rect 49874 425898 49916 426134
rect 50152 425898 50194 426134
rect 49874 425866 50194 425898
rect 55805 426454 56125 426486
rect 55805 426218 55847 426454
rect 56083 426218 56125 426454
rect 55805 426134 56125 426218
rect 55805 425898 55847 426134
rect 56083 425898 56125 426134
rect 55805 425866 56125 425898
rect 76874 426454 77194 426486
rect 76874 426218 76916 426454
rect 77152 426218 77194 426454
rect 76874 426134 77194 426218
rect 76874 425898 76916 426134
rect 77152 425898 77194 426134
rect 76874 425866 77194 425898
rect 82805 426454 83125 426486
rect 82805 426218 82847 426454
rect 83083 426218 83125 426454
rect 82805 426134 83125 426218
rect 82805 425898 82847 426134
rect 83083 425898 83125 426134
rect 82805 425866 83125 425898
rect 103874 426454 104194 426486
rect 103874 426218 103916 426454
rect 104152 426218 104194 426454
rect 103874 426134 104194 426218
rect 103874 425898 103916 426134
rect 104152 425898 104194 426134
rect 103874 425866 104194 425898
rect 109805 426454 110125 426486
rect 109805 426218 109847 426454
rect 110083 426218 110125 426454
rect 109805 426134 110125 426218
rect 109805 425898 109847 426134
rect 110083 425898 110125 426134
rect 109805 425866 110125 425898
rect 130874 426454 131194 426486
rect 130874 426218 130916 426454
rect 131152 426218 131194 426454
rect 130874 426134 131194 426218
rect 130874 425898 130916 426134
rect 131152 425898 131194 426134
rect 130874 425866 131194 425898
rect 136805 426454 137125 426486
rect 136805 426218 136847 426454
rect 137083 426218 137125 426454
rect 136805 426134 137125 426218
rect 136805 425898 136847 426134
rect 137083 425898 137125 426134
rect 136805 425866 137125 425898
rect 157874 426454 158194 426486
rect 157874 426218 157916 426454
rect 158152 426218 158194 426454
rect 157874 426134 158194 426218
rect 157874 425898 157916 426134
rect 158152 425898 158194 426134
rect 157874 425866 158194 425898
rect 163805 426454 164125 426486
rect 163805 426218 163847 426454
rect 164083 426218 164125 426454
rect 163805 426134 164125 426218
rect 163805 425898 163847 426134
rect 164083 425898 164125 426134
rect 163805 425866 164125 425898
rect 184874 426454 185194 426486
rect 184874 426218 184916 426454
rect 185152 426218 185194 426454
rect 184874 426134 185194 426218
rect 184874 425898 184916 426134
rect 185152 425898 185194 426134
rect 184874 425866 185194 425898
rect 190805 426454 191125 426486
rect 190805 426218 190847 426454
rect 191083 426218 191125 426454
rect 190805 426134 191125 426218
rect 190805 425898 190847 426134
rect 191083 425898 191125 426134
rect 190805 425866 191125 425898
rect 211874 426454 212194 426486
rect 211874 426218 211916 426454
rect 212152 426218 212194 426454
rect 211874 426134 212194 426218
rect 211874 425898 211916 426134
rect 212152 425898 212194 426134
rect 211874 425866 212194 425898
rect 217805 426454 218125 426486
rect 217805 426218 217847 426454
rect 218083 426218 218125 426454
rect 217805 426134 218125 426218
rect 217805 425898 217847 426134
rect 218083 425898 218125 426134
rect 217805 425866 218125 425898
rect 238874 426454 239194 426486
rect 238874 426218 238916 426454
rect 239152 426218 239194 426454
rect 238874 426134 239194 426218
rect 238874 425898 238916 426134
rect 239152 425898 239194 426134
rect 238874 425866 239194 425898
rect 244805 426454 245125 426486
rect 244805 426218 244847 426454
rect 245083 426218 245125 426454
rect 244805 426134 245125 426218
rect 244805 425898 244847 426134
rect 245083 425898 245125 426134
rect 244805 425866 245125 425898
rect 265874 426454 266194 426486
rect 265874 426218 265916 426454
rect 266152 426218 266194 426454
rect 265874 426134 266194 426218
rect 265874 425898 265916 426134
rect 266152 425898 266194 426134
rect 265874 425866 266194 425898
rect 271805 426454 272125 426486
rect 271805 426218 271847 426454
rect 272083 426218 272125 426454
rect 271805 426134 272125 426218
rect 271805 425898 271847 426134
rect 272083 425898 272125 426134
rect 271805 425866 272125 425898
rect 292874 426454 293194 426486
rect 292874 426218 292916 426454
rect 293152 426218 293194 426454
rect 292874 426134 293194 426218
rect 292874 425898 292916 426134
rect 293152 425898 293194 426134
rect 292874 425866 293194 425898
rect 298805 426454 299125 426486
rect 298805 426218 298847 426454
rect 299083 426218 299125 426454
rect 298805 426134 299125 426218
rect 298805 425898 298847 426134
rect 299083 425898 299125 426134
rect 298805 425866 299125 425898
rect 319874 426454 320194 426486
rect 319874 426218 319916 426454
rect 320152 426218 320194 426454
rect 319874 426134 320194 426218
rect 319874 425898 319916 426134
rect 320152 425898 320194 426134
rect 319874 425866 320194 425898
rect 325805 426454 326125 426486
rect 325805 426218 325847 426454
rect 326083 426218 326125 426454
rect 325805 426134 326125 426218
rect 325805 425898 325847 426134
rect 326083 425898 326125 426134
rect 325805 425866 326125 425898
rect 346874 426454 347194 426486
rect 346874 426218 346916 426454
rect 347152 426218 347194 426454
rect 346874 426134 347194 426218
rect 346874 425898 346916 426134
rect 347152 425898 347194 426134
rect 346874 425866 347194 425898
rect 352805 426454 353125 426486
rect 352805 426218 352847 426454
rect 353083 426218 353125 426454
rect 352805 426134 353125 426218
rect 352805 425898 352847 426134
rect 353083 425898 353125 426134
rect 352805 425866 353125 425898
rect 373874 426454 374194 426486
rect 373874 426218 373916 426454
rect 374152 426218 374194 426454
rect 373874 426134 374194 426218
rect 373874 425898 373916 426134
rect 374152 425898 374194 426134
rect 373874 425866 374194 425898
rect 379805 426454 380125 426486
rect 379805 426218 379847 426454
rect 380083 426218 380125 426454
rect 379805 426134 380125 426218
rect 379805 425898 379847 426134
rect 380083 425898 380125 426134
rect 379805 425866 380125 425898
rect 400874 426454 401194 426486
rect 400874 426218 400916 426454
rect 401152 426218 401194 426454
rect 400874 426134 401194 426218
rect 400874 425898 400916 426134
rect 401152 425898 401194 426134
rect 400874 425866 401194 425898
rect 406805 426454 407125 426486
rect 406805 426218 406847 426454
rect 407083 426218 407125 426454
rect 406805 426134 407125 426218
rect 406805 425898 406847 426134
rect 407083 425898 407125 426134
rect 406805 425866 407125 425898
rect 427874 426454 428194 426486
rect 427874 426218 427916 426454
rect 428152 426218 428194 426454
rect 427874 426134 428194 426218
rect 427874 425898 427916 426134
rect 428152 425898 428194 426134
rect 427874 425866 428194 425898
rect 433805 426454 434125 426486
rect 433805 426218 433847 426454
rect 434083 426218 434125 426454
rect 433805 426134 434125 426218
rect 433805 425898 433847 426134
rect 434083 425898 434125 426134
rect 433805 425866 434125 425898
rect 454874 426454 455194 426486
rect 454874 426218 454916 426454
rect 455152 426218 455194 426454
rect 454874 426134 455194 426218
rect 454874 425898 454916 426134
rect 455152 425898 455194 426134
rect 454874 425866 455194 425898
rect 460805 426454 461125 426486
rect 460805 426218 460847 426454
rect 461083 426218 461125 426454
rect 460805 426134 461125 426218
rect 460805 425898 460847 426134
rect 461083 425898 461125 426134
rect 460805 425866 461125 425898
rect 481874 426454 482194 426486
rect 481874 426218 481916 426454
rect 482152 426218 482194 426454
rect 481874 426134 482194 426218
rect 481874 425898 481916 426134
rect 482152 425898 482194 426134
rect 481874 425866 482194 425898
rect 487805 426454 488125 426486
rect 487805 426218 487847 426454
rect 488083 426218 488125 426454
rect 487805 426134 488125 426218
rect 487805 425898 487847 426134
rect 488083 425898 488125 426134
rect 487805 425866 488125 425898
rect 508874 426454 509194 426486
rect 508874 426218 508916 426454
rect 509152 426218 509194 426454
rect 508874 426134 509194 426218
rect 508874 425898 508916 426134
rect 509152 425898 509194 426134
rect 508874 425866 509194 425898
rect 514805 426454 515125 426486
rect 514805 426218 514847 426454
rect 515083 426218 515125 426454
rect 514805 426134 515125 426218
rect 514805 425898 514847 426134
rect 515083 425898 515125 426134
rect 514805 425866 515125 425898
rect 535874 426454 536194 426486
rect 535874 426218 535916 426454
rect 536152 426218 536194 426454
rect 535874 426134 536194 426218
rect 535874 425898 535916 426134
rect 536152 425898 536194 426134
rect 535874 425866 536194 425898
rect 541805 426454 542125 426486
rect 541805 426218 541847 426454
rect 542083 426218 542125 426454
rect 541805 426134 542125 426218
rect 541805 425898 541847 426134
rect 542083 425898 542125 426134
rect 541805 425866 542125 425898
rect 19794 417454 20414 419000
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 416000 20414 416898
rect 28794 418394 29414 419000
rect 28794 418158 28826 418394
rect 29062 418158 29146 418394
rect 29382 418158 29414 418394
rect 28794 418074 29414 418158
rect 28794 417838 28826 418074
rect 29062 417838 29146 418074
rect 29382 417838 29414 418074
rect 28794 416000 29414 417838
rect 37794 417454 38414 419000
rect 37794 417218 37826 417454
rect 38062 417218 38146 417454
rect 38382 417218 38414 417454
rect 37794 417134 38414 417218
rect 37794 416898 37826 417134
rect 38062 416898 38146 417134
rect 38382 416898 38414 417134
rect 37794 416000 38414 416898
rect 46794 418394 47414 419000
rect 46794 418158 46826 418394
rect 47062 418158 47146 418394
rect 47382 418158 47414 418394
rect 46794 418074 47414 418158
rect 46794 417838 46826 418074
rect 47062 417838 47146 418074
rect 47382 417838 47414 418074
rect 46794 416000 47414 417838
rect 55794 417454 56414 419000
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 416000 56414 416898
rect 64794 418394 65414 419000
rect 64794 418158 64826 418394
rect 65062 418158 65146 418394
rect 65382 418158 65414 418394
rect 64794 418074 65414 418158
rect 64794 417838 64826 418074
rect 65062 417838 65146 418074
rect 65382 417838 65414 418074
rect 64794 416000 65414 417838
rect 73794 417454 74414 419000
rect 73794 417218 73826 417454
rect 74062 417218 74146 417454
rect 74382 417218 74414 417454
rect 73794 417134 74414 417218
rect 73794 416898 73826 417134
rect 74062 416898 74146 417134
rect 74382 416898 74414 417134
rect 73794 416000 74414 416898
rect 82794 418394 83414 419000
rect 82794 418158 82826 418394
rect 83062 418158 83146 418394
rect 83382 418158 83414 418394
rect 82794 418074 83414 418158
rect 82794 417838 82826 418074
rect 83062 417838 83146 418074
rect 83382 417838 83414 418074
rect 82794 416000 83414 417838
rect 91794 417454 92414 419000
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 416000 92414 416898
rect 100794 418394 101414 419000
rect 100794 418158 100826 418394
rect 101062 418158 101146 418394
rect 101382 418158 101414 418394
rect 100794 418074 101414 418158
rect 100794 417838 100826 418074
rect 101062 417838 101146 418074
rect 101382 417838 101414 418074
rect 100794 416000 101414 417838
rect 109794 417454 110414 419000
rect 109794 417218 109826 417454
rect 110062 417218 110146 417454
rect 110382 417218 110414 417454
rect 109794 417134 110414 417218
rect 109794 416898 109826 417134
rect 110062 416898 110146 417134
rect 110382 416898 110414 417134
rect 109794 416000 110414 416898
rect 118794 418394 119414 419000
rect 118794 418158 118826 418394
rect 119062 418158 119146 418394
rect 119382 418158 119414 418394
rect 118794 418074 119414 418158
rect 118794 417838 118826 418074
rect 119062 417838 119146 418074
rect 119382 417838 119414 418074
rect 118794 416000 119414 417838
rect 127794 417454 128414 419000
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 416000 128414 416898
rect 136794 418394 137414 419000
rect 136794 418158 136826 418394
rect 137062 418158 137146 418394
rect 137382 418158 137414 418394
rect 136794 418074 137414 418158
rect 136794 417838 136826 418074
rect 137062 417838 137146 418074
rect 137382 417838 137414 418074
rect 136794 416000 137414 417838
rect 145794 417454 146414 419000
rect 145794 417218 145826 417454
rect 146062 417218 146146 417454
rect 146382 417218 146414 417454
rect 145794 417134 146414 417218
rect 145794 416898 145826 417134
rect 146062 416898 146146 417134
rect 146382 416898 146414 417134
rect 145794 416000 146414 416898
rect 154794 418394 155414 419000
rect 154794 418158 154826 418394
rect 155062 418158 155146 418394
rect 155382 418158 155414 418394
rect 154794 418074 155414 418158
rect 154794 417838 154826 418074
rect 155062 417838 155146 418074
rect 155382 417838 155414 418074
rect 154794 416000 155414 417838
rect 163794 417454 164414 419000
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 416000 164414 416898
rect 172794 418394 173414 419000
rect 172794 418158 172826 418394
rect 173062 418158 173146 418394
rect 173382 418158 173414 418394
rect 172794 418074 173414 418158
rect 172794 417838 172826 418074
rect 173062 417838 173146 418074
rect 173382 417838 173414 418074
rect 172794 416000 173414 417838
rect 181794 417454 182414 419000
rect 181794 417218 181826 417454
rect 182062 417218 182146 417454
rect 182382 417218 182414 417454
rect 181794 417134 182414 417218
rect 181794 416898 181826 417134
rect 182062 416898 182146 417134
rect 182382 416898 182414 417134
rect 181794 416000 182414 416898
rect 190794 418394 191414 419000
rect 190794 418158 190826 418394
rect 191062 418158 191146 418394
rect 191382 418158 191414 418394
rect 190794 418074 191414 418158
rect 190794 417838 190826 418074
rect 191062 417838 191146 418074
rect 191382 417838 191414 418074
rect 190794 416000 191414 417838
rect 199794 417454 200414 419000
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 416000 200414 416898
rect 208794 418394 209414 419000
rect 208794 418158 208826 418394
rect 209062 418158 209146 418394
rect 209382 418158 209414 418394
rect 208794 418074 209414 418158
rect 208794 417838 208826 418074
rect 209062 417838 209146 418074
rect 209382 417838 209414 418074
rect 208794 416000 209414 417838
rect 217794 417454 218414 419000
rect 217794 417218 217826 417454
rect 218062 417218 218146 417454
rect 218382 417218 218414 417454
rect 217794 417134 218414 417218
rect 217794 416898 217826 417134
rect 218062 416898 218146 417134
rect 218382 416898 218414 417134
rect 217794 416000 218414 416898
rect 226794 418394 227414 419000
rect 226794 418158 226826 418394
rect 227062 418158 227146 418394
rect 227382 418158 227414 418394
rect 226794 418074 227414 418158
rect 226794 417838 226826 418074
rect 227062 417838 227146 418074
rect 227382 417838 227414 418074
rect 226794 416000 227414 417838
rect 235794 417454 236414 419000
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 416000 236414 416898
rect 244794 418394 245414 419000
rect 244794 418158 244826 418394
rect 245062 418158 245146 418394
rect 245382 418158 245414 418394
rect 244794 418074 245414 418158
rect 244794 417838 244826 418074
rect 245062 417838 245146 418074
rect 245382 417838 245414 418074
rect 244794 416000 245414 417838
rect 253794 417454 254414 419000
rect 253794 417218 253826 417454
rect 254062 417218 254146 417454
rect 254382 417218 254414 417454
rect 253794 417134 254414 417218
rect 253794 416898 253826 417134
rect 254062 416898 254146 417134
rect 254382 416898 254414 417134
rect 253794 416000 254414 416898
rect 262794 418394 263414 419000
rect 262794 418158 262826 418394
rect 263062 418158 263146 418394
rect 263382 418158 263414 418394
rect 262794 418074 263414 418158
rect 262794 417838 262826 418074
rect 263062 417838 263146 418074
rect 263382 417838 263414 418074
rect 262794 416000 263414 417838
rect 271794 417454 272414 419000
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 416000 272414 416898
rect 280794 418394 281414 419000
rect 280794 418158 280826 418394
rect 281062 418158 281146 418394
rect 281382 418158 281414 418394
rect 280794 418074 281414 418158
rect 280794 417838 280826 418074
rect 281062 417838 281146 418074
rect 281382 417838 281414 418074
rect 280794 416000 281414 417838
rect 289794 417454 290414 419000
rect 289794 417218 289826 417454
rect 290062 417218 290146 417454
rect 290382 417218 290414 417454
rect 289794 417134 290414 417218
rect 289794 416898 289826 417134
rect 290062 416898 290146 417134
rect 290382 416898 290414 417134
rect 289794 416000 290414 416898
rect 298794 418394 299414 419000
rect 298794 418158 298826 418394
rect 299062 418158 299146 418394
rect 299382 418158 299414 418394
rect 298794 418074 299414 418158
rect 298794 417838 298826 418074
rect 299062 417838 299146 418074
rect 299382 417838 299414 418074
rect 298794 416000 299414 417838
rect 307794 417454 308414 419000
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 416000 308414 416898
rect 316794 418394 317414 419000
rect 316794 418158 316826 418394
rect 317062 418158 317146 418394
rect 317382 418158 317414 418394
rect 316794 418074 317414 418158
rect 316794 417838 316826 418074
rect 317062 417838 317146 418074
rect 317382 417838 317414 418074
rect 316794 416000 317414 417838
rect 325794 417454 326414 419000
rect 325794 417218 325826 417454
rect 326062 417218 326146 417454
rect 326382 417218 326414 417454
rect 325794 417134 326414 417218
rect 325794 416898 325826 417134
rect 326062 416898 326146 417134
rect 326382 416898 326414 417134
rect 325794 416000 326414 416898
rect 334794 418394 335414 419000
rect 334794 418158 334826 418394
rect 335062 418158 335146 418394
rect 335382 418158 335414 418394
rect 334794 418074 335414 418158
rect 334794 417838 334826 418074
rect 335062 417838 335146 418074
rect 335382 417838 335414 418074
rect 334794 416000 335414 417838
rect 343794 417454 344414 419000
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 416000 344414 416898
rect 352794 418394 353414 419000
rect 352794 418158 352826 418394
rect 353062 418158 353146 418394
rect 353382 418158 353414 418394
rect 352794 418074 353414 418158
rect 352794 417838 352826 418074
rect 353062 417838 353146 418074
rect 353382 417838 353414 418074
rect 352794 416000 353414 417838
rect 361794 417454 362414 419000
rect 361794 417218 361826 417454
rect 362062 417218 362146 417454
rect 362382 417218 362414 417454
rect 361794 417134 362414 417218
rect 361794 416898 361826 417134
rect 362062 416898 362146 417134
rect 362382 416898 362414 417134
rect 361794 416000 362414 416898
rect 370794 418394 371414 419000
rect 370794 418158 370826 418394
rect 371062 418158 371146 418394
rect 371382 418158 371414 418394
rect 370794 418074 371414 418158
rect 370794 417838 370826 418074
rect 371062 417838 371146 418074
rect 371382 417838 371414 418074
rect 370794 416000 371414 417838
rect 379794 417454 380414 419000
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 416000 380414 416898
rect 388794 418394 389414 419000
rect 388794 418158 388826 418394
rect 389062 418158 389146 418394
rect 389382 418158 389414 418394
rect 388794 418074 389414 418158
rect 388794 417838 388826 418074
rect 389062 417838 389146 418074
rect 389382 417838 389414 418074
rect 388794 416000 389414 417838
rect 397794 417454 398414 419000
rect 397794 417218 397826 417454
rect 398062 417218 398146 417454
rect 398382 417218 398414 417454
rect 397794 417134 398414 417218
rect 397794 416898 397826 417134
rect 398062 416898 398146 417134
rect 398382 416898 398414 417134
rect 397794 416000 398414 416898
rect 406794 418394 407414 419000
rect 406794 418158 406826 418394
rect 407062 418158 407146 418394
rect 407382 418158 407414 418394
rect 406794 418074 407414 418158
rect 406794 417838 406826 418074
rect 407062 417838 407146 418074
rect 407382 417838 407414 418074
rect 406794 416000 407414 417838
rect 415794 417454 416414 419000
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 416000 416414 416898
rect 424794 418394 425414 419000
rect 424794 418158 424826 418394
rect 425062 418158 425146 418394
rect 425382 418158 425414 418394
rect 424794 418074 425414 418158
rect 424794 417838 424826 418074
rect 425062 417838 425146 418074
rect 425382 417838 425414 418074
rect 424794 416000 425414 417838
rect 433794 417454 434414 419000
rect 433794 417218 433826 417454
rect 434062 417218 434146 417454
rect 434382 417218 434414 417454
rect 433794 417134 434414 417218
rect 433794 416898 433826 417134
rect 434062 416898 434146 417134
rect 434382 416898 434414 417134
rect 433794 416000 434414 416898
rect 442794 418394 443414 419000
rect 442794 418158 442826 418394
rect 443062 418158 443146 418394
rect 443382 418158 443414 418394
rect 442794 418074 443414 418158
rect 442794 417838 442826 418074
rect 443062 417838 443146 418074
rect 443382 417838 443414 418074
rect 442794 416000 443414 417838
rect 451794 417454 452414 419000
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 416000 452414 416898
rect 460794 418394 461414 419000
rect 460794 418158 460826 418394
rect 461062 418158 461146 418394
rect 461382 418158 461414 418394
rect 460794 418074 461414 418158
rect 460794 417838 460826 418074
rect 461062 417838 461146 418074
rect 461382 417838 461414 418074
rect 460794 416000 461414 417838
rect 469794 417454 470414 419000
rect 469794 417218 469826 417454
rect 470062 417218 470146 417454
rect 470382 417218 470414 417454
rect 469794 417134 470414 417218
rect 469794 416898 469826 417134
rect 470062 416898 470146 417134
rect 470382 416898 470414 417134
rect 469794 416000 470414 416898
rect 478794 418394 479414 419000
rect 478794 418158 478826 418394
rect 479062 418158 479146 418394
rect 479382 418158 479414 418394
rect 478794 418074 479414 418158
rect 478794 417838 478826 418074
rect 479062 417838 479146 418074
rect 479382 417838 479414 418074
rect 478794 416000 479414 417838
rect 487794 417454 488414 419000
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 416000 488414 416898
rect 496794 418394 497414 419000
rect 496794 418158 496826 418394
rect 497062 418158 497146 418394
rect 497382 418158 497414 418394
rect 496794 418074 497414 418158
rect 496794 417838 496826 418074
rect 497062 417838 497146 418074
rect 497382 417838 497414 418074
rect 496794 416000 497414 417838
rect 505794 417454 506414 419000
rect 505794 417218 505826 417454
rect 506062 417218 506146 417454
rect 506382 417218 506414 417454
rect 505794 417134 506414 417218
rect 505794 416898 505826 417134
rect 506062 416898 506146 417134
rect 506382 416898 506414 417134
rect 505794 416000 506414 416898
rect 514794 418394 515414 419000
rect 514794 418158 514826 418394
rect 515062 418158 515146 418394
rect 515382 418158 515414 418394
rect 514794 418074 515414 418158
rect 514794 417838 514826 418074
rect 515062 417838 515146 418074
rect 515382 417838 515414 418074
rect 514794 416000 515414 417838
rect 523794 417454 524414 419000
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 416000 524414 416898
rect 532794 418394 533414 419000
rect 532794 418158 532826 418394
rect 533062 418158 533146 418394
rect 533382 418158 533414 418394
rect 532794 418074 533414 418158
rect 532794 417838 532826 418074
rect 533062 417838 533146 418074
rect 533382 417838 533414 418074
rect 532794 416000 533414 417838
rect 541794 417454 542414 419000
rect 541794 417218 541826 417454
rect 542062 417218 542146 417454
rect 542382 417218 542414 417454
rect 541794 417134 542414 417218
rect 541794 416898 541826 417134
rect 542062 416898 542146 417134
rect 542382 416898 542414 417134
rect 541794 416000 542414 416898
rect 550794 418394 551414 419000
rect 550794 418158 550826 418394
rect 551062 418158 551146 418394
rect 551382 418158 551414 418394
rect 550794 418074 551414 418158
rect 550794 417838 550826 418074
rect 551062 417838 551146 418074
rect 551382 417838 551414 418074
rect 550794 416000 551414 417838
rect 559794 417454 560414 434898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 390454 11414 407898
rect 22874 408454 23194 408486
rect 22874 408218 22916 408454
rect 23152 408218 23194 408454
rect 22874 408134 23194 408218
rect 22874 407898 22916 408134
rect 23152 407898 23194 408134
rect 22874 407866 23194 407898
rect 28805 408454 29125 408486
rect 28805 408218 28847 408454
rect 29083 408218 29125 408454
rect 28805 408134 29125 408218
rect 28805 407898 28847 408134
rect 29083 407898 29125 408134
rect 28805 407866 29125 407898
rect 49874 408454 50194 408486
rect 49874 408218 49916 408454
rect 50152 408218 50194 408454
rect 49874 408134 50194 408218
rect 49874 407898 49916 408134
rect 50152 407898 50194 408134
rect 49874 407866 50194 407898
rect 55805 408454 56125 408486
rect 55805 408218 55847 408454
rect 56083 408218 56125 408454
rect 55805 408134 56125 408218
rect 55805 407898 55847 408134
rect 56083 407898 56125 408134
rect 55805 407866 56125 407898
rect 76874 408454 77194 408486
rect 76874 408218 76916 408454
rect 77152 408218 77194 408454
rect 76874 408134 77194 408218
rect 76874 407898 76916 408134
rect 77152 407898 77194 408134
rect 76874 407866 77194 407898
rect 82805 408454 83125 408486
rect 82805 408218 82847 408454
rect 83083 408218 83125 408454
rect 82805 408134 83125 408218
rect 82805 407898 82847 408134
rect 83083 407898 83125 408134
rect 82805 407866 83125 407898
rect 103874 408454 104194 408486
rect 103874 408218 103916 408454
rect 104152 408218 104194 408454
rect 103874 408134 104194 408218
rect 103874 407898 103916 408134
rect 104152 407898 104194 408134
rect 103874 407866 104194 407898
rect 109805 408454 110125 408486
rect 109805 408218 109847 408454
rect 110083 408218 110125 408454
rect 109805 408134 110125 408218
rect 109805 407898 109847 408134
rect 110083 407898 110125 408134
rect 109805 407866 110125 407898
rect 130874 408454 131194 408486
rect 130874 408218 130916 408454
rect 131152 408218 131194 408454
rect 130874 408134 131194 408218
rect 130874 407898 130916 408134
rect 131152 407898 131194 408134
rect 130874 407866 131194 407898
rect 136805 408454 137125 408486
rect 136805 408218 136847 408454
rect 137083 408218 137125 408454
rect 136805 408134 137125 408218
rect 136805 407898 136847 408134
rect 137083 407898 137125 408134
rect 136805 407866 137125 407898
rect 157874 408454 158194 408486
rect 157874 408218 157916 408454
rect 158152 408218 158194 408454
rect 157874 408134 158194 408218
rect 157874 407898 157916 408134
rect 158152 407898 158194 408134
rect 157874 407866 158194 407898
rect 163805 408454 164125 408486
rect 163805 408218 163847 408454
rect 164083 408218 164125 408454
rect 163805 408134 164125 408218
rect 163805 407898 163847 408134
rect 164083 407898 164125 408134
rect 163805 407866 164125 407898
rect 184874 408454 185194 408486
rect 184874 408218 184916 408454
rect 185152 408218 185194 408454
rect 184874 408134 185194 408218
rect 184874 407898 184916 408134
rect 185152 407898 185194 408134
rect 184874 407866 185194 407898
rect 190805 408454 191125 408486
rect 190805 408218 190847 408454
rect 191083 408218 191125 408454
rect 190805 408134 191125 408218
rect 190805 407898 190847 408134
rect 191083 407898 191125 408134
rect 190805 407866 191125 407898
rect 211874 408454 212194 408486
rect 211874 408218 211916 408454
rect 212152 408218 212194 408454
rect 211874 408134 212194 408218
rect 211874 407898 211916 408134
rect 212152 407898 212194 408134
rect 211874 407866 212194 407898
rect 217805 408454 218125 408486
rect 217805 408218 217847 408454
rect 218083 408218 218125 408454
rect 217805 408134 218125 408218
rect 217805 407898 217847 408134
rect 218083 407898 218125 408134
rect 217805 407866 218125 407898
rect 238874 408454 239194 408486
rect 238874 408218 238916 408454
rect 239152 408218 239194 408454
rect 238874 408134 239194 408218
rect 238874 407898 238916 408134
rect 239152 407898 239194 408134
rect 238874 407866 239194 407898
rect 244805 408454 245125 408486
rect 244805 408218 244847 408454
rect 245083 408218 245125 408454
rect 244805 408134 245125 408218
rect 244805 407898 244847 408134
rect 245083 407898 245125 408134
rect 244805 407866 245125 407898
rect 265874 408454 266194 408486
rect 265874 408218 265916 408454
rect 266152 408218 266194 408454
rect 265874 408134 266194 408218
rect 265874 407898 265916 408134
rect 266152 407898 266194 408134
rect 265874 407866 266194 407898
rect 271805 408454 272125 408486
rect 271805 408218 271847 408454
rect 272083 408218 272125 408454
rect 271805 408134 272125 408218
rect 271805 407898 271847 408134
rect 272083 407898 272125 408134
rect 271805 407866 272125 407898
rect 292874 408454 293194 408486
rect 292874 408218 292916 408454
rect 293152 408218 293194 408454
rect 292874 408134 293194 408218
rect 292874 407898 292916 408134
rect 293152 407898 293194 408134
rect 292874 407866 293194 407898
rect 298805 408454 299125 408486
rect 298805 408218 298847 408454
rect 299083 408218 299125 408454
rect 298805 408134 299125 408218
rect 298805 407898 298847 408134
rect 299083 407898 299125 408134
rect 298805 407866 299125 407898
rect 319874 408454 320194 408486
rect 319874 408218 319916 408454
rect 320152 408218 320194 408454
rect 319874 408134 320194 408218
rect 319874 407898 319916 408134
rect 320152 407898 320194 408134
rect 319874 407866 320194 407898
rect 325805 408454 326125 408486
rect 325805 408218 325847 408454
rect 326083 408218 326125 408454
rect 325805 408134 326125 408218
rect 325805 407898 325847 408134
rect 326083 407898 326125 408134
rect 325805 407866 326125 407898
rect 346874 408454 347194 408486
rect 346874 408218 346916 408454
rect 347152 408218 347194 408454
rect 346874 408134 347194 408218
rect 346874 407898 346916 408134
rect 347152 407898 347194 408134
rect 346874 407866 347194 407898
rect 352805 408454 353125 408486
rect 352805 408218 352847 408454
rect 353083 408218 353125 408454
rect 352805 408134 353125 408218
rect 352805 407898 352847 408134
rect 353083 407898 353125 408134
rect 352805 407866 353125 407898
rect 373874 408454 374194 408486
rect 373874 408218 373916 408454
rect 374152 408218 374194 408454
rect 373874 408134 374194 408218
rect 373874 407898 373916 408134
rect 374152 407898 374194 408134
rect 373874 407866 374194 407898
rect 379805 408454 380125 408486
rect 379805 408218 379847 408454
rect 380083 408218 380125 408454
rect 379805 408134 380125 408218
rect 379805 407898 379847 408134
rect 380083 407898 380125 408134
rect 379805 407866 380125 407898
rect 400874 408454 401194 408486
rect 400874 408218 400916 408454
rect 401152 408218 401194 408454
rect 400874 408134 401194 408218
rect 400874 407898 400916 408134
rect 401152 407898 401194 408134
rect 400874 407866 401194 407898
rect 406805 408454 407125 408486
rect 406805 408218 406847 408454
rect 407083 408218 407125 408454
rect 406805 408134 407125 408218
rect 406805 407898 406847 408134
rect 407083 407898 407125 408134
rect 406805 407866 407125 407898
rect 427874 408454 428194 408486
rect 427874 408218 427916 408454
rect 428152 408218 428194 408454
rect 427874 408134 428194 408218
rect 427874 407898 427916 408134
rect 428152 407898 428194 408134
rect 427874 407866 428194 407898
rect 433805 408454 434125 408486
rect 433805 408218 433847 408454
rect 434083 408218 434125 408454
rect 433805 408134 434125 408218
rect 433805 407898 433847 408134
rect 434083 407898 434125 408134
rect 433805 407866 434125 407898
rect 454874 408454 455194 408486
rect 454874 408218 454916 408454
rect 455152 408218 455194 408454
rect 454874 408134 455194 408218
rect 454874 407898 454916 408134
rect 455152 407898 455194 408134
rect 454874 407866 455194 407898
rect 460805 408454 461125 408486
rect 460805 408218 460847 408454
rect 461083 408218 461125 408454
rect 460805 408134 461125 408218
rect 460805 407898 460847 408134
rect 461083 407898 461125 408134
rect 460805 407866 461125 407898
rect 481874 408454 482194 408486
rect 481874 408218 481916 408454
rect 482152 408218 482194 408454
rect 481874 408134 482194 408218
rect 481874 407898 481916 408134
rect 482152 407898 482194 408134
rect 481874 407866 482194 407898
rect 487805 408454 488125 408486
rect 487805 408218 487847 408454
rect 488083 408218 488125 408454
rect 487805 408134 488125 408218
rect 487805 407898 487847 408134
rect 488083 407898 488125 408134
rect 487805 407866 488125 407898
rect 508874 408454 509194 408486
rect 508874 408218 508916 408454
rect 509152 408218 509194 408454
rect 508874 408134 509194 408218
rect 508874 407898 508916 408134
rect 509152 407898 509194 408134
rect 508874 407866 509194 407898
rect 514805 408454 515125 408486
rect 514805 408218 514847 408454
rect 515083 408218 515125 408454
rect 514805 408134 515125 408218
rect 514805 407898 514847 408134
rect 515083 407898 515125 408134
rect 514805 407866 515125 407898
rect 535874 408454 536194 408486
rect 535874 408218 535916 408454
rect 536152 408218 536194 408454
rect 535874 408134 536194 408218
rect 535874 407898 535916 408134
rect 536152 407898 536194 408134
rect 535874 407866 536194 407898
rect 541805 408454 542125 408486
rect 541805 408218 541847 408454
rect 542083 408218 542125 408454
rect 541805 408134 542125 408218
rect 541805 407898 541847 408134
rect 542083 407898 542125 408134
rect 541805 407866 542125 407898
rect 19910 399454 20230 399486
rect 19910 399218 19952 399454
rect 20188 399218 20230 399454
rect 19910 399134 20230 399218
rect 19910 398898 19952 399134
rect 20188 398898 20230 399134
rect 19910 398866 20230 398898
rect 25840 399454 26160 399486
rect 25840 399218 25882 399454
rect 26118 399218 26160 399454
rect 25840 399134 26160 399218
rect 25840 398898 25882 399134
rect 26118 398898 26160 399134
rect 25840 398866 26160 398898
rect 31771 399454 32091 399486
rect 31771 399218 31813 399454
rect 32049 399218 32091 399454
rect 31771 399134 32091 399218
rect 31771 398898 31813 399134
rect 32049 398898 32091 399134
rect 31771 398866 32091 398898
rect 46910 399454 47230 399486
rect 46910 399218 46952 399454
rect 47188 399218 47230 399454
rect 46910 399134 47230 399218
rect 46910 398898 46952 399134
rect 47188 398898 47230 399134
rect 46910 398866 47230 398898
rect 52840 399454 53160 399486
rect 52840 399218 52882 399454
rect 53118 399218 53160 399454
rect 52840 399134 53160 399218
rect 52840 398898 52882 399134
rect 53118 398898 53160 399134
rect 52840 398866 53160 398898
rect 58771 399454 59091 399486
rect 58771 399218 58813 399454
rect 59049 399218 59091 399454
rect 58771 399134 59091 399218
rect 58771 398898 58813 399134
rect 59049 398898 59091 399134
rect 58771 398866 59091 398898
rect 73910 399454 74230 399486
rect 73910 399218 73952 399454
rect 74188 399218 74230 399454
rect 73910 399134 74230 399218
rect 73910 398898 73952 399134
rect 74188 398898 74230 399134
rect 73910 398866 74230 398898
rect 79840 399454 80160 399486
rect 79840 399218 79882 399454
rect 80118 399218 80160 399454
rect 79840 399134 80160 399218
rect 79840 398898 79882 399134
rect 80118 398898 80160 399134
rect 79840 398866 80160 398898
rect 85771 399454 86091 399486
rect 85771 399218 85813 399454
rect 86049 399218 86091 399454
rect 85771 399134 86091 399218
rect 85771 398898 85813 399134
rect 86049 398898 86091 399134
rect 85771 398866 86091 398898
rect 100910 399454 101230 399486
rect 100910 399218 100952 399454
rect 101188 399218 101230 399454
rect 100910 399134 101230 399218
rect 100910 398898 100952 399134
rect 101188 398898 101230 399134
rect 100910 398866 101230 398898
rect 106840 399454 107160 399486
rect 106840 399218 106882 399454
rect 107118 399218 107160 399454
rect 106840 399134 107160 399218
rect 106840 398898 106882 399134
rect 107118 398898 107160 399134
rect 106840 398866 107160 398898
rect 112771 399454 113091 399486
rect 112771 399218 112813 399454
rect 113049 399218 113091 399454
rect 112771 399134 113091 399218
rect 112771 398898 112813 399134
rect 113049 398898 113091 399134
rect 112771 398866 113091 398898
rect 127910 399454 128230 399486
rect 127910 399218 127952 399454
rect 128188 399218 128230 399454
rect 127910 399134 128230 399218
rect 127910 398898 127952 399134
rect 128188 398898 128230 399134
rect 127910 398866 128230 398898
rect 133840 399454 134160 399486
rect 133840 399218 133882 399454
rect 134118 399218 134160 399454
rect 133840 399134 134160 399218
rect 133840 398898 133882 399134
rect 134118 398898 134160 399134
rect 133840 398866 134160 398898
rect 139771 399454 140091 399486
rect 139771 399218 139813 399454
rect 140049 399218 140091 399454
rect 139771 399134 140091 399218
rect 139771 398898 139813 399134
rect 140049 398898 140091 399134
rect 139771 398866 140091 398898
rect 154910 399454 155230 399486
rect 154910 399218 154952 399454
rect 155188 399218 155230 399454
rect 154910 399134 155230 399218
rect 154910 398898 154952 399134
rect 155188 398898 155230 399134
rect 154910 398866 155230 398898
rect 160840 399454 161160 399486
rect 160840 399218 160882 399454
rect 161118 399218 161160 399454
rect 160840 399134 161160 399218
rect 160840 398898 160882 399134
rect 161118 398898 161160 399134
rect 160840 398866 161160 398898
rect 166771 399454 167091 399486
rect 166771 399218 166813 399454
rect 167049 399218 167091 399454
rect 166771 399134 167091 399218
rect 166771 398898 166813 399134
rect 167049 398898 167091 399134
rect 166771 398866 167091 398898
rect 181910 399454 182230 399486
rect 181910 399218 181952 399454
rect 182188 399218 182230 399454
rect 181910 399134 182230 399218
rect 181910 398898 181952 399134
rect 182188 398898 182230 399134
rect 181910 398866 182230 398898
rect 187840 399454 188160 399486
rect 187840 399218 187882 399454
rect 188118 399218 188160 399454
rect 187840 399134 188160 399218
rect 187840 398898 187882 399134
rect 188118 398898 188160 399134
rect 187840 398866 188160 398898
rect 193771 399454 194091 399486
rect 193771 399218 193813 399454
rect 194049 399218 194091 399454
rect 193771 399134 194091 399218
rect 193771 398898 193813 399134
rect 194049 398898 194091 399134
rect 193771 398866 194091 398898
rect 208910 399454 209230 399486
rect 208910 399218 208952 399454
rect 209188 399218 209230 399454
rect 208910 399134 209230 399218
rect 208910 398898 208952 399134
rect 209188 398898 209230 399134
rect 208910 398866 209230 398898
rect 214840 399454 215160 399486
rect 214840 399218 214882 399454
rect 215118 399218 215160 399454
rect 214840 399134 215160 399218
rect 214840 398898 214882 399134
rect 215118 398898 215160 399134
rect 214840 398866 215160 398898
rect 220771 399454 221091 399486
rect 220771 399218 220813 399454
rect 221049 399218 221091 399454
rect 220771 399134 221091 399218
rect 220771 398898 220813 399134
rect 221049 398898 221091 399134
rect 220771 398866 221091 398898
rect 235910 399454 236230 399486
rect 235910 399218 235952 399454
rect 236188 399218 236230 399454
rect 235910 399134 236230 399218
rect 235910 398898 235952 399134
rect 236188 398898 236230 399134
rect 235910 398866 236230 398898
rect 241840 399454 242160 399486
rect 241840 399218 241882 399454
rect 242118 399218 242160 399454
rect 241840 399134 242160 399218
rect 241840 398898 241882 399134
rect 242118 398898 242160 399134
rect 241840 398866 242160 398898
rect 247771 399454 248091 399486
rect 247771 399218 247813 399454
rect 248049 399218 248091 399454
rect 247771 399134 248091 399218
rect 247771 398898 247813 399134
rect 248049 398898 248091 399134
rect 247771 398866 248091 398898
rect 262910 399454 263230 399486
rect 262910 399218 262952 399454
rect 263188 399218 263230 399454
rect 262910 399134 263230 399218
rect 262910 398898 262952 399134
rect 263188 398898 263230 399134
rect 262910 398866 263230 398898
rect 268840 399454 269160 399486
rect 268840 399218 268882 399454
rect 269118 399218 269160 399454
rect 268840 399134 269160 399218
rect 268840 398898 268882 399134
rect 269118 398898 269160 399134
rect 268840 398866 269160 398898
rect 274771 399454 275091 399486
rect 274771 399218 274813 399454
rect 275049 399218 275091 399454
rect 274771 399134 275091 399218
rect 274771 398898 274813 399134
rect 275049 398898 275091 399134
rect 274771 398866 275091 398898
rect 289910 399454 290230 399486
rect 289910 399218 289952 399454
rect 290188 399218 290230 399454
rect 289910 399134 290230 399218
rect 289910 398898 289952 399134
rect 290188 398898 290230 399134
rect 289910 398866 290230 398898
rect 295840 399454 296160 399486
rect 295840 399218 295882 399454
rect 296118 399218 296160 399454
rect 295840 399134 296160 399218
rect 295840 398898 295882 399134
rect 296118 398898 296160 399134
rect 295840 398866 296160 398898
rect 301771 399454 302091 399486
rect 301771 399218 301813 399454
rect 302049 399218 302091 399454
rect 301771 399134 302091 399218
rect 301771 398898 301813 399134
rect 302049 398898 302091 399134
rect 301771 398866 302091 398898
rect 316910 399454 317230 399486
rect 316910 399218 316952 399454
rect 317188 399218 317230 399454
rect 316910 399134 317230 399218
rect 316910 398898 316952 399134
rect 317188 398898 317230 399134
rect 316910 398866 317230 398898
rect 322840 399454 323160 399486
rect 322840 399218 322882 399454
rect 323118 399218 323160 399454
rect 322840 399134 323160 399218
rect 322840 398898 322882 399134
rect 323118 398898 323160 399134
rect 322840 398866 323160 398898
rect 328771 399454 329091 399486
rect 328771 399218 328813 399454
rect 329049 399218 329091 399454
rect 328771 399134 329091 399218
rect 328771 398898 328813 399134
rect 329049 398898 329091 399134
rect 328771 398866 329091 398898
rect 343910 399454 344230 399486
rect 343910 399218 343952 399454
rect 344188 399218 344230 399454
rect 343910 399134 344230 399218
rect 343910 398898 343952 399134
rect 344188 398898 344230 399134
rect 343910 398866 344230 398898
rect 349840 399454 350160 399486
rect 349840 399218 349882 399454
rect 350118 399218 350160 399454
rect 349840 399134 350160 399218
rect 349840 398898 349882 399134
rect 350118 398898 350160 399134
rect 349840 398866 350160 398898
rect 355771 399454 356091 399486
rect 355771 399218 355813 399454
rect 356049 399218 356091 399454
rect 355771 399134 356091 399218
rect 355771 398898 355813 399134
rect 356049 398898 356091 399134
rect 355771 398866 356091 398898
rect 370910 399454 371230 399486
rect 370910 399218 370952 399454
rect 371188 399218 371230 399454
rect 370910 399134 371230 399218
rect 370910 398898 370952 399134
rect 371188 398898 371230 399134
rect 370910 398866 371230 398898
rect 376840 399454 377160 399486
rect 376840 399218 376882 399454
rect 377118 399218 377160 399454
rect 376840 399134 377160 399218
rect 376840 398898 376882 399134
rect 377118 398898 377160 399134
rect 376840 398866 377160 398898
rect 382771 399454 383091 399486
rect 382771 399218 382813 399454
rect 383049 399218 383091 399454
rect 382771 399134 383091 399218
rect 382771 398898 382813 399134
rect 383049 398898 383091 399134
rect 382771 398866 383091 398898
rect 397910 399454 398230 399486
rect 397910 399218 397952 399454
rect 398188 399218 398230 399454
rect 397910 399134 398230 399218
rect 397910 398898 397952 399134
rect 398188 398898 398230 399134
rect 397910 398866 398230 398898
rect 403840 399454 404160 399486
rect 403840 399218 403882 399454
rect 404118 399218 404160 399454
rect 403840 399134 404160 399218
rect 403840 398898 403882 399134
rect 404118 398898 404160 399134
rect 403840 398866 404160 398898
rect 409771 399454 410091 399486
rect 409771 399218 409813 399454
rect 410049 399218 410091 399454
rect 409771 399134 410091 399218
rect 409771 398898 409813 399134
rect 410049 398898 410091 399134
rect 409771 398866 410091 398898
rect 424910 399454 425230 399486
rect 424910 399218 424952 399454
rect 425188 399218 425230 399454
rect 424910 399134 425230 399218
rect 424910 398898 424952 399134
rect 425188 398898 425230 399134
rect 424910 398866 425230 398898
rect 430840 399454 431160 399486
rect 430840 399218 430882 399454
rect 431118 399218 431160 399454
rect 430840 399134 431160 399218
rect 430840 398898 430882 399134
rect 431118 398898 431160 399134
rect 430840 398866 431160 398898
rect 436771 399454 437091 399486
rect 436771 399218 436813 399454
rect 437049 399218 437091 399454
rect 436771 399134 437091 399218
rect 436771 398898 436813 399134
rect 437049 398898 437091 399134
rect 436771 398866 437091 398898
rect 451910 399454 452230 399486
rect 451910 399218 451952 399454
rect 452188 399218 452230 399454
rect 451910 399134 452230 399218
rect 451910 398898 451952 399134
rect 452188 398898 452230 399134
rect 451910 398866 452230 398898
rect 457840 399454 458160 399486
rect 457840 399218 457882 399454
rect 458118 399218 458160 399454
rect 457840 399134 458160 399218
rect 457840 398898 457882 399134
rect 458118 398898 458160 399134
rect 457840 398866 458160 398898
rect 463771 399454 464091 399486
rect 463771 399218 463813 399454
rect 464049 399218 464091 399454
rect 463771 399134 464091 399218
rect 463771 398898 463813 399134
rect 464049 398898 464091 399134
rect 463771 398866 464091 398898
rect 478910 399454 479230 399486
rect 478910 399218 478952 399454
rect 479188 399218 479230 399454
rect 478910 399134 479230 399218
rect 478910 398898 478952 399134
rect 479188 398898 479230 399134
rect 478910 398866 479230 398898
rect 484840 399454 485160 399486
rect 484840 399218 484882 399454
rect 485118 399218 485160 399454
rect 484840 399134 485160 399218
rect 484840 398898 484882 399134
rect 485118 398898 485160 399134
rect 484840 398866 485160 398898
rect 490771 399454 491091 399486
rect 490771 399218 490813 399454
rect 491049 399218 491091 399454
rect 490771 399134 491091 399218
rect 490771 398898 490813 399134
rect 491049 398898 491091 399134
rect 490771 398866 491091 398898
rect 505910 399454 506230 399486
rect 505910 399218 505952 399454
rect 506188 399218 506230 399454
rect 505910 399134 506230 399218
rect 505910 398898 505952 399134
rect 506188 398898 506230 399134
rect 505910 398866 506230 398898
rect 511840 399454 512160 399486
rect 511840 399218 511882 399454
rect 512118 399218 512160 399454
rect 511840 399134 512160 399218
rect 511840 398898 511882 399134
rect 512118 398898 512160 399134
rect 511840 398866 512160 398898
rect 517771 399454 518091 399486
rect 517771 399218 517813 399454
rect 518049 399218 518091 399454
rect 517771 399134 518091 399218
rect 517771 398898 517813 399134
rect 518049 398898 518091 399134
rect 517771 398866 518091 398898
rect 532910 399454 533230 399486
rect 532910 399218 532952 399454
rect 533188 399218 533230 399454
rect 532910 399134 533230 399218
rect 532910 398898 532952 399134
rect 533188 398898 533230 399134
rect 532910 398866 533230 398898
rect 538840 399454 539160 399486
rect 538840 399218 538882 399454
rect 539118 399218 539160 399454
rect 538840 399134 539160 399218
rect 538840 398898 538882 399134
rect 539118 398898 539160 399134
rect 538840 398866 539160 398898
rect 544771 399454 545091 399486
rect 544771 399218 544813 399454
rect 545049 399218 545091 399454
rect 544771 399134 545091 399218
rect 544771 398898 544813 399134
rect 545049 398898 545091 399134
rect 544771 398866 545091 398898
rect 559794 399454 560414 416898
rect 559794 399218 559826 399454
rect 560062 399218 560146 399454
rect 560382 399218 560414 399454
rect 559794 399134 560414 399218
rect 559794 398898 559826 399134
rect 560062 398898 560146 399134
rect 560382 398898 560414 399134
rect 10794 390218 10826 390454
rect 11062 390218 11146 390454
rect 11382 390218 11414 390454
rect 10794 390134 11414 390218
rect 10794 389898 10826 390134
rect 11062 389898 11146 390134
rect 11382 389898 11414 390134
rect 10794 372454 11414 389898
rect 19794 391394 20414 392000
rect 19794 391158 19826 391394
rect 20062 391158 20146 391394
rect 20382 391158 20414 391394
rect 19794 391074 20414 391158
rect 19794 390838 19826 391074
rect 20062 390838 20146 391074
rect 20382 390838 20414 391074
rect 19794 389000 20414 390838
rect 28794 390454 29414 392000
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 389000 29414 389898
rect 37794 391394 38414 392000
rect 37794 391158 37826 391394
rect 38062 391158 38146 391394
rect 38382 391158 38414 391394
rect 37794 391074 38414 391158
rect 37794 390838 37826 391074
rect 38062 390838 38146 391074
rect 38382 390838 38414 391074
rect 37794 389000 38414 390838
rect 46794 390454 47414 392000
rect 46794 390218 46826 390454
rect 47062 390218 47146 390454
rect 47382 390218 47414 390454
rect 46794 390134 47414 390218
rect 46794 389898 46826 390134
rect 47062 389898 47146 390134
rect 47382 389898 47414 390134
rect 46794 389000 47414 389898
rect 55794 391394 56414 392000
rect 55794 391158 55826 391394
rect 56062 391158 56146 391394
rect 56382 391158 56414 391394
rect 55794 391074 56414 391158
rect 55794 390838 55826 391074
rect 56062 390838 56146 391074
rect 56382 390838 56414 391074
rect 55794 389000 56414 390838
rect 64794 390454 65414 392000
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 389000 65414 389898
rect 73794 391394 74414 392000
rect 73794 391158 73826 391394
rect 74062 391158 74146 391394
rect 74382 391158 74414 391394
rect 73794 391074 74414 391158
rect 73794 390838 73826 391074
rect 74062 390838 74146 391074
rect 74382 390838 74414 391074
rect 73794 389000 74414 390838
rect 82794 390454 83414 392000
rect 82794 390218 82826 390454
rect 83062 390218 83146 390454
rect 83382 390218 83414 390454
rect 82794 390134 83414 390218
rect 82794 389898 82826 390134
rect 83062 389898 83146 390134
rect 83382 389898 83414 390134
rect 82794 389000 83414 389898
rect 91794 391394 92414 392000
rect 91794 391158 91826 391394
rect 92062 391158 92146 391394
rect 92382 391158 92414 391394
rect 91794 391074 92414 391158
rect 91794 390838 91826 391074
rect 92062 390838 92146 391074
rect 92382 390838 92414 391074
rect 91794 389000 92414 390838
rect 100794 390454 101414 392000
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 389000 101414 389898
rect 109794 391394 110414 392000
rect 109794 391158 109826 391394
rect 110062 391158 110146 391394
rect 110382 391158 110414 391394
rect 109794 391074 110414 391158
rect 109794 390838 109826 391074
rect 110062 390838 110146 391074
rect 110382 390838 110414 391074
rect 109794 389000 110414 390838
rect 118794 390454 119414 392000
rect 118794 390218 118826 390454
rect 119062 390218 119146 390454
rect 119382 390218 119414 390454
rect 118794 390134 119414 390218
rect 118794 389898 118826 390134
rect 119062 389898 119146 390134
rect 119382 389898 119414 390134
rect 118794 389000 119414 389898
rect 127794 391394 128414 392000
rect 127794 391158 127826 391394
rect 128062 391158 128146 391394
rect 128382 391158 128414 391394
rect 127794 391074 128414 391158
rect 127794 390838 127826 391074
rect 128062 390838 128146 391074
rect 128382 390838 128414 391074
rect 127794 389000 128414 390838
rect 136794 390454 137414 392000
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 389000 137414 389898
rect 145794 391394 146414 392000
rect 145794 391158 145826 391394
rect 146062 391158 146146 391394
rect 146382 391158 146414 391394
rect 145794 391074 146414 391158
rect 145794 390838 145826 391074
rect 146062 390838 146146 391074
rect 146382 390838 146414 391074
rect 145794 389000 146414 390838
rect 154794 390454 155414 392000
rect 154794 390218 154826 390454
rect 155062 390218 155146 390454
rect 155382 390218 155414 390454
rect 154794 390134 155414 390218
rect 154794 389898 154826 390134
rect 155062 389898 155146 390134
rect 155382 389898 155414 390134
rect 154794 389000 155414 389898
rect 163794 391394 164414 392000
rect 163794 391158 163826 391394
rect 164062 391158 164146 391394
rect 164382 391158 164414 391394
rect 163794 391074 164414 391158
rect 163794 390838 163826 391074
rect 164062 390838 164146 391074
rect 164382 390838 164414 391074
rect 163794 389000 164414 390838
rect 172794 390454 173414 392000
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 389000 173414 389898
rect 181794 391394 182414 392000
rect 181794 391158 181826 391394
rect 182062 391158 182146 391394
rect 182382 391158 182414 391394
rect 181794 391074 182414 391158
rect 181794 390838 181826 391074
rect 182062 390838 182146 391074
rect 182382 390838 182414 391074
rect 181794 389000 182414 390838
rect 190794 390454 191414 392000
rect 190794 390218 190826 390454
rect 191062 390218 191146 390454
rect 191382 390218 191414 390454
rect 190794 390134 191414 390218
rect 190794 389898 190826 390134
rect 191062 389898 191146 390134
rect 191382 389898 191414 390134
rect 190794 389000 191414 389898
rect 199794 391394 200414 392000
rect 199794 391158 199826 391394
rect 200062 391158 200146 391394
rect 200382 391158 200414 391394
rect 199794 391074 200414 391158
rect 199794 390838 199826 391074
rect 200062 390838 200146 391074
rect 200382 390838 200414 391074
rect 199794 389000 200414 390838
rect 208794 390454 209414 392000
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 389000 209414 389898
rect 217794 391394 218414 392000
rect 217794 391158 217826 391394
rect 218062 391158 218146 391394
rect 218382 391158 218414 391394
rect 217794 391074 218414 391158
rect 217794 390838 217826 391074
rect 218062 390838 218146 391074
rect 218382 390838 218414 391074
rect 217794 389000 218414 390838
rect 226794 390454 227414 392000
rect 226794 390218 226826 390454
rect 227062 390218 227146 390454
rect 227382 390218 227414 390454
rect 226794 390134 227414 390218
rect 226794 389898 226826 390134
rect 227062 389898 227146 390134
rect 227382 389898 227414 390134
rect 226794 389000 227414 389898
rect 235794 391394 236414 392000
rect 235794 391158 235826 391394
rect 236062 391158 236146 391394
rect 236382 391158 236414 391394
rect 235794 391074 236414 391158
rect 235794 390838 235826 391074
rect 236062 390838 236146 391074
rect 236382 390838 236414 391074
rect 235794 389000 236414 390838
rect 244794 390454 245414 392000
rect 244794 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 245414 390454
rect 244794 390134 245414 390218
rect 244794 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 245414 390134
rect 244794 389000 245414 389898
rect 253794 391394 254414 392000
rect 253794 391158 253826 391394
rect 254062 391158 254146 391394
rect 254382 391158 254414 391394
rect 253794 391074 254414 391158
rect 253794 390838 253826 391074
rect 254062 390838 254146 391074
rect 254382 390838 254414 391074
rect 253794 389000 254414 390838
rect 262794 390454 263414 392000
rect 262794 390218 262826 390454
rect 263062 390218 263146 390454
rect 263382 390218 263414 390454
rect 262794 390134 263414 390218
rect 262794 389898 262826 390134
rect 263062 389898 263146 390134
rect 263382 389898 263414 390134
rect 262794 389000 263414 389898
rect 271794 391394 272414 392000
rect 271794 391158 271826 391394
rect 272062 391158 272146 391394
rect 272382 391158 272414 391394
rect 271794 391074 272414 391158
rect 271794 390838 271826 391074
rect 272062 390838 272146 391074
rect 272382 390838 272414 391074
rect 271794 389000 272414 390838
rect 280794 390454 281414 392000
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 389000 281414 389898
rect 289794 391394 290414 392000
rect 289794 391158 289826 391394
rect 290062 391158 290146 391394
rect 290382 391158 290414 391394
rect 289794 391074 290414 391158
rect 289794 390838 289826 391074
rect 290062 390838 290146 391074
rect 290382 390838 290414 391074
rect 289794 389000 290414 390838
rect 298794 390454 299414 392000
rect 298794 390218 298826 390454
rect 299062 390218 299146 390454
rect 299382 390218 299414 390454
rect 298794 390134 299414 390218
rect 298794 389898 298826 390134
rect 299062 389898 299146 390134
rect 299382 389898 299414 390134
rect 298794 389000 299414 389898
rect 307794 391394 308414 392000
rect 307794 391158 307826 391394
rect 308062 391158 308146 391394
rect 308382 391158 308414 391394
rect 307794 391074 308414 391158
rect 307794 390838 307826 391074
rect 308062 390838 308146 391074
rect 308382 390838 308414 391074
rect 307794 389000 308414 390838
rect 316794 390454 317414 392000
rect 316794 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 317414 390454
rect 316794 390134 317414 390218
rect 316794 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 317414 390134
rect 316794 389000 317414 389898
rect 325794 391394 326414 392000
rect 325794 391158 325826 391394
rect 326062 391158 326146 391394
rect 326382 391158 326414 391394
rect 325794 391074 326414 391158
rect 325794 390838 325826 391074
rect 326062 390838 326146 391074
rect 326382 390838 326414 391074
rect 325794 389000 326414 390838
rect 334794 390454 335414 392000
rect 334794 390218 334826 390454
rect 335062 390218 335146 390454
rect 335382 390218 335414 390454
rect 334794 390134 335414 390218
rect 334794 389898 334826 390134
rect 335062 389898 335146 390134
rect 335382 389898 335414 390134
rect 334794 389000 335414 389898
rect 343794 391394 344414 392000
rect 343794 391158 343826 391394
rect 344062 391158 344146 391394
rect 344382 391158 344414 391394
rect 343794 391074 344414 391158
rect 343794 390838 343826 391074
rect 344062 390838 344146 391074
rect 344382 390838 344414 391074
rect 343794 389000 344414 390838
rect 352794 390454 353414 392000
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 389000 353414 389898
rect 361794 391394 362414 392000
rect 361794 391158 361826 391394
rect 362062 391158 362146 391394
rect 362382 391158 362414 391394
rect 361794 391074 362414 391158
rect 361794 390838 361826 391074
rect 362062 390838 362146 391074
rect 362382 390838 362414 391074
rect 361794 389000 362414 390838
rect 370794 390454 371414 392000
rect 370794 390218 370826 390454
rect 371062 390218 371146 390454
rect 371382 390218 371414 390454
rect 370794 390134 371414 390218
rect 370794 389898 370826 390134
rect 371062 389898 371146 390134
rect 371382 389898 371414 390134
rect 370794 389000 371414 389898
rect 379794 391394 380414 392000
rect 379794 391158 379826 391394
rect 380062 391158 380146 391394
rect 380382 391158 380414 391394
rect 379794 391074 380414 391158
rect 379794 390838 379826 391074
rect 380062 390838 380146 391074
rect 380382 390838 380414 391074
rect 379794 389000 380414 390838
rect 388794 390454 389414 392000
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 389000 389414 389898
rect 397794 391394 398414 392000
rect 397794 391158 397826 391394
rect 398062 391158 398146 391394
rect 398382 391158 398414 391394
rect 397794 391074 398414 391158
rect 397794 390838 397826 391074
rect 398062 390838 398146 391074
rect 398382 390838 398414 391074
rect 397794 389000 398414 390838
rect 406794 390454 407414 392000
rect 406794 390218 406826 390454
rect 407062 390218 407146 390454
rect 407382 390218 407414 390454
rect 406794 390134 407414 390218
rect 406794 389898 406826 390134
rect 407062 389898 407146 390134
rect 407382 389898 407414 390134
rect 406794 389000 407414 389898
rect 415794 391394 416414 392000
rect 415794 391158 415826 391394
rect 416062 391158 416146 391394
rect 416382 391158 416414 391394
rect 415794 391074 416414 391158
rect 415794 390838 415826 391074
rect 416062 390838 416146 391074
rect 416382 390838 416414 391074
rect 415794 389000 416414 390838
rect 424794 390454 425414 392000
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 389000 425414 389898
rect 433794 391394 434414 392000
rect 433794 391158 433826 391394
rect 434062 391158 434146 391394
rect 434382 391158 434414 391394
rect 433794 391074 434414 391158
rect 433794 390838 433826 391074
rect 434062 390838 434146 391074
rect 434382 390838 434414 391074
rect 433794 389000 434414 390838
rect 442794 390454 443414 392000
rect 442794 390218 442826 390454
rect 443062 390218 443146 390454
rect 443382 390218 443414 390454
rect 442794 390134 443414 390218
rect 442794 389898 442826 390134
rect 443062 389898 443146 390134
rect 443382 389898 443414 390134
rect 442794 389000 443414 389898
rect 451794 391394 452414 392000
rect 451794 391158 451826 391394
rect 452062 391158 452146 391394
rect 452382 391158 452414 391394
rect 451794 391074 452414 391158
rect 451794 390838 451826 391074
rect 452062 390838 452146 391074
rect 452382 390838 452414 391074
rect 451794 389000 452414 390838
rect 460794 390454 461414 392000
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 389000 461414 389898
rect 469794 391394 470414 392000
rect 469794 391158 469826 391394
rect 470062 391158 470146 391394
rect 470382 391158 470414 391394
rect 469794 391074 470414 391158
rect 469794 390838 469826 391074
rect 470062 390838 470146 391074
rect 470382 390838 470414 391074
rect 469794 389000 470414 390838
rect 478794 390454 479414 392000
rect 478794 390218 478826 390454
rect 479062 390218 479146 390454
rect 479382 390218 479414 390454
rect 478794 390134 479414 390218
rect 478794 389898 478826 390134
rect 479062 389898 479146 390134
rect 479382 389898 479414 390134
rect 478794 389000 479414 389898
rect 487794 391394 488414 392000
rect 487794 391158 487826 391394
rect 488062 391158 488146 391394
rect 488382 391158 488414 391394
rect 487794 391074 488414 391158
rect 487794 390838 487826 391074
rect 488062 390838 488146 391074
rect 488382 390838 488414 391074
rect 487794 389000 488414 390838
rect 496794 390454 497414 392000
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 389000 497414 389898
rect 505794 391394 506414 392000
rect 505794 391158 505826 391394
rect 506062 391158 506146 391394
rect 506382 391158 506414 391394
rect 505794 391074 506414 391158
rect 505794 390838 505826 391074
rect 506062 390838 506146 391074
rect 506382 390838 506414 391074
rect 505794 389000 506414 390838
rect 514794 390454 515414 392000
rect 514794 390218 514826 390454
rect 515062 390218 515146 390454
rect 515382 390218 515414 390454
rect 514794 390134 515414 390218
rect 514794 389898 514826 390134
rect 515062 389898 515146 390134
rect 515382 389898 515414 390134
rect 514794 389000 515414 389898
rect 523794 391394 524414 392000
rect 523794 391158 523826 391394
rect 524062 391158 524146 391394
rect 524382 391158 524414 391394
rect 523794 391074 524414 391158
rect 523794 390838 523826 391074
rect 524062 390838 524146 391074
rect 524382 390838 524414 391074
rect 523794 389000 524414 390838
rect 532794 390454 533414 392000
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 389000 533414 389898
rect 541794 391394 542414 392000
rect 541794 391158 541826 391394
rect 542062 391158 542146 391394
rect 542382 391158 542414 391394
rect 541794 391074 542414 391158
rect 541794 390838 541826 391074
rect 542062 390838 542146 391074
rect 542382 390838 542414 391074
rect 541794 389000 542414 390838
rect 550794 390454 551414 392000
rect 550794 390218 550826 390454
rect 551062 390218 551146 390454
rect 551382 390218 551414 390454
rect 550794 390134 551414 390218
rect 550794 389898 550826 390134
rect 551062 389898 551146 390134
rect 551382 389898 551414 390134
rect 550794 389000 551414 389898
rect 19910 381454 20230 381486
rect 19910 381218 19952 381454
rect 20188 381218 20230 381454
rect 19910 381134 20230 381218
rect 19910 380898 19952 381134
rect 20188 380898 20230 381134
rect 19910 380866 20230 380898
rect 25840 381454 26160 381486
rect 25840 381218 25882 381454
rect 26118 381218 26160 381454
rect 25840 381134 26160 381218
rect 25840 380898 25882 381134
rect 26118 380898 26160 381134
rect 25840 380866 26160 380898
rect 31771 381454 32091 381486
rect 31771 381218 31813 381454
rect 32049 381218 32091 381454
rect 31771 381134 32091 381218
rect 31771 380898 31813 381134
rect 32049 380898 32091 381134
rect 31771 380866 32091 380898
rect 46910 381454 47230 381486
rect 46910 381218 46952 381454
rect 47188 381218 47230 381454
rect 46910 381134 47230 381218
rect 46910 380898 46952 381134
rect 47188 380898 47230 381134
rect 46910 380866 47230 380898
rect 52840 381454 53160 381486
rect 52840 381218 52882 381454
rect 53118 381218 53160 381454
rect 52840 381134 53160 381218
rect 52840 380898 52882 381134
rect 53118 380898 53160 381134
rect 52840 380866 53160 380898
rect 58771 381454 59091 381486
rect 58771 381218 58813 381454
rect 59049 381218 59091 381454
rect 58771 381134 59091 381218
rect 58771 380898 58813 381134
rect 59049 380898 59091 381134
rect 58771 380866 59091 380898
rect 73910 381454 74230 381486
rect 73910 381218 73952 381454
rect 74188 381218 74230 381454
rect 73910 381134 74230 381218
rect 73910 380898 73952 381134
rect 74188 380898 74230 381134
rect 73910 380866 74230 380898
rect 79840 381454 80160 381486
rect 79840 381218 79882 381454
rect 80118 381218 80160 381454
rect 79840 381134 80160 381218
rect 79840 380898 79882 381134
rect 80118 380898 80160 381134
rect 79840 380866 80160 380898
rect 85771 381454 86091 381486
rect 85771 381218 85813 381454
rect 86049 381218 86091 381454
rect 85771 381134 86091 381218
rect 85771 380898 85813 381134
rect 86049 380898 86091 381134
rect 85771 380866 86091 380898
rect 100910 381454 101230 381486
rect 100910 381218 100952 381454
rect 101188 381218 101230 381454
rect 100910 381134 101230 381218
rect 100910 380898 100952 381134
rect 101188 380898 101230 381134
rect 100910 380866 101230 380898
rect 106840 381454 107160 381486
rect 106840 381218 106882 381454
rect 107118 381218 107160 381454
rect 106840 381134 107160 381218
rect 106840 380898 106882 381134
rect 107118 380898 107160 381134
rect 106840 380866 107160 380898
rect 112771 381454 113091 381486
rect 112771 381218 112813 381454
rect 113049 381218 113091 381454
rect 112771 381134 113091 381218
rect 112771 380898 112813 381134
rect 113049 380898 113091 381134
rect 112771 380866 113091 380898
rect 127910 381454 128230 381486
rect 127910 381218 127952 381454
rect 128188 381218 128230 381454
rect 127910 381134 128230 381218
rect 127910 380898 127952 381134
rect 128188 380898 128230 381134
rect 127910 380866 128230 380898
rect 133840 381454 134160 381486
rect 133840 381218 133882 381454
rect 134118 381218 134160 381454
rect 133840 381134 134160 381218
rect 133840 380898 133882 381134
rect 134118 380898 134160 381134
rect 133840 380866 134160 380898
rect 139771 381454 140091 381486
rect 139771 381218 139813 381454
rect 140049 381218 140091 381454
rect 139771 381134 140091 381218
rect 139771 380898 139813 381134
rect 140049 380898 140091 381134
rect 139771 380866 140091 380898
rect 154910 381454 155230 381486
rect 154910 381218 154952 381454
rect 155188 381218 155230 381454
rect 154910 381134 155230 381218
rect 154910 380898 154952 381134
rect 155188 380898 155230 381134
rect 154910 380866 155230 380898
rect 160840 381454 161160 381486
rect 160840 381218 160882 381454
rect 161118 381218 161160 381454
rect 160840 381134 161160 381218
rect 160840 380898 160882 381134
rect 161118 380898 161160 381134
rect 160840 380866 161160 380898
rect 166771 381454 167091 381486
rect 166771 381218 166813 381454
rect 167049 381218 167091 381454
rect 166771 381134 167091 381218
rect 166771 380898 166813 381134
rect 167049 380898 167091 381134
rect 166771 380866 167091 380898
rect 181910 381454 182230 381486
rect 181910 381218 181952 381454
rect 182188 381218 182230 381454
rect 181910 381134 182230 381218
rect 181910 380898 181952 381134
rect 182188 380898 182230 381134
rect 181910 380866 182230 380898
rect 187840 381454 188160 381486
rect 187840 381218 187882 381454
rect 188118 381218 188160 381454
rect 187840 381134 188160 381218
rect 187840 380898 187882 381134
rect 188118 380898 188160 381134
rect 187840 380866 188160 380898
rect 193771 381454 194091 381486
rect 193771 381218 193813 381454
rect 194049 381218 194091 381454
rect 193771 381134 194091 381218
rect 193771 380898 193813 381134
rect 194049 380898 194091 381134
rect 193771 380866 194091 380898
rect 208910 381454 209230 381486
rect 208910 381218 208952 381454
rect 209188 381218 209230 381454
rect 208910 381134 209230 381218
rect 208910 380898 208952 381134
rect 209188 380898 209230 381134
rect 208910 380866 209230 380898
rect 214840 381454 215160 381486
rect 214840 381218 214882 381454
rect 215118 381218 215160 381454
rect 214840 381134 215160 381218
rect 214840 380898 214882 381134
rect 215118 380898 215160 381134
rect 214840 380866 215160 380898
rect 220771 381454 221091 381486
rect 220771 381218 220813 381454
rect 221049 381218 221091 381454
rect 220771 381134 221091 381218
rect 220771 380898 220813 381134
rect 221049 380898 221091 381134
rect 220771 380866 221091 380898
rect 235910 381454 236230 381486
rect 235910 381218 235952 381454
rect 236188 381218 236230 381454
rect 235910 381134 236230 381218
rect 235910 380898 235952 381134
rect 236188 380898 236230 381134
rect 235910 380866 236230 380898
rect 241840 381454 242160 381486
rect 241840 381218 241882 381454
rect 242118 381218 242160 381454
rect 241840 381134 242160 381218
rect 241840 380898 241882 381134
rect 242118 380898 242160 381134
rect 241840 380866 242160 380898
rect 247771 381454 248091 381486
rect 247771 381218 247813 381454
rect 248049 381218 248091 381454
rect 247771 381134 248091 381218
rect 247771 380898 247813 381134
rect 248049 380898 248091 381134
rect 247771 380866 248091 380898
rect 262910 381454 263230 381486
rect 262910 381218 262952 381454
rect 263188 381218 263230 381454
rect 262910 381134 263230 381218
rect 262910 380898 262952 381134
rect 263188 380898 263230 381134
rect 262910 380866 263230 380898
rect 268840 381454 269160 381486
rect 268840 381218 268882 381454
rect 269118 381218 269160 381454
rect 268840 381134 269160 381218
rect 268840 380898 268882 381134
rect 269118 380898 269160 381134
rect 268840 380866 269160 380898
rect 274771 381454 275091 381486
rect 274771 381218 274813 381454
rect 275049 381218 275091 381454
rect 274771 381134 275091 381218
rect 274771 380898 274813 381134
rect 275049 380898 275091 381134
rect 274771 380866 275091 380898
rect 289910 381454 290230 381486
rect 289910 381218 289952 381454
rect 290188 381218 290230 381454
rect 289910 381134 290230 381218
rect 289910 380898 289952 381134
rect 290188 380898 290230 381134
rect 289910 380866 290230 380898
rect 295840 381454 296160 381486
rect 295840 381218 295882 381454
rect 296118 381218 296160 381454
rect 295840 381134 296160 381218
rect 295840 380898 295882 381134
rect 296118 380898 296160 381134
rect 295840 380866 296160 380898
rect 301771 381454 302091 381486
rect 301771 381218 301813 381454
rect 302049 381218 302091 381454
rect 301771 381134 302091 381218
rect 301771 380898 301813 381134
rect 302049 380898 302091 381134
rect 301771 380866 302091 380898
rect 316910 381454 317230 381486
rect 316910 381218 316952 381454
rect 317188 381218 317230 381454
rect 316910 381134 317230 381218
rect 316910 380898 316952 381134
rect 317188 380898 317230 381134
rect 316910 380866 317230 380898
rect 322840 381454 323160 381486
rect 322840 381218 322882 381454
rect 323118 381218 323160 381454
rect 322840 381134 323160 381218
rect 322840 380898 322882 381134
rect 323118 380898 323160 381134
rect 322840 380866 323160 380898
rect 328771 381454 329091 381486
rect 328771 381218 328813 381454
rect 329049 381218 329091 381454
rect 328771 381134 329091 381218
rect 328771 380898 328813 381134
rect 329049 380898 329091 381134
rect 328771 380866 329091 380898
rect 343910 381454 344230 381486
rect 343910 381218 343952 381454
rect 344188 381218 344230 381454
rect 343910 381134 344230 381218
rect 343910 380898 343952 381134
rect 344188 380898 344230 381134
rect 343910 380866 344230 380898
rect 349840 381454 350160 381486
rect 349840 381218 349882 381454
rect 350118 381218 350160 381454
rect 349840 381134 350160 381218
rect 349840 380898 349882 381134
rect 350118 380898 350160 381134
rect 349840 380866 350160 380898
rect 355771 381454 356091 381486
rect 355771 381218 355813 381454
rect 356049 381218 356091 381454
rect 355771 381134 356091 381218
rect 355771 380898 355813 381134
rect 356049 380898 356091 381134
rect 355771 380866 356091 380898
rect 370910 381454 371230 381486
rect 370910 381218 370952 381454
rect 371188 381218 371230 381454
rect 370910 381134 371230 381218
rect 370910 380898 370952 381134
rect 371188 380898 371230 381134
rect 370910 380866 371230 380898
rect 376840 381454 377160 381486
rect 376840 381218 376882 381454
rect 377118 381218 377160 381454
rect 376840 381134 377160 381218
rect 376840 380898 376882 381134
rect 377118 380898 377160 381134
rect 376840 380866 377160 380898
rect 382771 381454 383091 381486
rect 382771 381218 382813 381454
rect 383049 381218 383091 381454
rect 382771 381134 383091 381218
rect 382771 380898 382813 381134
rect 383049 380898 383091 381134
rect 382771 380866 383091 380898
rect 397910 381454 398230 381486
rect 397910 381218 397952 381454
rect 398188 381218 398230 381454
rect 397910 381134 398230 381218
rect 397910 380898 397952 381134
rect 398188 380898 398230 381134
rect 397910 380866 398230 380898
rect 403840 381454 404160 381486
rect 403840 381218 403882 381454
rect 404118 381218 404160 381454
rect 403840 381134 404160 381218
rect 403840 380898 403882 381134
rect 404118 380898 404160 381134
rect 403840 380866 404160 380898
rect 409771 381454 410091 381486
rect 409771 381218 409813 381454
rect 410049 381218 410091 381454
rect 409771 381134 410091 381218
rect 409771 380898 409813 381134
rect 410049 380898 410091 381134
rect 409771 380866 410091 380898
rect 424910 381454 425230 381486
rect 424910 381218 424952 381454
rect 425188 381218 425230 381454
rect 424910 381134 425230 381218
rect 424910 380898 424952 381134
rect 425188 380898 425230 381134
rect 424910 380866 425230 380898
rect 430840 381454 431160 381486
rect 430840 381218 430882 381454
rect 431118 381218 431160 381454
rect 430840 381134 431160 381218
rect 430840 380898 430882 381134
rect 431118 380898 431160 381134
rect 430840 380866 431160 380898
rect 436771 381454 437091 381486
rect 436771 381218 436813 381454
rect 437049 381218 437091 381454
rect 436771 381134 437091 381218
rect 436771 380898 436813 381134
rect 437049 380898 437091 381134
rect 436771 380866 437091 380898
rect 451910 381454 452230 381486
rect 451910 381218 451952 381454
rect 452188 381218 452230 381454
rect 451910 381134 452230 381218
rect 451910 380898 451952 381134
rect 452188 380898 452230 381134
rect 451910 380866 452230 380898
rect 457840 381454 458160 381486
rect 457840 381218 457882 381454
rect 458118 381218 458160 381454
rect 457840 381134 458160 381218
rect 457840 380898 457882 381134
rect 458118 380898 458160 381134
rect 457840 380866 458160 380898
rect 463771 381454 464091 381486
rect 463771 381218 463813 381454
rect 464049 381218 464091 381454
rect 463771 381134 464091 381218
rect 463771 380898 463813 381134
rect 464049 380898 464091 381134
rect 463771 380866 464091 380898
rect 478910 381454 479230 381486
rect 478910 381218 478952 381454
rect 479188 381218 479230 381454
rect 478910 381134 479230 381218
rect 478910 380898 478952 381134
rect 479188 380898 479230 381134
rect 478910 380866 479230 380898
rect 484840 381454 485160 381486
rect 484840 381218 484882 381454
rect 485118 381218 485160 381454
rect 484840 381134 485160 381218
rect 484840 380898 484882 381134
rect 485118 380898 485160 381134
rect 484840 380866 485160 380898
rect 490771 381454 491091 381486
rect 490771 381218 490813 381454
rect 491049 381218 491091 381454
rect 490771 381134 491091 381218
rect 490771 380898 490813 381134
rect 491049 380898 491091 381134
rect 490771 380866 491091 380898
rect 505910 381454 506230 381486
rect 505910 381218 505952 381454
rect 506188 381218 506230 381454
rect 505910 381134 506230 381218
rect 505910 380898 505952 381134
rect 506188 380898 506230 381134
rect 505910 380866 506230 380898
rect 511840 381454 512160 381486
rect 511840 381218 511882 381454
rect 512118 381218 512160 381454
rect 511840 381134 512160 381218
rect 511840 380898 511882 381134
rect 512118 380898 512160 381134
rect 511840 380866 512160 380898
rect 517771 381454 518091 381486
rect 517771 381218 517813 381454
rect 518049 381218 518091 381454
rect 517771 381134 518091 381218
rect 517771 380898 517813 381134
rect 518049 380898 518091 381134
rect 517771 380866 518091 380898
rect 532910 381454 533230 381486
rect 532910 381218 532952 381454
rect 533188 381218 533230 381454
rect 532910 381134 533230 381218
rect 532910 380898 532952 381134
rect 533188 380898 533230 381134
rect 532910 380866 533230 380898
rect 538840 381454 539160 381486
rect 538840 381218 538882 381454
rect 539118 381218 539160 381454
rect 538840 381134 539160 381218
rect 538840 380898 538882 381134
rect 539118 380898 539160 381134
rect 538840 380866 539160 380898
rect 544771 381454 545091 381486
rect 544771 381218 544813 381454
rect 545049 381218 545091 381454
rect 544771 381134 545091 381218
rect 544771 380898 544813 381134
rect 545049 380898 545091 381134
rect 544771 380866 545091 380898
rect 559794 381454 560414 398898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 354454 11414 371898
rect 22874 372454 23194 372486
rect 22874 372218 22916 372454
rect 23152 372218 23194 372454
rect 22874 372134 23194 372218
rect 22874 371898 22916 372134
rect 23152 371898 23194 372134
rect 22874 371866 23194 371898
rect 28805 372454 29125 372486
rect 28805 372218 28847 372454
rect 29083 372218 29125 372454
rect 28805 372134 29125 372218
rect 28805 371898 28847 372134
rect 29083 371898 29125 372134
rect 28805 371866 29125 371898
rect 49874 372454 50194 372486
rect 49874 372218 49916 372454
rect 50152 372218 50194 372454
rect 49874 372134 50194 372218
rect 49874 371898 49916 372134
rect 50152 371898 50194 372134
rect 49874 371866 50194 371898
rect 55805 372454 56125 372486
rect 55805 372218 55847 372454
rect 56083 372218 56125 372454
rect 55805 372134 56125 372218
rect 55805 371898 55847 372134
rect 56083 371898 56125 372134
rect 55805 371866 56125 371898
rect 76874 372454 77194 372486
rect 76874 372218 76916 372454
rect 77152 372218 77194 372454
rect 76874 372134 77194 372218
rect 76874 371898 76916 372134
rect 77152 371898 77194 372134
rect 76874 371866 77194 371898
rect 82805 372454 83125 372486
rect 82805 372218 82847 372454
rect 83083 372218 83125 372454
rect 82805 372134 83125 372218
rect 82805 371898 82847 372134
rect 83083 371898 83125 372134
rect 82805 371866 83125 371898
rect 103874 372454 104194 372486
rect 103874 372218 103916 372454
rect 104152 372218 104194 372454
rect 103874 372134 104194 372218
rect 103874 371898 103916 372134
rect 104152 371898 104194 372134
rect 103874 371866 104194 371898
rect 109805 372454 110125 372486
rect 109805 372218 109847 372454
rect 110083 372218 110125 372454
rect 109805 372134 110125 372218
rect 109805 371898 109847 372134
rect 110083 371898 110125 372134
rect 109805 371866 110125 371898
rect 130874 372454 131194 372486
rect 130874 372218 130916 372454
rect 131152 372218 131194 372454
rect 130874 372134 131194 372218
rect 130874 371898 130916 372134
rect 131152 371898 131194 372134
rect 130874 371866 131194 371898
rect 136805 372454 137125 372486
rect 136805 372218 136847 372454
rect 137083 372218 137125 372454
rect 136805 372134 137125 372218
rect 136805 371898 136847 372134
rect 137083 371898 137125 372134
rect 136805 371866 137125 371898
rect 157874 372454 158194 372486
rect 157874 372218 157916 372454
rect 158152 372218 158194 372454
rect 157874 372134 158194 372218
rect 157874 371898 157916 372134
rect 158152 371898 158194 372134
rect 157874 371866 158194 371898
rect 163805 372454 164125 372486
rect 163805 372218 163847 372454
rect 164083 372218 164125 372454
rect 163805 372134 164125 372218
rect 163805 371898 163847 372134
rect 164083 371898 164125 372134
rect 163805 371866 164125 371898
rect 184874 372454 185194 372486
rect 184874 372218 184916 372454
rect 185152 372218 185194 372454
rect 184874 372134 185194 372218
rect 184874 371898 184916 372134
rect 185152 371898 185194 372134
rect 184874 371866 185194 371898
rect 190805 372454 191125 372486
rect 190805 372218 190847 372454
rect 191083 372218 191125 372454
rect 190805 372134 191125 372218
rect 190805 371898 190847 372134
rect 191083 371898 191125 372134
rect 190805 371866 191125 371898
rect 211874 372454 212194 372486
rect 211874 372218 211916 372454
rect 212152 372218 212194 372454
rect 211874 372134 212194 372218
rect 211874 371898 211916 372134
rect 212152 371898 212194 372134
rect 211874 371866 212194 371898
rect 217805 372454 218125 372486
rect 217805 372218 217847 372454
rect 218083 372218 218125 372454
rect 217805 372134 218125 372218
rect 217805 371898 217847 372134
rect 218083 371898 218125 372134
rect 217805 371866 218125 371898
rect 238874 372454 239194 372486
rect 238874 372218 238916 372454
rect 239152 372218 239194 372454
rect 238874 372134 239194 372218
rect 238874 371898 238916 372134
rect 239152 371898 239194 372134
rect 238874 371866 239194 371898
rect 244805 372454 245125 372486
rect 244805 372218 244847 372454
rect 245083 372218 245125 372454
rect 244805 372134 245125 372218
rect 244805 371898 244847 372134
rect 245083 371898 245125 372134
rect 244805 371866 245125 371898
rect 265874 372454 266194 372486
rect 265874 372218 265916 372454
rect 266152 372218 266194 372454
rect 265874 372134 266194 372218
rect 265874 371898 265916 372134
rect 266152 371898 266194 372134
rect 265874 371866 266194 371898
rect 271805 372454 272125 372486
rect 271805 372218 271847 372454
rect 272083 372218 272125 372454
rect 271805 372134 272125 372218
rect 271805 371898 271847 372134
rect 272083 371898 272125 372134
rect 271805 371866 272125 371898
rect 292874 372454 293194 372486
rect 292874 372218 292916 372454
rect 293152 372218 293194 372454
rect 292874 372134 293194 372218
rect 292874 371898 292916 372134
rect 293152 371898 293194 372134
rect 292874 371866 293194 371898
rect 298805 372454 299125 372486
rect 298805 372218 298847 372454
rect 299083 372218 299125 372454
rect 298805 372134 299125 372218
rect 298805 371898 298847 372134
rect 299083 371898 299125 372134
rect 298805 371866 299125 371898
rect 319874 372454 320194 372486
rect 319874 372218 319916 372454
rect 320152 372218 320194 372454
rect 319874 372134 320194 372218
rect 319874 371898 319916 372134
rect 320152 371898 320194 372134
rect 319874 371866 320194 371898
rect 325805 372454 326125 372486
rect 325805 372218 325847 372454
rect 326083 372218 326125 372454
rect 325805 372134 326125 372218
rect 325805 371898 325847 372134
rect 326083 371898 326125 372134
rect 325805 371866 326125 371898
rect 346874 372454 347194 372486
rect 346874 372218 346916 372454
rect 347152 372218 347194 372454
rect 346874 372134 347194 372218
rect 346874 371898 346916 372134
rect 347152 371898 347194 372134
rect 346874 371866 347194 371898
rect 352805 372454 353125 372486
rect 352805 372218 352847 372454
rect 353083 372218 353125 372454
rect 352805 372134 353125 372218
rect 352805 371898 352847 372134
rect 353083 371898 353125 372134
rect 352805 371866 353125 371898
rect 373874 372454 374194 372486
rect 373874 372218 373916 372454
rect 374152 372218 374194 372454
rect 373874 372134 374194 372218
rect 373874 371898 373916 372134
rect 374152 371898 374194 372134
rect 373874 371866 374194 371898
rect 379805 372454 380125 372486
rect 379805 372218 379847 372454
rect 380083 372218 380125 372454
rect 379805 372134 380125 372218
rect 379805 371898 379847 372134
rect 380083 371898 380125 372134
rect 379805 371866 380125 371898
rect 400874 372454 401194 372486
rect 400874 372218 400916 372454
rect 401152 372218 401194 372454
rect 400874 372134 401194 372218
rect 400874 371898 400916 372134
rect 401152 371898 401194 372134
rect 400874 371866 401194 371898
rect 406805 372454 407125 372486
rect 406805 372218 406847 372454
rect 407083 372218 407125 372454
rect 406805 372134 407125 372218
rect 406805 371898 406847 372134
rect 407083 371898 407125 372134
rect 406805 371866 407125 371898
rect 427874 372454 428194 372486
rect 427874 372218 427916 372454
rect 428152 372218 428194 372454
rect 427874 372134 428194 372218
rect 427874 371898 427916 372134
rect 428152 371898 428194 372134
rect 427874 371866 428194 371898
rect 433805 372454 434125 372486
rect 433805 372218 433847 372454
rect 434083 372218 434125 372454
rect 433805 372134 434125 372218
rect 433805 371898 433847 372134
rect 434083 371898 434125 372134
rect 433805 371866 434125 371898
rect 454874 372454 455194 372486
rect 454874 372218 454916 372454
rect 455152 372218 455194 372454
rect 454874 372134 455194 372218
rect 454874 371898 454916 372134
rect 455152 371898 455194 372134
rect 454874 371866 455194 371898
rect 460805 372454 461125 372486
rect 460805 372218 460847 372454
rect 461083 372218 461125 372454
rect 460805 372134 461125 372218
rect 460805 371898 460847 372134
rect 461083 371898 461125 372134
rect 460805 371866 461125 371898
rect 481874 372454 482194 372486
rect 481874 372218 481916 372454
rect 482152 372218 482194 372454
rect 481874 372134 482194 372218
rect 481874 371898 481916 372134
rect 482152 371898 482194 372134
rect 481874 371866 482194 371898
rect 487805 372454 488125 372486
rect 487805 372218 487847 372454
rect 488083 372218 488125 372454
rect 487805 372134 488125 372218
rect 487805 371898 487847 372134
rect 488083 371898 488125 372134
rect 487805 371866 488125 371898
rect 508874 372454 509194 372486
rect 508874 372218 508916 372454
rect 509152 372218 509194 372454
rect 508874 372134 509194 372218
rect 508874 371898 508916 372134
rect 509152 371898 509194 372134
rect 508874 371866 509194 371898
rect 514805 372454 515125 372486
rect 514805 372218 514847 372454
rect 515083 372218 515125 372454
rect 514805 372134 515125 372218
rect 514805 371898 514847 372134
rect 515083 371898 515125 372134
rect 514805 371866 515125 371898
rect 535874 372454 536194 372486
rect 535874 372218 535916 372454
rect 536152 372218 536194 372454
rect 535874 372134 536194 372218
rect 535874 371898 535916 372134
rect 536152 371898 536194 372134
rect 535874 371866 536194 371898
rect 541805 372454 542125 372486
rect 541805 372218 541847 372454
rect 542083 372218 542125 372454
rect 541805 372134 542125 372218
rect 541805 371898 541847 372134
rect 542083 371898 542125 372134
rect 541805 371866 542125 371898
rect 19794 363454 20414 365000
rect 19794 363218 19826 363454
rect 20062 363218 20146 363454
rect 20382 363218 20414 363454
rect 19794 363134 20414 363218
rect 19794 362898 19826 363134
rect 20062 362898 20146 363134
rect 20382 362898 20414 363134
rect 19794 362000 20414 362898
rect 28794 364394 29414 365000
rect 28794 364158 28826 364394
rect 29062 364158 29146 364394
rect 29382 364158 29414 364394
rect 28794 364074 29414 364158
rect 28794 363838 28826 364074
rect 29062 363838 29146 364074
rect 29382 363838 29414 364074
rect 28794 362000 29414 363838
rect 37794 363454 38414 365000
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 362000 38414 362898
rect 46794 364394 47414 365000
rect 46794 364158 46826 364394
rect 47062 364158 47146 364394
rect 47382 364158 47414 364394
rect 46794 364074 47414 364158
rect 46794 363838 46826 364074
rect 47062 363838 47146 364074
rect 47382 363838 47414 364074
rect 46794 362000 47414 363838
rect 55794 363454 56414 365000
rect 55794 363218 55826 363454
rect 56062 363218 56146 363454
rect 56382 363218 56414 363454
rect 55794 363134 56414 363218
rect 55794 362898 55826 363134
rect 56062 362898 56146 363134
rect 56382 362898 56414 363134
rect 55794 362000 56414 362898
rect 64794 364394 65414 365000
rect 64794 364158 64826 364394
rect 65062 364158 65146 364394
rect 65382 364158 65414 364394
rect 64794 364074 65414 364158
rect 64794 363838 64826 364074
rect 65062 363838 65146 364074
rect 65382 363838 65414 364074
rect 64794 362000 65414 363838
rect 73794 363454 74414 365000
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 362000 74414 362898
rect 82794 364394 83414 365000
rect 82794 364158 82826 364394
rect 83062 364158 83146 364394
rect 83382 364158 83414 364394
rect 82794 364074 83414 364158
rect 82794 363838 82826 364074
rect 83062 363838 83146 364074
rect 83382 363838 83414 364074
rect 82794 362000 83414 363838
rect 91794 363454 92414 365000
rect 91794 363218 91826 363454
rect 92062 363218 92146 363454
rect 92382 363218 92414 363454
rect 91794 363134 92414 363218
rect 91794 362898 91826 363134
rect 92062 362898 92146 363134
rect 92382 362898 92414 363134
rect 91794 362000 92414 362898
rect 100794 364394 101414 365000
rect 100794 364158 100826 364394
rect 101062 364158 101146 364394
rect 101382 364158 101414 364394
rect 100794 364074 101414 364158
rect 100794 363838 100826 364074
rect 101062 363838 101146 364074
rect 101382 363838 101414 364074
rect 100794 362000 101414 363838
rect 109794 363454 110414 365000
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 362000 110414 362898
rect 118794 364394 119414 365000
rect 118794 364158 118826 364394
rect 119062 364158 119146 364394
rect 119382 364158 119414 364394
rect 118794 364074 119414 364158
rect 118794 363838 118826 364074
rect 119062 363838 119146 364074
rect 119382 363838 119414 364074
rect 118794 362000 119414 363838
rect 127794 363454 128414 365000
rect 127794 363218 127826 363454
rect 128062 363218 128146 363454
rect 128382 363218 128414 363454
rect 127794 363134 128414 363218
rect 127794 362898 127826 363134
rect 128062 362898 128146 363134
rect 128382 362898 128414 363134
rect 127794 362000 128414 362898
rect 136794 364394 137414 365000
rect 136794 364158 136826 364394
rect 137062 364158 137146 364394
rect 137382 364158 137414 364394
rect 136794 364074 137414 364158
rect 136794 363838 136826 364074
rect 137062 363838 137146 364074
rect 137382 363838 137414 364074
rect 136794 362000 137414 363838
rect 145794 363454 146414 365000
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 362000 146414 362898
rect 154794 364394 155414 365000
rect 154794 364158 154826 364394
rect 155062 364158 155146 364394
rect 155382 364158 155414 364394
rect 154794 364074 155414 364158
rect 154794 363838 154826 364074
rect 155062 363838 155146 364074
rect 155382 363838 155414 364074
rect 154794 362000 155414 363838
rect 163794 363454 164414 365000
rect 163794 363218 163826 363454
rect 164062 363218 164146 363454
rect 164382 363218 164414 363454
rect 163794 363134 164414 363218
rect 163794 362898 163826 363134
rect 164062 362898 164146 363134
rect 164382 362898 164414 363134
rect 163794 362000 164414 362898
rect 172794 364394 173414 365000
rect 172794 364158 172826 364394
rect 173062 364158 173146 364394
rect 173382 364158 173414 364394
rect 172794 364074 173414 364158
rect 172794 363838 172826 364074
rect 173062 363838 173146 364074
rect 173382 363838 173414 364074
rect 172794 362000 173414 363838
rect 181794 363454 182414 365000
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 362000 182414 362898
rect 190794 364394 191414 365000
rect 190794 364158 190826 364394
rect 191062 364158 191146 364394
rect 191382 364158 191414 364394
rect 190794 364074 191414 364158
rect 190794 363838 190826 364074
rect 191062 363838 191146 364074
rect 191382 363838 191414 364074
rect 190794 362000 191414 363838
rect 199794 363454 200414 365000
rect 199794 363218 199826 363454
rect 200062 363218 200146 363454
rect 200382 363218 200414 363454
rect 199794 363134 200414 363218
rect 199794 362898 199826 363134
rect 200062 362898 200146 363134
rect 200382 362898 200414 363134
rect 199794 362000 200414 362898
rect 208794 364394 209414 365000
rect 208794 364158 208826 364394
rect 209062 364158 209146 364394
rect 209382 364158 209414 364394
rect 208794 364074 209414 364158
rect 208794 363838 208826 364074
rect 209062 363838 209146 364074
rect 209382 363838 209414 364074
rect 208794 362000 209414 363838
rect 217794 363454 218414 365000
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 362000 218414 362898
rect 226794 364394 227414 365000
rect 226794 364158 226826 364394
rect 227062 364158 227146 364394
rect 227382 364158 227414 364394
rect 226794 364074 227414 364158
rect 226794 363838 226826 364074
rect 227062 363838 227146 364074
rect 227382 363838 227414 364074
rect 226794 362000 227414 363838
rect 235794 363454 236414 365000
rect 235794 363218 235826 363454
rect 236062 363218 236146 363454
rect 236382 363218 236414 363454
rect 235794 363134 236414 363218
rect 235794 362898 235826 363134
rect 236062 362898 236146 363134
rect 236382 362898 236414 363134
rect 235794 362000 236414 362898
rect 244794 364394 245414 365000
rect 244794 364158 244826 364394
rect 245062 364158 245146 364394
rect 245382 364158 245414 364394
rect 244794 364074 245414 364158
rect 244794 363838 244826 364074
rect 245062 363838 245146 364074
rect 245382 363838 245414 364074
rect 244794 362000 245414 363838
rect 253794 363454 254414 365000
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 362000 254414 362898
rect 262794 364394 263414 365000
rect 262794 364158 262826 364394
rect 263062 364158 263146 364394
rect 263382 364158 263414 364394
rect 262794 364074 263414 364158
rect 262794 363838 262826 364074
rect 263062 363838 263146 364074
rect 263382 363838 263414 364074
rect 262794 362000 263414 363838
rect 271794 363454 272414 365000
rect 271794 363218 271826 363454
rect 272062 363218 272146 363454
rect 272382 363218 272414 363454
rect 271794 363134 272414 363218
rect 271794 362898 271826 363134
rect 272062 362898 272146 363134
rect 272382 362898 272414 363134
rect 271794 362000 272414 362898
rect 280794 364394 281414 365000
rect 280794 364158 280826 364394
rect 281062 364158 281146 364394
rect 281382 364158 281414 364394
rect 280794 364074 281414 364158
rect 280794 363838 280826 364074
rect 281062 363838 281146 364074
rect 281382 363838 281414 364074
rect 280794 362000 281414 363838
rect 289794 363454 290414 365000
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 362000 290414 362898
rect 298794 364394 299414 365000
rect 298794 364158 298826 364394
rect 299062 364158 299146 364394
rect 299382 364158 299414 364394
rect 298794 364074 299414 364158
rect 298794 363838 298826 364074
rect 299062 363838 299146 364074
rect 299382 363838 299414 364074
rect 298794 362000 299414 363838
rect 307794 363454 308414 365000
rect 307794 363218 307826 363454
rect 308062 363218 308146 363454
rect 308382 363218 308414 363454
rect 307794 363134 308414 363218
rect 307794 362898 307826 363134
rect 308062 362898 308146 363134
rect 308382 362898 308414 363134
rect 307794 362000 308414 362898
rect 316794 364394 317414 365000
rect 316794 364158 316826 364394
rect 317062 364158 317146 364394
rect 317382 364158 317414 364394
rect 316794 364074 317414 364158
rect 316794 363838 316826 364074
rect 317062 363838 317146 364074
rect 317382 363838 317414 364074
rect 316794 362000 317414 363838
rect 325794 363454 326414 365000
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 362000 326414 362898
rect 334794 364394 335414 365000
rect 334794 364158 334826 364394
rect 335062 364158 335146 364394
rect 335382 364158 335414 364394
rect 334794 364074 335414 364158
rect 334794 363838 334826 364074
rect 335062 363838 335146 364074
rect 335382 363838 335414 364074
rect 334794 362000 335414 363838
rect 343794 363454 344414 365000
rect 343794 363218 343826 363454
rect 344062 363218 344146 363454
rect 344382 363218 344414 363454
rect 343794 363134 344414 363218
rect 343794 362898 343826 363134
rect 344062 362898 344146 363134
rect 344382 362898 344414 363134
rect 343794 362000 344414 362898
rect 352794 364394 353414 365000
rect 352794 364158 352826 364394
rect 353062 364158 353146 364394
rect 353382 364158 353414 364394
rect 352794 364074 353414 364158
rect 352794 363838 352826 364074
rect 353062 363838 353146 364074
rect 353382 363838 353414 364074
rect 352794 362000 353414 363838
rect 361794 363454 362414 365000
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 362000 362414 362898
rect 370794 364394 371414 365000
rect 370794 364158 370826 364394
rect 371062 364158 371146 364394
rect 371382 364158 371414 364394
rect 370794 364074 371414 364158
rect 370794 363838 370826 364074
rect 371062 363838 371146 364074
rect 371382 363838 371414 364074
rect 370794 362000 371414 363838
rect 379794 363454 380414 365000
rect 379794 363218 379826 363454
rect 380062 363218 380146 363454
rect 380382 363218 380414 363454
rect 379794 363134 380414 363218
rect 379794 362898 379826 363134
rect 380062 362898 380146 363134
rect 380382 362898 380414 363134
rect 379794 362000 380414 362898
rect 388794 364394 389414 365000
rect 388794 364158 388826 364394
rect 389062 364158 389146 364394
rect 389382 364158 389414 364394
rect 388794 364074 389414 364158
rect 388794 363838 388826 364074
rect 389062 363838 389146 364074
rect 389382 363838 389414 364074
rect 388794 362000 389414 363838
rect 397794 363454 398414 365000
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 362000 398414 362898
rect 406794 364394 407414 365000
rect 406794 364158 406826 364394
rect 407062 364158 407146 364394
rect 407382 364158 407414 364394
rect 406794 364074 407414 364158
rect 406794 363838 406826 364074
rect 407062 363838 407146 364074
rect 407382 363838 407414 364074
rect 406794 362000 407414 363838
rect 415794 363454 416414 365000
rect 415794 363218 415826 363454
rect 416062 363218 416146 363454
rect 416382 363218 416414 363454
rect 415794 363134 416414 363218
rect 415794 362898 415826 363134
rect 416062 362898 416146 363134
rect 416382 362898 416414 363134
rect 415794 362000 416414 362898
rect 424794 364394 425414 365000
rect 424794 364158 424826 364394
rect 425062 364158 425146 364394
rect 425382 364158 425414 364394
rect 424794 364074 425414 364158
rect 424794 363838 424826 364074
rect 425062 363838 425146 364074
rect 425382 363838 425414 364074
rect 424794 362000 425414 363838
rect 433794 363454 434414 365000
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 362000 434414 362898
rect 442794 364394 443414 365000
rect 442794 364158 442826 364394
rect 443062 364158 443146 364394
rect 443382 364158 443414 364394
rect 442794 364074 443414 364158
rect 442794 363838 442826 364074
rect 443062 363838 443146 364074
rect 443382 363838 443414 364074
rect 442794 362000 443414 363838
rect 451794 363454 452414 365000
rect 451794 363218 451826 363454
rect 452062 363218 452146 363454
rect 452382 363218 452414 363454
rect 451794 363134 452414 363218
rect 451794 362898 451826 363134
rect 452062 362898 452146 363134
rect 452382 362898 452414 363134
rect 451794 362000 452414 362898
rect 460794 364394 461414 365000
rect 460794 364158 460826 364394
rect 461062 364158 461146 364394
rect 461382 364158 461414 364394
rect 460794 364074 461414 364158
rect 460794 363838 460826 364074
rect 461062 363838 461146 364074
rect 461382 363838 461414 364074
rect 460794 362000 461414 363838
rect 469794 363454 470414 365000
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 362000 470414 362898
rect 478794 364394 479414 365000
rect 478794 364158 478826 364394
rect 479062 364158 479146 364394
rect 479382 364158 479414 364394
rect 478794 364074 479414 364158
rect 478794 363838 478826 364074
rect 479062 363838 479146 364074
rect 479382 363838 479414 364074
rect 478794 362000 479414 363838
rect 487794 363454 488414 365000
rect 487794 363218 487826 363454
rect 488062 363218 488146 363454
rect 488382 363218 488414 363454
rect 487794 363134 488414 363218
rect 487794 362898 487826 363134
rect 488062 362898 488146 363134
rect 488382 362898 488414 363134
rect 487794 362000 488414 362898
rect 496794 364394 497414 365000
rect 496794 364158 496826 364394
rect 497062 364158 497146 364394
rect 497382 364158 497414 364394
rect 496794 364074 497414 364158
rect 496794 363838 496826 364074
rect 497062 363838 497146 364074
rect 497382 363838 497414 364074
rect 496794 362000 497414 363838
rect 505794 363454 506414 365000
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 362000 506414 362898
rect 514794 364394 515414 365000
rect 514794 364158 514826 364394
rect 515062 364158 515146 364394
rect 515382 364158 515414 364394
rect 514794 364074 515414 364158
rect 514794 363838 514826 364074
rect 515062 363838 515146 364074
rect 515382 363838 515414 364074
rect 514794 362000 515414 363838
rect 523794 363454 524414 365000
rect 523794 363218 523826 363454
rect 524062 363218 524146 363454
rect 524382 363218 524414 363454
rect 523794 363134 524414 363218
rect 523794 362898 523826 363134
rect 524062 362898 524146 363134
rect 524382 362898 524414 363134
rect 523794 362000 524414 362898
rect 532794 364394 533414 365000
rect 532794 364158 532826 364394
rect 533062 364158 533146 364394
rect 533382 364158 533414 364394
rect 532794 364074 533414 364158
rect 532794 363838 532826 364074
rect 533062 363838 533146 364074
rect 533382 363838 533414 364074
rect 532794 362000 533414 363838
rect 541794 363454 542414 365000
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 362000 542414 362898
rect 550794 364394 551414 365000
rect 550794 364158 550826 364394
rect 551062 364158 551146 364394
rect 551382 364158 551414 364394
rect 550794 364074 551414 364158
rect 550794 363838 550826 364074
rect 551062 363838 551146 364074
rect 551382 363838 551414 364074
rect 550794 362000 551414 363838
rect 559794 363454 560414 380898
rect 559794 363218 559826 363454
rect 560062 363218 560146 363454
rect 560382 363218 560414 363454
rect 559794 363134 560414 363218
rect 559794 362898 559826 363134
rect 560062 362898 560146 363134
rect 560382 362898 560414 363134
rect 10794 354218 10826 354454
rect 11062 354218 11146 354454
rect 11382 354218 11414 354454
rect 10794 354134 11414 354218
rect 10794 353898 10826 354134
rect 11062 353898 11146 354134
rect 11382 353898 11414 354134
rect 10794 336454 11414 353898
rect 22874 354454 23194 354486
rect 22874 354218 22916 354454
rect 23152 354218 23194 354454
rect 22874 354134 23194 354218
rect 22874 353898 22916 354134
rect 23152 353898 23194 354134
rect 22874 353866 23194 353898
rect 28805 354454 29125 354486
rect 28805 354218 28847 354454
rect 29083 354218 29125 354454
rect 28805 354134 29125 354218
rect 28805 353898 28847 354134
rect 29083 353898 29125 354134
rect 28805 353866 29125 353898
rect 49874 354454 50194 354486
rect 49874 354218 49916 354454
rect 50152 354218 50194 354454
rect 49874 354134 50194 354218
rect 49874 353898 49916 354134
rect 50152 353898 50194 354134
rect 49874 353866 50194 353898
rect 55805 354454 56125 354486
rect 55805 354218 55847 354454
rect 56083 354218 56125 354454
rect 55805 354134 56125 354218
rect 55805 353898 55847 354134
rect 56083 353898 56125 354134
rect 55805 353866 56125 353898
rect 76874 354454 77194 354486
rect 76874 354218 76916 354454
rect 77152 354218 77194 354454
rect 76874 354134 77194 354218
rect 76874 353898 76916 354134
rect 77152 353898 77194 354134
rect 76874 353866 77194 353898
rect 82805 354454 83125 354486
rect 82805 354218 82847 354454
rect 83083 354218 83125 354454
rect 82805 354134 83125 354218
rect 82805 353898 82847 354134
rect 83083 353898 83125 354134
rect 82805 353866 83125 353898
rect 103874 354454 104194 354486
rect 103874 354218 103916 354454
rect 104152 354218 104194 354454
rect 103874 354134 104194 354218
rect 103874 353898 103916 354134
rect 104152 353898 104194 354134
rect 103874 353866 104194 353898
rect 109805 354454 110125 354486
rect 109805 354218 109847 354454
rect 110083 354218 110125 354454
rect 109805 354134 110125 354218
rect 109805 353898 109847 354134
rect 110083 353898 110125 354134
rect 109805 353866 110125 353898
rect 130874 354454 131194 354486
rect 130874 354218 130916 354454
rect 131152 354218 131194 354454
rect 130874 354134 131194 354218
rect 130874 353898 130916 354134
rect 131152 353898 131194 354134
rect 130874 353866 131194 353898
rect 136805 354454 137125 354486
rect 136805 354218 136847 354454
rect 137083 354218 137125 354454
rect 136805 354134 137125 354218
rect 136805 353898 136847 354134
rect 137083 353898 137125 354134
rect 136805 353866 137125 353898
rect 157874 354454 158194 354486
rect 157874 354218 157916 354454
rect 158152 354218 158194 354454
rect 157874 354134 158194 354218
rect 157874 353898 157916 354134
rect 158152 353898 158194 354134
rect 157874 353866 158194 353898
rect 163805 354454 164125 354486
rect 163805 354218 163847 354454
rect 164083 354218 164125 354454
rect 163805 354134 164125 354218
rect 163805 353898 163847 354134
rect 164083 353898 164125 354134
rect 163805 353866 164125 353898
rect 184874 354454 185194 354486
rect 184874 354218 184916 354454
rect 185152 354218 185194 354454
rect 184874 354134 185194 354218
rect 184874 353898 184916 354134
rect 185152 353898 185194 354134
rect 184874 353866 185194 353898
rect 190805 354454 191125 354486
rect 190805 354218 190847 354454
rect 191083 354218 191125 354454
rect 190805 354134 191125 354218
rect 190805 353898 190847 354134
rect 191083 353898 191125 354134
rect 190805 353866 191125 353898
rect 211874 354454 212194 354486
rect 211874 354218 211916 354454
rect 212152 354218 212194 354454
rect 211874 354134 212194 354218
rect 211874 353898 211916 354134
rect 212152 353898 212194 354134
rect 211874 353866 212194 353898
rect 217805 354454 218125 354486
rect 217805 354218 217847 354454
rect 218083 354218 218125 354454
rect 217805 354134 218125 354218
rect 217805 353898 217847 354134
rect 218083 353898 218125 354134
rect 217805 353866 218125 353898
rect 238874 354454 239194 354486
rect 238874 354218 238916 354454
rect 239152 354218 239194 354454
rect 238874 354134 239194 354218
rect 238874 353898 238916 354134
rect 239152 353898 239194 354134
rect 238874 353866 239194 353898
rect 244805 354454 245125 354486
rect 244805 354218 244847 354454
rect 245083 354218 245125 354454
rect 244805 354134 245125 354218
rect 244805 353898 244847 354134
rect 245083 353898 245125 354134
rect 244805 353866 245125 353898
rect 265874 354454 266194 354486
rect 265874 354218 265916 354454
rect 266152 354218 266194 354454
rect 265874 354134 266194 354218
rect 265874 353898 265916 354134
rect 266152 353898 266194 354134
rect 265874 353866 266194 353898
rect 271805 354454 272125 354486
rect 271805 354218 271847 354454
rect 272083 354218 272125 354454
rect 271805 354134 272125 354218
rect 271805 353898 271847 354134
rect 272083 353898 272125 354134
rect 271805 353866 272125 353898
rect 292874 354454 293194 354486
rect 292874 354218 292916 354454
rect 293152 354218 293194 354454
rect 292874 354134 293194 354218
rect 292874 353898 292916 354134
rect 293152 353898 293194 354134
rect 292874 353866 293194 353898
rect 298805 354454 299125 354486
rect 298805 354218 298847 354454
rect 299083 354218 299125 354454
rect 298805 354134 299125 354218
rect 298805 353898 298847 354134
rect 299083 353898 299125 354134
rect 298805 353866 299125 353898
rect 319874 354454 320194 354486
rect 319874 354218 319916 354454
rect 320152 354218 320194 354454
rect 319874 354134 320194 354218
rect 319874 353898 319916 354134
rect 320152 353898 320194 354134
rect 319874 353866 320194 353898
rect 325805 354454 326125 354486
rect 325805 354218 325847 354454
rect 326083 354218 326125 354454
rect 325805 354134 326125 354218
rect 325805 353898 325847 354134
rect 326083 353898 326125 354134
rect 325805 353866 326125 353898
rect 346874 354454 347194 354486
rect 346874 354218 346916 354454
rect 347152 354218 347194 354454
rect 346874 354134 347194 354218
rect 346874 353898 346916 354134
rect 347152 353898 347194 354134
rect 346874 353866 347194 353898
rect 352805 354454 353125 354486
rect 352805 354218 352847 354454
rect 353083 354218 353125 354454
rect 352805 354134 353125 354218
rect 352805 353898 352847 354134
rect 353083 353898 353125 354134
rect 352805 353866 353125 353898
rect 373874 354454 374194 354486
rect 373874 354218 373916 354454
rect 374152 354218 374194 354454
rect 373874 354134 374194 354218
rect 373874 353898 373916 354134
rect 374152 353898 374194 354134
rect 373874 353866 374194 353898
rect 379805 354454 380125 354486
rect 379805 354218 379847 354454
rect 380083 354218 380125 354454
rect 379805 354134 380125 354218
rect 379805 353898 379847 354134
rect 380083 353898 380125 354134
rect 379805 353866 380125 353898
rect 400874 354454 401194 354486
rect 400874 354218 400916 354454
rect 401152 354218 401194 354454
rect 400874 354134 401194 354218
rect 400874 353898 400916 354134
rect 401152 353898 401194 354134
rect 400874 353866 401194 353898
rect 406805 354454 407125 354486
rect 406805 354218 406847 354454
rect 407083 354218 407125 354454
rect 406805 354134 407125 354218
rect 406805 353898 406847 354134
rect 407083 353898 407125 354134
rect 406805 353866 407125 353898
rect 427874 354454 428194 354486
rect 427874 354218 427916 354454
rect 428152 354218 428194 354454
rect 427874 354134 428194 354218
rect 427874 353898 427916 354134
rect 428152 353898 428194 354134
rect 427874 353866 428194 353898
rect 433805 354454 434125 354486
rect 433805 354218 433847 354454
rect 434083 354218 434125 354454
rect 433805 354134 434125 354218
rect 433805 353898 433847 354134
rect 434083 353898 434125 354134
rect 433805 353866 434125 353898
rect 454874 354454 455194 354486
rect 454874 354218 454916 354454
rect 455152 354218 455194 354454
rect 454874 354134 455194 354218
rect 454874 353898 454916 354134
rect 455152 353898 455194 354134
rect 454874 353866 455194 353898
rect 460805 354454 461125 354486
rect 460805 354218 460847 354454
rect 461083 354218 461125 354454
rect 460805 354134 461125 354218
rect 460805 353898 460847 354134
rect 461083 353898 461125 354134
rect 460805 353866 461125 353898
rect 481874 354454 482194 354486
rect 481874 354218 481916 354454
rect 482152 354218 482194 354454
rect 481874 354134 482194 354218
rect 481874 353898 481916 354134
rect 482152 353898 482194 354134
rect 481874 353866 482194 353898
rect 487805 354454 488125 354486
rect 487805 354218 487847 354454
rect 488083 354218 488125 354454
rect 487805 354134 488125 354218
rect 487805 353898 487847 354134
rect 488083 353898 488125 354134
rect 487805 353866 488125 353898
rect 508874 354454 509194 354486
rect 508874 354218 508916 354454
rect 509152 354218 509194 354454
rect 508874 354134 509194 354218
rect 508874 353898 508916 354134
rect 509152 353898 509194 354134
rect 508874 353866 509194 353898
rect 514805 354454 515125 354486
rect 514805 354218 514847 354454
rect 515083 354218 515125 354454
rect 514805 354134 515125 354218
rect 514805 353898 514847 354134
rect 515083 353898 515125 354134
rect 514805 353866 515125 353898
rect 535874 354454 536194 354486
rect 535874 354218 535916 354454
rect 536152 354218 536194 354454
rect 535874 354134 536194 354218
rect 535874 353898 535916 354134
rect 536152 353898 536194 354134
rect 535874 353866 536194 353898
rect 541805 354454 542125 354486
rect 541805 354218 541847 354454
rect 542083 354218 542125 354454
rect 541805 354134 542125 354218
rect 541805 353898 541847 354134
rect 542083 353898 542125 354134
rect 541805 353866 542125 353898
rect 19910 345454 20230 345486
rect 19910 345218 19952 345454
rect 20188 345218 20230 345454
rect 19910 345134 20230 345218
rect 19910 344898 19952 345134
rect 20188 344898 20230 345134
rect 19910 344866 20230 344898
rect 25840 345454 26160 345486
rect 25840 345218 25882 345454
rect 26118 345218 26160 345454
rect 25840 345134 26160 345218
rect 25840 344898 25882 345134
rect 26118 344898 26160 345134
rect 25840 344866 26160 344898
rect 31771 345454 32091 345486
rect 31771 345218 31813 345454
rect 32049 345218 32091 345454
rect 31771 345134 32091 345218
rect 31771 344898 31813 345134
rect 32049 344898 32091 345134
rect 31771 344866 32091 344898
rect 46910 345454 47230 345486
rect 46910 345218 46952 345454
rect 47188 345218 47230 345454
rect 46910 345134 47230 345218
rect 46910 344898 46952 345134
rect 47188 344898 47230 345134
rect 46910 344866 47230 344898
rect 52840 345454 53160 345486
rect 52840 345218 52882 345454
rect 53118 345218 53160 345454
rect 52840 345134 53160 345218
rect 52840 344898 52882 345134
rect 53118 344898 53160 345134
rect 52840 344866 53160 344898
rect 58771 345454 59091 345486
rect 58771 345218 58813 345454
rect 59049 345218 59091 345454
rect 58771 345134 59091 345218
rect 58771 344898 58813 345134
rect 59049 344898 59091 345134
rect 58771 344866 59091 344898
rect 73910 345454 74230 345486
rect 73910 345218 73952 345454
rect 74188 345218 74230 345454
rect 73910 345134 74230 345218
rect 73910 344898 73952 345134
rect 74188 344898 74230 345134
rect 73910 344866 74230 344898
rect 79840 345454 80160 345486
rect 79840 345218 79882 345454
rect 80118 345218 80160 345454
rect 79840 345134 80160 345218
rect 79840 344898 79882 345134
rect 80118 344898 80160 345134
rect 79840 344866 80160 344898
rect 85771 345454 86091 345486
rect 85771 345218 85813 345454
rect 86049 345218 86091 345454
rect 85771 345134 86091 345218
rect 85771 344898 85813 345134
rect 86049 344898 86091 345134
rect 85771 344866 86091 344898
rect 100910 345454 101230 345486
rect 100910 345218 100952 345454
rect 101188 345218 101230 345454
rect 100910 345134 101230 345218
rect 100910 344898 100952 345134
rect 101188 344898 101230 345134
rect 100910 344866 101230 344898
rect 106840 345454 107160 345486
rect 106840 345218 106882 345454
rect 107118 345218 107160 345454
rect 106840 345134 107160 345218
rect 106840 344898 106882 345134
rect 107118 344898 107160 345134
rect 106840 344866 107160 344898
rect 112771 345454 113091 345486
rect 112771 345218 112813 345454
rect 113049 345218 113091 345454
rect 112771 345134 113091 345218
rect 112771 344898 112813 345134
rect 113049 344898 113091 345134
rect 112771 344866 113091 344898
rect 127910 345454 128230 345486
rect 127910 345218 127952 345454
rect 128188 345218 128230 345454
rect 127910 345134 128230 345218
rect 127910 344898 127952 345134
rect 128188 344898 128230 345134
rect 127910 344866 128230 344898
rect 133840 345454 134160 345486
rect 133840 345218 133882 345454
rect 134118 345218 134160 345454
rect 133840 345134 134160 345218
rect 133840 344898 133882 345134
rect 134118 344898 134160 345134
rect 133840 344866 134160 344898
rect 139771 345454 140091 345486
rect 139771 345218 139813 345454
rect 140049 345218 140091 345454
rect 139771 345134 140091 345218
rect 139771 344898 139813 345134
rect 140049 344898 140091 345134
rect 139771 344866 140091 344898
rect 154910 345454 155230 345486
rect 154910 345218 154952 345454
rect 155188 345218 155230 345454
rect 154910 345134 155230 345218
rect 154910 344898 154952 345134
rect 155188 344898 155230 345134
rect 154910 344866 155230 344898
rect 160840 345454 161160 345486
rect 160840 345218 160882 345454
rect 161118 345218 161160 345454
rect 160840 345134 161160 345218
rect 160840 344898 160882 345134
rect 161118 344898 161160 345134
rect 160840 344866 161160 344898
rect 166771 345454 167091 345486
rect 166771 345218 166813 345454
rect 167049 345218 167091 345454
rect 166771 345134 167091 345218
rect 166771 344898 166813 345134
rect 167049 344898 167091 345134
rect 166771 344866 167091 344898
rect 181910 345454 182230 345486
rect 181910 345218 181952 345454
rect 182188 345218 182230 345454
rect 181910 345134 182230 345218
rect 181910 344898 181952 345134
rect 182188 344898 182230 345134
rect 181910 344866 182230 344898
rect 187840 345454 188160 345486
rect 187840 345218 187882 345454
rect 188118 345218 188160 345454
rect 187840 345134 188160 345218
rect 187840 344898 187882 345134
rect 188118 344898 188160 345134
rect 187840 344866 188160 344898
rect 193771 345454 194091 345486
rect 193771 345218 193813 345454
rect 194049 345218 194091 345454
rect 193771 345134 194091 345218
rect 193771 344898 193813 345134
rect 194049 344898 194091 345134
rect 193771 344866 194091 344898
rect 208910 345454 209230 345486
rect 208910 345218 208952 345454
rect 209188 345218 209230 345454
rect 208910 345134 209230 345218
rect 208910 344898 208952 345134
rect 209188 344898 209230 345134
rect 208910 344866 209230 344898
rect 214840 345454 215160 345486
rect 214840 345218 214882 345454
rect 215118 345218 215160 345454
rect 214840 345134 215160 345218
rect 214840 344898 214882 345134
rect 215118 344898 215160 345134
rect 214840 344866 215160 344898
rect 220771 345454 221091 345486
rect 220771 345218 220813 345454
rect 221049 345218 221091 345454
rect 220771 345134 221091 345218
rect 220771 344898 220813 345134
rect 221049 344898 221091 345134
rect 220771 344866 221091 344898
rect 235910 345454 236230 345486
rect 235910 345218 235952 345454
rect 236188 345218 236230 345454
rect 235910 345134 236230 345218
rect 235910 344898 235952 345134
rect 236188 344898 236230 345134
rect 235910 344866 236230 344898
rect 241840 345454 242160 345486
rect 241840 345218 241882 345454
rect 242118 345218 242160 345454
rect 241840 345134 242160 345218
rect 241840 344898 241882 345134
rect 242118 344898 242160 345134
rect 241840 344866 242160 344898
rect 247771 345454 248091 345486
rect 247771 345218 247813 345454
rect 248049 345218 248091 345454
rect 247771 345134 248091 345218
rect 247771 344898 247813 345134
rect 248049 344898 248091 345134
rect 247771 344866 248091 344898
rect 262910 345454 263230 345486
rect 262910 345218 262952 345454
rect 263188 345218 263230 345454
rect 262910 345134 263230 345218
rect 262910 344898 262952 345134
rect 263188 344898 263230 345134
rect 262910 344866 263230 344898
rect 268840 345454 269160 345486
rect 268840 345218 268882 345454
rect 269118 345218 269160 345454
rect 268840 345134 269160 345218
rect 268840 344898 268882 345134
rect 269118 344898 269160 345134
rect 268840 344866 269160 344898
rect 274771 345454 275091 345486
rect 274771 345218 274813 345454
rect 275049 345218 275091 345454
rect 274771 345134 275091 345218
rect 274771 344898 274813 345134
rect 275049 344898 275091 345134
rect 274771 344866 275091 344898
rect 289910 345454 290230 345486
rect 289910 345218 289952 345454
rect 290188 345218 290230 345454
rect 289910 345134 290230 345218
rect 289910 344898 289952 345134
rect 290188 344898 290230 345134
rect 289910 344866 290230 344898
rect 295840 345454 296160 345486
rect 295840 345218 295882 345454
rect 296118 345218 296160 345454
rect 295840 345134 296160 345218
rect 295840 344898 295882 345134
rect 296118 344898 296160 345134
rect 295840 344866 296160 344898
rect 301771 345454 302091 345486
rect 301771 345218 301813 345454
rect 302049 345218 302091 345454
rect 301771 345134 302091 345218
rect 301771 344898 301813 345134
rect 302049 344898 302091 345134
rect 301771 344866 302091 344898
rect 316910 345454 317230 345486
rect 316910 345218 316952 345454
rect 317188 345218 317230 345454
rect 316910 345134 317230 345218
rect 316910 344898 316952 345134
rect 317188 344898 317230 345134
rect 316910 344866 317230 344898
rect 322840 345454 323160 345486
rect 322840 345218 322882 345454
rect 323118 345218 323160 345454
rect 322840 345134 323160 345218
rect 322840 344898 322882 345134
rect 323118 344898 323160 345134
rect 322840 344866 323160 344898
rect 328771 345454 329091 345486
rect 328771 345218 328813 345454
rect 329049 345218 329091 345454
rect 328771 345134 329091 345218
rect 328771 344898 328813 345134
rect 329049 344898 329091 345134
rect 328771 344866 329091 344898
rect 343910 345454 344230 345486
rect 343910 345218 343952 345454
rect 344188 345218 344230 345454
rect 343910 345134 344230 345218
rect 343910 344898 343952 345134
rect 344188 344898 344230 345134
rect 343910 344866 344230 344898
rect 349840 345454 350160 345486
rect 349840 345218 349882 345454
rect 350118 345218 350160 345454
rect 349840 345134 350160 345218
rect 349840 344898 349882 345134
rect 350118 344898 350160 345134
rect 349840 344866 350160 344898
rect 355771 345454 356091 345486
rect 355771 345218 355813 345454
rect 356049 345218 356091 345454
rect 355771 345134 356091 345218
rect 355771 344898 355813 345134
rect 356049 344898 356091 345134
rect 355771 344866 356091 344898
rect 370910 345454 371230 345486
rect 370910 345218 370952 345454
rect 371188 345218 371230 345454
rect 370910 345134 371230 345218
rect 370910 344898 370952 345134
rect 371188 344898 371230 345134
rect 370910 344866 371230 344898
rect 376840 345454 377160 345486
rect 376840 345218 376882 345454
rect 377118 345218 377160 345454
rect 376840 345134 377160 345218
rect 376840 344898 376882 345134
rect 377118 344898 377160 345134
rect 376840 344866 377160 344898
rect 382771 345454 383091 345486
rect 382771 345218 382813 345454
rect 383049 345218 383091 345454
rect 382771 345134 383091 345218
rect 382771 344898 382813 345134
rect 383049 344898 383091 345134
rect 382771 344866 383091 344898
rect 397910 345454 398230 345486
rect 397910 345218 397952 345454
rect 398188 345218 398230 345454
rect 397910 345134 398230 345218
rect 397910 344898 397952 345134
rect 398188 344898 398230 345134
rect 397910 344866 398230 344898
rect 403840 345454 404160 345486
rect 403840 345218 403882 345454
rect 404118 345218 404160 345454
rect 403840 345134 404160 345218
rect 403840 344898 403882 345134
rect 404118 344898 404160 345134
rect 403840 344866 404160 344898
rect 409771 345454 410091 345486
rect 409771 345218 409813 345454
rect 410049 345218 410091 345454
rect 409771 345134 410091 345218
rect 409771 344898 409813 345134
rect 410049 344898 410091 345134
rect 409771 344866 410091 344898
rect 424910 345454 425230 345486
rect 424910 345218 424952 345454
rect 425188 345218 425230 345454
rect 424910 345134 425230 345218
rect 424910 344898 424952 345134
rect 425188 344898 425230 345134
rect 424910 344866 425230 344898
rect 430840 345454 431160 345486
rect 430840 345218 430882 345454
rect 431118 345218 431160 345454
rect 430840 345134 431160 345218
rect 430840 344898 430882 345134
rect 431118 344898 431160 345134
rect 430840 344866 431160 344898
rect 436771 345454 437091 345486
rect 436771 345218 436813 345454
rect 437049 345218 437091 345454
rect 436771 345134 437091 345218
rect 436771 344898 436813 345134
rect 437049 344898 437091 345134
rect 436771 344866 437091 344898
rect 451910 345454 452230 345486
rect 451910 345218 451952 345454
rect 452188 345218 452230 345454
rect 451910 345134 452230 345218
rect 451910 344898 451952 345134
rect 452188 344898 452230 345134
rect 451910 344866 452230 344898
rect 457840 345454 458160 345486
rect 457840 345218 457882 345454
rect 458118 345218 458160 345454
rect 457840 345134 458160 345218
rect 457840 344898 457882 345134
rect 458118 344898 458160 345134
rect 457840 344866 458160 344898
rect 463771 345454 464091 345486
rect 463771 345218 463813 345454
rect 464049 345218 464091 345454
rect 463771 345134 464091 345218
rect 463771 344898 463813 345134
rect 464049 344898 464091 345134
rect 463771 344866 464091 344898
rect 478910 345454 479230 345486
rect 478910 345218 478952 345454
rect 479188 345218 479230 345454
rect 478910 345134 479230 345218
rect 478910 344898 478952 345134
rect 479188 344898 479230 345134
rect 478910 344866 479230 344898
rect 484840 345454 485160 345486
rect 484840 345218 484882 345454
rect 485118 345218 485160 345454
rect 484840 345134 485160 345218
rect 484840 344898 484882 345134
rect 485118 344898 485160 345134
rect 484840 344866 485160 344898
rect 490771 345454 491091 345486
rect 490771 345218 490813 345454
rect 491049 345218 491091 345454
rect 490771 345134 491091 345218
rect 490771 344898 490813 345134
rect 491049 344898 491091 345134
rect 490771 344866 491091 344898
rect 505910 345454 506230 345486
rect 505910 345218 505952 345454
rect 506188 345218 506230 345454
rect 505910 345134 506230 345218
rect 505910 344898 505952 345134
rect 506188 344898 506230 345134
rect 505910 344866 506230 344898
rect 511840 345454 512160 345486
rect 511840 345218 511882 345454
rect 512118 345218 512160 345454
rect 511840 345134 512160 345218
rect 511840 344898 511882 345134
rect 512118 344898 512160 345134
rect 511840 344866 512160 344898
rect 517771 345454 518091 345486
rect 517771 345218 517813 345454
rect 518049 345218 518091 345454
rect 517771 345134 518091 345218
rect 517771 344898 517813 345134
rect 518049 344898 518091 345134
rect 517771 344866 518091 344898
rect 532910 345454 533230 345486
rect 532910 345218 532952 345454
rect 533188 345218 533230 345454
rect 532910 345134 533230 345218
rect 532910 344898 532952 345134
rect 533188 344898 533230 345134
rect 532910 344866 533230 344898
rect 538840 345454 539160 345486
rect 538840 345218 538882 345454
rect 539118 345218 539160 345454
rect 538840 345134 539160 345218
rect 538840 344898 538882 345134
rect 539118 344898 539160 345134
rect 538840 344866 539160 344898
rect 544771 345454 545091 345486
rect 544771 345218 544813 345454
rect 545049 345218 545091 345454
rect 544771 345134 545091 345218
rect 544771 344898 544813 345134
rect 545049 344898 545091 345134
rect 544771 344866 545091 344898
rect 559794 345454 560414 362898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 318454 11414 335898
rect 19794 337394 20414 338000
rect 19794 337158 19826 337394
rect 20062 337158 20146 337394
rect 20382 337158 20414 337394
rect 19794 337074 20414 337158
rect 19794 336838 19826 337074
rect 20062 336838 20146 337074
rect 20382 336838 20414 337074
rect 19794 335000 20414 336838
rect 28794 336454 29414 338000
rect 28794 336218 28826 336454
rect 29062 336218 29146 336454
rect 29382 336218 29414 336454
rect 28794 336134 29414 336218
rect 28794 335898 28826 336134
rect 29062 335898 29146 336134
rect 29382 335898 29414 336134
rect 28794 335000 29414 335898
rect 37794 337394 38414 338000
rect 37794 337158 37826 337394
rect 38062 337158 38146 337394
rect 38382 337158 38414 337394
rect 37794 337074 38414 337158
rect 37794 336838 37826 337074
rect 38062 336838 38146 337074
rect 38382 336838 38414 337074
rect 37794 335000 38414 336838
rect 46794 336454 47414 338000
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 335000 47414 335898
rect 55794 337394 56414 338000
rect 55794 337158 55826 337394
rect 56062 337158 56146 337394
rect 56382 337158 56414 337394
rect 55794 337074 56414 337158
rect 55794 336838 55826 337074
rect 56062 336838 56146 337074
rect 56382 336838 56414 337074
rect 55794 335000 56414 336838
rect 64794 336454 65414 338000
rect 64794 336218 64826 336454
rect 65062 336218 65146 336454
rect 65382 336218 65414 336454
rect 64794 336134 65414 336218
rect 64794 335898 64826 336134
rect 65062 335898 65146 336134
rect 65382 335898 65414 336134
rect 64794 335000 65414 335898
rect 73794 337394 74414 338000
rect 73794 337158 73826 337394
rect 74062 337158 74146 337394
rect 74382 337158 74414 337394
rect 73794 337074 74414 337158
rect 73794 336838 73826 337074
rect 74062 336838 74146 337074
rect 74382 336838 74414 337074
rect 73794 335000 74414 336838
rect 82794 336454 83414 338000
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 335000 83414 335898
rect 91794 337394 92414 338000
rect 91794 337158 91826 337394
rect 92062 337158 92146 337394
rect 92382 337158 92414 337394
rect 91794 337074 92414 337158
rect 91794 336838 91826 337074
rect 92062 336838 92146 337074
rect 92382 336838 92414 337074
rect 91794 335000 92414 336838
rect 100794 336454 101414 338000
rect 100794 336218 100826 336454
rect 101062 336218 101146 336454
rect 101382 336218 101414 336454
rect 100794 336134 101414 336218
rect 100794 335898 100826 336134
rect 101062 335898 101146 336134
rect 101382 335898 101414 336134
rect 100794 335000 101414 335898
rect 109794 337394 110414 338000
rect 109794 337158 109826 337394
rect 110062 337158 110146 337394
rect 110382 337158 110414 337394
rect 109794 337074 110414 337158
rect 109794 336838 109826 337074
rect 110062 336838 110146 337074
rect 110382 336838 110414 337074
rect 109794 335000 110414 336838
rect 118794 336454 119414 338000
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 335000 119414 335898
rect 127794 337394 128414 338000
rect 127794 337158 127826 337394
rect 128062 337158 128146 337394
rect 128382 337158 128414 337394
rect 127794 337074 128414 337158
rect 127794 336838 127826 337074
rect 128062 336838 128146 337074
rect 128382 336838 128414 337074
rect 127794 335000 128414 336838
rect 136794 336454 137414 338000
rect 136794 336218 136826 336454
rect 137062 336218 137146 336454
rect 137382 336218 137414 336454
rect 136794 336134 137414 336218
rect 136794 335898 136826 336134
rect 137062 335898 137146 336134
rect 137382 335898 137414 336134
rect 136794 335000 137414 335898
rect 145794 337394 146414 338000
rect 145794 337158 145826 337394
rect 146062 337158 146146 337394
rect 146382 337158 146414 337394
rect 145794 337074 146414 337158
rect 145794 336838 145826 337074
rect 146062 336838 146146 337074
rect 146382 336838 146414 337074
rect 145794 335000 146414 336838
rect 154794 336454 155414 338000
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 335000 155414 335898
rect 163794 337394 164414 338000
rect 163794 337158 163826 337394
rect 164062 337158 164146 337394
rect 164382 337158 164414 337394
rect 163794 337074 164414 337158
rect 163794 336838 163826 337074
rect 164062 336838 164146 337074
rect 164382 336838 164414 337074
rect 163794 335000 164414 336838
rect 172794 336454 173414 338000
rect 172794 336218 172826 336454
rect 173062 336218 173146 336454
rect 173382 336218 173414 336454
rect 172794 336134 173414 336218
rect 172794 335898 172826 336134
rect 173062 335898 173146 336134
rect 173382 335898 173414 336134
rect 172794 335000 173414 335898
rect 181794 337394 182414 338000
rect 181794 337158 181826 337394
rect 182062 337158 182146 337394
rect 182382 337158 182414 337394
rect 181794 337074 182414 337158
rect 181794 336838 181826 337074
rect 182062 336838 182146 337074
rect 182382 336838 182414 337074
rect 181794 335000 182414 336838
rect 190794 336454 191414 338000
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 335000 191414 335898
rect 199794 337394 200414 338000
rect 199794 337158 199826 337394
rect 200062 337158 200146 337394
rect 200382 337158 200414 337394
rect 199794 337074 200414 337158
rect 199794 336838 199826 337074
rect 200062 336838 200146 337074
rect 200382 336838 200414 337074
rect 199794 335000 200414 336838
rect 208794 336454 209414 338000
rect 208794 336218 208826 336454
rect 209062 336218 209146 336454
rect 209382 336218 209414 336454
rect 208794 336134 209414 336218
rect 208794 335898 208826 336134
rect 209062 335898 209146 336134
rect 209382 335898 209414 336134
rect 208794 335000 209414 335898
rect 217794 337394 218414 338000
rect 217794 337158 217826 337394
rect 218062 337158 218146 337394
rect 218382 337158 218414 337394
rect 217794 337074 218414 337158
rect 217794 336838 217826 337074
rect 218062 336838 218146 337074
rect 218382 336838 218414 337074
rect 217794 335000 218414 336838
rect 226794 336454 227414 338000
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 335000 227414 335898
rect 235794 337394 236414 338000
rect 235794 337158 235826 337394
rect 236062 337158 236146 337394
rect 236382 337158 236414 337394
rect 235794 337074 236414 337158
rect 235794 336838 235826 337074
rect 236062 336838 236146 337074
rect 236382 336838 236414 337074
rect 235794 335000 236414 336838
rect 244794 336454 245414 338000
rect 244794 336218 244826 336454
rect 245062 336218 245146 336454
rect 245382 336218 245414 336454
rect 244794 336134 245414 336218
rect 244794 335898 244826 336134
rect 245062 335898 245146 336134
rect 245382 335898 245414 336134
rect 244794 335000 245414 335898
rect 253794 337394 254414 338000
rect 253794 337158 253826 337394
rect 254062 337158 254146 337394
rect 254382 337158 254414 337394
rect 253794 337074 254414 337158
rect 253794 336838 253826 337074
rect 254062 336838 254146 337074
rect 254382 336838 254414 337074
rect 253794 335000 254414 336838
rect 262794 336454 263414 338000
rect 262794 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 263414 336454
rect 262794 336134 263414 336218
rect 262794 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 263414 336134
rect 262794 335000 263414 335898
rect 271794 337394 272414 338000
rect 271794 337158 271826 337394
rect 272062 337158 272146 337394
rect 272382 337158 272414 337394
rect 271794 337074 272414 337158
rect 271794 336838 271826 337074
rect 272062 336838 272146 337074
rect 272382 336838 272414 337074
rect 271794 335000 272414 336838
rect 280794 336454 281414 338000
rect 280794 336218 280826 336454
rect 281062 336218 281146 336454
rect 281382 336218 281414 336454
rect 280794 336134 281414 336218
rect 280794 335898 280826 336134
rect 281062 335898 281146 336134
rect 281382 335898 281414 336134
rect 280794 335000 281414 335898
rect 289794 337394 290414 338000
rect 289794 337158 289826 337394
rect 290062 337158 290146 337394
rect 290382 337158 290414 337394
rect 289794 337074 290414 337158
rect 289794 336838 289826 337074
rect 290062 336838 290146 337074
rect 290382 336838 290414 337074
rect 289794 335000 290414 336838
rect 298794 336454 299414 338000
rect 298794 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 299414 336454
rect 298794 336134 299414 336218
rect 298794 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 299414 336134
rect 298794 335000 299414 335898
rect 307794 337394 308414 338000
rect 307794 337158 307826 337394
rect 308062 337158 308146 337394
rect 308382 337158 308414 337394
rect 307794 337074 308414 337158
rect 307794 336838 307826 337074
rect 308062 336838 308146 337074
rect 308382 336838 308414 337074
rect 307794 335000 308414 336838
rect 316794 336454 317414 338000
rect 316794 336218 316826 336454
rect 317062 336218 317146 336454
rect 317382 336218 317414 336454
rect 316794 336134 317414 336218
rect 316794 335898 316826 336134
rect 317062 335898 317146 336134
rect 317382 335898 317414 336134
rect 316794 335000 317414 335898
rect 325794 337394 326414 338000
rect 325794 337158 325826 337394
rect 326062 337158 326146 337394
rect 326382 337158 326414 337394
rect 325794 337074 326414 337158
rect 325794 336838 325826 337074
rect 326062 336838 326146 337074
rect 326382 336838 326414 337074
rect 325794 335000 326414 336838
rect 334794 336454 335414 338000
rect 334794 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 335414 336454
rect 334794 336134 335414 336218
rect 334794 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 335414 336134
rect 334794 335000 335414 335898
rect 343794 337394 344414 338000
rect 343794 337158 343826 337394
rect 344062 337158 344146 337394
rect 344382 337158 344414 337394
rect 343794 337074 344414 337158
rect 343794 336838 343826 337074
rect 344062 336838 344146 337074
rect 344382 336838 344414 337074
rect 343794 335000 344414 336838
rect 352794 336454 353414 338000
rect 352794 336218 352826 336454
rect 353062 336218 353146 336454
rect 353382 336218 353414 336454
rect 352794 336134 353414 336218
rect 352794 335898 352826 336134
rect 353062 335898 353146 336134
rect 353382 335898 353414 336134
rect 352794 335000 353414 335898
rect 361794 337394 362414 338000
rect 361794 337158 361826 337394
rect 362062 337158 362146 337394
rect 362382 337158 362414 337394
rect 361794 337074 362414 337158
rect 361794 336838 361826 337074
rect 362062 336838 362146 337074
rect 362382 336838 362414 337074
rect 361794 335000 362414 336838
rect 370794 336454 371414 338000
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 335000 371414 335898
rect 379794 337394 380414 338000
rect 379794 337158 379826 337394
rect 380062 337158 380146 337394
rect 380382 337158 380414 337394
rect 379794 337074 380414 337158
rect 379794 336838 379826 337074
rect 380062 336838 380146 337074
rect 380382 336838 380414 337074
rect 379794 335000 380414 336838
rect 388794 336454 389414 338000
rect 388794 336218 388826 336454
rect 389062 336218 389146 336454
rect 389382 336218 389414 336454
rect 388794 336134 389414 336218
rect 388794 335898 388826 336134
rect 389062 335898 389146 336134
rect 389382 335898 389414 336134
rect 388794 335000 389414 335898
rect 397794 337394 398414 338000
rect 397794 337158 397826 337394
rect 398062 337158 398146 337394
rect 398382 337158 398414 337394
rect 397794 337074 398414 337158
rect 397794 336838 397826 337074
rect 398062 336838 398146 337074
rect 398382 336838 398414 337074
rect 397794 335000 398414 336838
rect 406794 336454 407414 338000
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 335000 407414 335898
rect 415794 337394 416414 338000
rect 415794 337158 415826 337394
rect 416062 337158 416146 337394
rect 416382 337158 416414 337394
rect 415794 337074 416414 337158
rect 415794 336838 415826 337074
rect 416062 336838 416146 337074
rect 416382 336838 416414 337074
rect 415794 335000 416414 336838
rect 424794 336454 425414 338000
rect 424794 336218 424826 336454
rect 425062 336218 425146 336454
rect 425382 336218 425414 336454
rect 424794 336134 425414 336218
rect 424794 335898 424826 336134
rect 425062 335898 425146 336134
rect 425382 335898 425414 336134
rect 424794 335000 425414 335898
rect 433794 337394 434414 338000
rect 433794 337158 433826 337394
rect 434062 337158 434146 337394
rect 434382 337158 434414 337394
rect 433794 337074 434414 337158
rect 433794 336838 433826 337074
rect 434062 336838 434146 337074
rect 434382 336838 434414 337074
rect 433794 335000 434414 336838
rect 442794 336454 443414 338000
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 335000 443414 335898
rect 451794 337394 452414 338000
rect 451794 337158 451826 337394
rect 452062 337158 452146 337394
rect 452382 337158 452414 337394
rect 451794 337074 452414 337158
rect 451794 336838 451826 337074
rect 452062 336838 452146 337074
rect 452382 336838 452414 337074
rect 451794 335000 452414 336838
rect 460794 336454 461414 338000
rect 460794 336218 460826 336454
rect 461062 336218 461146 336454
rect 461382 336218 461414 336454
rect 460794 336134 461414 336218
rect 460794 335898 460826 336134
rect 461062 335898 461146 336134
rect 461382 335898 461414 336134
rect 460794 335000 461414 335898
rect 469794 337394 470414 338000
rect 469794 337158 469826 337394
rect 470062 337158 470146 337394
rect 470382 337158 470414 337394
rect 469794 337074 470414 337158
rect 469794 336838 469826 337074
rect 470062 336838 470146 337074
rect 470382 336838 470414 337074
rect 469794 335000 470414 336838
rect 478794 336454 479414 338000
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 335000 479414 335898
rect 487794 337394 488414 338000
rect 487794 337158 487826 337394
rect 488062 337158 488146 337394
rect 488382 337158 488414 337394
rect 487794 337074 488414 337158
rect 487794 336838 487826 337074
rect 488062 336838 488146 337074
rect 488382 336838 488414 337074
rect 487794 335000 488414 336838
rect 496794 336454 497414 338000
rect 496794 336218 496826 336454
rect 497062 336218 497146 336454
rect 497382 336218 497414 336454
rect 496794 336134 497414 336218
rect 496794 335898 496826 336134
rect 497062 335898 497146 336134
rect 497382 335898 497414 336134
rect 496794 335000 497414 335898
rect 505794 337394 506414 338000
rect 505794 337158 505826 337394
rect 506062 337158 506146 337394
rect 506382 337158 506414 337394
rect 505794 337074 506414 337158
rect 505794 336838 505826 337074
rect 506062 336838 506146 337074
rect 506382 336838 506414 337074
rect 505794 335000 506414 336838
rect 514794 336454 515414 338000
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 335000 515414 335898
rect 523794 337394 524414 338000
rect 523794 337158 523826 337394
rect 524062 337158 524146 337394
rect 524382 337158 524414 337394
rect 523794 337074 524414 337158
rect 523794 336838 523826 337074
rect 524062 336838 524146 337074
rect 524382 336838 524414 337074
rect 523794 335000 524414 336838
rect 532794 336454 533414 338000
rect 532794 336218 532826 336454
rect 533062 336218 533146 336454
rect 533382 336218 533414 336454
rect 532794 336134 533414 336218
rect 532794 335898 532826 336134
rect 533062 335898 533146 336134
rect 533382 335898 533414 336134
rect 532794 335000 533414 335898
rect 541794 337394 542414 338000
rect 541794 337158 541826 337394
rect 542062 337158 542146 337394
rect 542382 337158 542414 337394
rect 541794 337074 542414 337158
rect 541794 336838 541826 337074
rect 542062 336838 542146 337074
rect 542382 336838 542414 337074
rect 541794 335000 542414 336838
rect 550794 336454 551414 338000
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 335000 551414 335898
rect 19910 327454 20230 327486
rect 19910 327218 19952 327454
rect 20188 327218 20230 327454
rect 19910 327134 20230 327218
rect 19910 326898 19952 327134
rect 20188 326898 20230 327134
rect 19910 326866 20230 326898
rect 25840 327454 26160 327486
rect 25840 327218 25882 327454
rect 26118 327218 26160 327454
rect 25840 327134 26160 327218
rect 25840 326898 25882 327134
rect 26118 326898 26160 327134
rect 25840 326866 26160 326898
rect 31771 327454 32091 327486
rect 31771 327218 31813 327454
rect 32049 327218 32091 327454
rect 31771 327134 32091 327218
rect 31771 326898 31813 327134
rect 32049 326898 32091 327134
rect 31771 326866 32091 326898
rect 46910 327454 47230 327486
rect 46910 327218 46952 327454
rect 47188 327218 47230 327454
rect 46910 327134 47230 327218
rect 46910 326898 46952 327134
rect 47188 326898 47230 327134
rect 46910 326866 47230 326898
rect 52840 327454 53160 327486
rect 52840 327218 52882 327454
rect 53118 327218 53160 327454
rect 52840 327134 53160 327218
rect 52840 326898 52882 327134
rect 53118 326898 53160 327134
rect 52840 326866 53160 326898
rect 58771 327454 59091 327486
rect 58771 327218 58813 327454
rect 59049 327218 59091 327454
rect 58771 327134 59091 327218
rect 58771 326898 58813 327134
rect 59049 326898 59091 327134
rect 58771 326866 59091 326898
rect 73910 327454 74230 327486
rect 73910 327218 73952 327454
rect 74188 327218 74230 327454
rect 73910 327134 74230 327218
rect 73910 326898 73952 327134
rect 74188 326898 74230 327134
rect 73910 326866 74230 326898
rect 79840 327454 80160 327486
rect 79840 327218 79882 327454
rect 80118 327218 80160 327454
rect 79840 327134 80160 327218
rect 79840 326898 79882 327134
rect 80118 326898 80160 327134
rect 79840 326866 80160 326898
rect 85771 327454 86091 327486
rect 85771 327218 85813 327454
rect 86049 327218 86091 327454
rect 85771 327134 86091 327218
rect 85771 326898 85813 327134
rect 86049 326898 86091 327134
rect 85771 326866 86091 326898
rect 100910 327454 101230 327486
rect 100910 327218 100952 327454
rect 101188 327218 101230 327454
rect 100910 327134 101230 327218
rect 100910 326898 100952 327134
rect 101188 326898 101230 327134
rect 100910 326866 101230 326898
rect 106840 327454 107160 327486
rect 106840 327218 106882 327454
rect 107118 327218 107160 327454
rect 106840 327134 107160 327218
rect 106840 326898 106882 327134
rect 107118 326898 107160 327134
rect 106840 326866 107160 326898
rect 112771 327454 113091 327486
rect 112771 327218 112813 327454
rect 113049 327218 113091 327454
rect 112771 327134 113091 327218
rect 112771 326898 112813 327134
rect 113049 326898 113091 327134
rect 112771 326866 113091 326898
rect 127910 327454 128230 327486
rect 127910 327218 127952 327454
rect 128188 327218 128230 327454
rect 127910 327134 128230 327218
rect 127910 326898 127952 327134
rect 128188 326898 128230 327134
rect 127910 326866 128230 326898
rect 133840 327454 134160 327486
rect 133840 327218 133882 327454
rect 134118 327218 134160 327454
rect 133840 327134 134160 327218
rect 133840 326898 133882 327134
rect 134118 326898 134160 327134
rect 133840 326866 134160 326898
rect 139771 327454 140091 327486
rect 139771 327218 139813 327454
rect 140049 327218 140091 327454
rect 139771 327134 140091 327218
rect 139771 326898 139813 327134
rect 140049 326898 140091 327134
rect 139771 326866 140091 326898
rect 154910 327454 155230 327486
rect 154910 327218 154952 327454
rect 155188 327218 155230 327454
rect 154910 327134 155230 327218
rect 154910 326898 154952 327134
rect 155188 326898 155230 327134
rect 154910 326866 155230 326898
rect 160840 327454 161160 327486
rect 160840 327218 160882 327454
rect 161118 327218 161160 327454
rect 160840 327134 161160 327218
rect 160840 326898 160882 327134
rect 161118 326898 161160 327134
rect 160840 326866 161160 326898
rect 166771 327454 167091 327486
rect 166771 327218 166813 327454
rect 167049 327218 167091 327454
rect 166771 327134 167091 327218
rect 166771 326898 166813 327134
rect 167049 326898 167091 327134
rect 166771 326866 167091 326898
rect 181910 327454 182230 327486
rect 181910 327218 181952 327454
rect 182188 327218 182230 327454
rect 181910 327134 182230 327218
rect 181910 326898 181952 327134
rect 182188 326898 182230 327134
rect 181910 326866 182230 326898
rect 187840 327454 188160 327486
rect 187840 327218 187882 327454
rect 188118 327218 188160 327454
rect 187840 327134 188160 327218
rect 187840 326898 187882 327134
rect 188118 326898 188160 327134
rect 187840 326866 188160 326898
rect 193771 327454 194091 327486
rect 193771 327218 193813 327454
rect 194049 327218 194091 327454
rect 193771 327134 194091 327218
rect 193771 326898 193813 327134
rect 194049 326898 194091 327134
rect 193771 326866 194091 326898
rect 208910 327454 209230 327486
rect 208910 327218 208952 327454
rect 209188 327218 209230 327454
rect 208910 327134 209230 327218
rect 208910 326898 208952 327134
rect 209188 326898 209230 327134
rect 208910 326866 209230 326898
rect 214840 327454 215160 327486
rect 214840 327218 214882 327454
rect 215118 327218 215160 327454
rect 214840 327134 215160 327218
rect 214840 326898 214882 327134
rect 215118 326898 215160 327134
rect 214840 326866 215160 326898
rect 220771 327454 221091 327486
rect 220771 327218 220813 327454
rect 221049 327218 221091 327454
rect 220771 327134 221091 327218
rect 220771 326898 220813 327134
rect 221049 326898 221091 327134
rect 220771 326866 221091 326898
rect 235910 327454 236230 327486
rect 235910 327218 235952 327454
rect 236188 327218 236230 327454
rect 235910 327134 236230 327218
rect 235910 326898 235952 327134
rect 236188 326898 236230 327134
rect 235910 326866 236230 326898
rect 241840 327454 242160 327486
rect 241840 327218 241882 327454
rect 242118 327218 242160 327454
rect 241840 327134 242160 327218
rect 241840 326898 241882 327134
rect 242118 326898 242160 327134
rect 241840 326866 242160 326898
rect 247771 327454 248091 327486
rect 247771 327218 247813 327454
rect 248049 327218 248091 327454
rect 247771 327134 248091 327218
rect 247771 326898 247813 327134
rect 248049 326898 248091 327134
rect 247771 326866 248091 326898
rect 262910 327454 263230 327486
rect 262910 327218 262952 327454
rect 263188 327218 263230 327454
rect 262910 327134 263230 327218
rect 262910 326898 262952 327134
rect 263188 326898 263230 327134
rect 262910 326866 263230 326898
rect 268840 327454 269160 327486
rect 268840 327218 268882 327454
rect 269118 327218 269160 327454
rect 268840 327134 269160 327218
rect 268840 326898 268882 327134
rect 269118 326898 269160 327134
rect 268840 326866 269160 326898
rect 274771 327454 275091 327486
rect 274771 327218 274813 327454
rect 275049 327218 275091 327454
rect 274771 327134 275091 327218
rect 274771 326898 274813 327134
rect 275049 326898 275091 327134
rect 274771 326866 275091 326898
rect 289910 327454 290230 327486
rect 289910 327218 289952 327454
rect 290188 327218 290230 327454
rect 289910 327134 290230 327218
rect 289910 326898 289952 327134
rect 290188 326898 290230 327134
rect 289910 326866 290230 326898
rect 295840 327454 296160 327486
rect 295840 327218 295882 327454
rect 296118 327218 296160 327454
rect 295840 327134 296160 327218
rect 295840 326898 295882 327134
rect 296118 326898 296160 327134
rect 295840 326866 296160 326898
rect 301771 327454 302091 327486
rect 301771 327218 301813 327454
rect 302049 327218 302091 327454
rect 301771 327134 302091 327218
rect 301771 326898 301813 327134
rect 302049 326898 302091 327134
rect 301771 326866 302091 326898
rect 316910 327454 317230 327486
rect 316910 327218 316952 327454
rect 317188 327218 317230 327454
rect 316910 327134 317230 327218
rect 316910 326898 316952 327134
rect 317188 326898 317230 327134
rect 316910 326866 317230 326898
rect 322840 327454 323160 327486
rect 322840 327218 322882 327454
rect 323118 327218 323160 327454
rect 322840 327134 323160 327218
rect 322840 326898 322882 327134
rect 323118 326898 323160 327134
rect 322840 326866 323160 326898
rect 328771 327454 329091 327486
rect 328771 327218 328813 327454
rect 329049 327218 329091 327454
rect 328771 327134 329091 327218
rect 328771 326898 328813 327134
rect 329049 326898 329091 327134
rect 328771 326866 329091 326898
rect 343910 327454 344230 327486
rect 343910 327218 343952 327454
rect 344188 327218 344230 327454
rect 343910 327134 344230 327218
rect 343910 326898 343952 327134
rect 344188 326898 344230 327134
rect 343910 326866 344230 326898
rect 349840 327454 350160 327486
rect 349840 327218 349882 327454
rect 350118 327218 350160 327454
rect 349840 327134 350160 327218
rect 349840 326898 349882 327134
rect 350118 326898 350160 327134
rect 349840 326866 350160 326898
rect 355771 327454 356091 327486
rect 355771 327218 355813 327454
rect 356049 327218 356091 327454
rect 355771 327134 356091 327218
rect 355771 326898 355813 327134
rect 356049 326898 356091 327134
rect 355771 326866 356091 326898
rect 370910 327454 371230 327486
rect 370910 327218 370952 327454
rect 371188 327218 371230 327454
rect 370910 327134 371230 327218
rect 370910 326898 370952 327134
rect 371188 326898 371230 327134
rect 370910 326866 371230 326898
rect 376840 327454 377160 327486
rect 376840 327218 376882 327454
rect 377118 327218 377160 327454
rect 376840 327134 377160 327218
rect 376840 326898 376882 327134
rect 377118 326898 377160 327134
rect 376840 326866 377160 326898
rect 382771 327454 383091 327486
rect 382771 327218 382813 327454
rect 383049 327218 383091 327454
rect 382771 327134 383091 327218
rect 382771 326898 382813 327134
rect 383049 326898 383091 327134
rect 382771 326866 383091 326898
rect 397910 327454 398230 327486
rect 397910 327218 397952 327454
rect 398188 327218 398230 327454
rect 397910 327134 398230 327218
rect 397910 326898 397952 327134
rect 398188 326898 398230 327134
rect 397910 326866 398230 326898
rect 403840 327454 404160 327486
rect 403840 327218 403882 327454
rect 404118 327218 404160 327454
rect 403840 327134 404160 327218
rect 403840 326898 403882 327134
rect 404118 326898 404160 327134
rect 403840 326866 404160 326898
rect 409771 327454 410091 327486
rect 409771 327218 409813 327454
rect 410049 327218 410091 327454
rect 409771 327134 410091 327218
rect 409771 326898 409813 327134
rect 410049 326898 410091 327134
rect 409771 326866 410091 326898
rect 424910 327454 425230 327486
rect 424910 327218 424952 327454
rect 425188 327218 425230 327454
rect 424910 327134 425230 327218
rect 424910 326898 424952 327134
rect 425188 326898 425230 327134
rect 424910 326866 425230 326898
rect 430840 327454 431160 327486
rect 430840 327218 430882 327454
rect 431118 327218 431160 327454
rect 430840 327134 431160 327218
rect 430840 326898 430882 327134
rect 431118 326898 431160 327134
rect 430840 326866 431160 326898
rect 436771 327454 437091 327486
rect 436771 327218 436813 327454
rect 437049 327218 437091 327454
rect 436771 327134 437091 327218
rect 436771 326898 436813 327134
rect 437049 326898 437091 327134
rect 436771 326866 437091 326898
rect 451910 327454 452230 327486
rect 451910 327218 451952 327454
rect 452188 327218 452230 327454
rect 451910 327134 452230 327218
rect 451910 326898 451952 327134
rect 452188 326898 452230 327134
rect 451910 326866 452230 326898
rect 457840 327454 458160 327486
rect 457840 327218 457882 327454
rect 458118 327218 458160 327454
rect 457840 327134 458160 327218
rect 457840 326898 457882 327134
rect 458118 326898 458160 327134
rect 457840 326866 458160 326898
rect 463771 327454 464091 327486
rect 463771 327218 463813 327454
rect 464049 327218 464091 327454
rect 463771 327134 464091 327218
rect 463771 326898 463813 327134
rect 464049 326898 464091 327134
rect 463771 326866 464091 326898
rect 478910 327454 479230 327486
rect 478910 327218 478952 327454
rect 479188 327218 479230 327454
rect 478910 327134 479230 327218
rect 478910 326898 478952 327134
rect 479188 326898 479230 327134
rect 478910 326866 479230 326898
rect 484840 327454 485160 327486
rect 484840 327218 484882 327454
rect 485118 327218 485160 327454
rect 484840 327134 485160 327218
rect 484840 326898 484882 327134
rect 485118 326898 485160 327134
rect 484840 326866 485160 326898
rect 490771 327454 491091 327486
rect 490771 327218 490813 327454
rect 491049 327218 491091 327454
rect 490771 327134 491091 327218
rect 490771 326898 490813 327134
rect 491049 326898 491091 327134
rect 490771 326866 491091 326898
rect 505910 327454 506230 327486
rect 505910 327218 505952 327454
rect 506188 327218 506230 327454
rect 505910 327134 506230 327218
rect 505910 326898 505952 327134
rect 506188 326898 506230 327134
rect 505910 326866 506230 326898
rect 511840 327454 512160 327486
rect 511840 327218 511882 327454
rect 512118 327218 512160 327454
rect 511840 327134 512160 327218
rect 511840 326898 511882 327134
rect 512118 326898 512160 327134
rect 511840 326866 512160 326898
rect 517771 327454 518091 327486
rect 517771 327218 517813 327454
rect 518049 327218 518091 327454
rect 517771 327134 518091 327218
rect 517771 326898 517813 327134
rect 518049 326898 518091 327134
rect 517771 326866 518091 326898
rect 532910 327454 533230 327486
rect 532910 327218 532952 327454
rect 533188 327218 533230 327454
rect 532910 327134 533230 327218
rect 532910 326898 532952 327134
rect 533188 326898 533230 327134
rect 532910 326866 533230 326898
rect 538840 327454 539160 327486
rect 538840 327218 538882 327454
rect 539118 327218 539160 327454
rect 538840 327134 539160 327218
rect 538840 326898 538882 327134
rect 539118 326898 539160 327134
rect 538840 326866 539160 326898
rect 544771 327454 545091 327486
rect 544771 327218 544813 327454
rect 545049 327218 545091 327454
rect 544771 327134 545091 327218
rect 544771 326898 544813 327134
rect 545049 326898 545091 327134
rect 544771 326866 545091 326898
rect 559794 327454 560414 344898
rect 559794 327218 559826 327454
rect 560062 327218 560146 327454
rect 560382 327218 560414 327454
rect 559794 327134 560414 327218
rect 559794 326898 559826 327134
rect 560062 326898 560146 327134
rect 560382 326898 560414 327134
rect 10794 318218 10826 318454
rect 11062 318218 11146 318454
rect 11382 318218 11414 318454
rect 10794 318134 11414 318218
rect 10794 317898 10826 318134
rect 11062 317898 11146 318134
rect 11382 317898 11414 318134
rect 10794 300454 11414 317898
rect 22874 318454 23194 318486
rect 22874 318218 22916 318454
rect 23152 318218 23194 318454
rect 22874 318134 23194 318218
rect 22874 317898 22916 318134
rect 23152 317898 23194 318134
rect 22874 317866 23194 317898
rect 28805 318454 29125 318486
rect 28805 318218 28847 318454
rect 29083 318218 29125 318454
rect 28805 318134 29125 318218
rect 28805 317898 28847 318134
rect 29083 317898 29125 318134
rect 28805 317866 29125 317898
rect 49874 318454 50194 318486
rect 49874 318218 49916 318454
rect 50152 318218 50194 318454
rect 49874 318134 50194 318218
rect 49874 317898 49916 318134
rect 50152 317898 50194 318134
rect 49874 317866 50194 317898
rect 55805 318454 56125 318486
rect 55805 318218 55847 318454
rect 56083 318218 56125 318454
rect 55805 318134 56125 318218
rect 55805 317898 55847 318134
rect 56083 317898 56125 318134
rect 55805 317866 56125 317898
rect 76874 318454 77194 318486
rect 76874 318218 76916 318454
rect 77152 318218 77194 318454
rect 76874 318134 77194 318218
rect 76874 317898 76916 318134
rect 77152 317898 77194 318134
rect 76874 317866 77194 317898
rect 82805 318454 83125 318486
rect 82805 318218 82847 318454
rect 83083 318218 83125 318454
rect 82805 318134 83125 318218
rect 82805 317898 82847 318134
rect 83083 317898 83125 318134
rect 82805 317866 83125 317898
rect 103874 318454 104194 318486
rect 103874 318218 103916 318454
rect 104152 318218 104194 318454
rect 103874 318134 104194 318218
rect 103874 317898 103916 318134
rect 104152 317898 104194 318134
rect 103874 317866 104194 317898
rect 109805 318454 110125 318486
rect 109805 318218 109847 318454
rect 110083 318218 110125 318454
rect 109805 318134 110125 318218
rect 109805 317898 109847 318134
rect 110083 317898 110125 318134
rect 109805 317866 110125 317898
rect 130874 318454 131194 318486
rect 130874 318218 130916 318454
rect 131152 318218 131194 318454
rect 130874 318134 131194 318218
rect 130874 317898 130916 318134
rect 131152 317898 131194 318134
rect 130874 317866 131194 317898
rect 136805 318454 137125 318486
rect 136805 318218 136847 318454
rect 137083 318218 137125 318454
rect 136805 318134 137125 318218
rect 136805 317898 136847 318134
rect 137083 317898 137125 318134
rect 136805 317866 137125 317898
rect 157874 318454 158194 318486
rect 157874 318218 157916 318454
rect 158152 318218 158194 318454
rect 157874 318134 158194 318218
rect 157874 317898 157916 318134
rect 158152 317898 158194 318134
rect 157874 317866 158194 317898
rect 163805 318454 164125 318486
rect 163805 318218 163847 318454
rect 164083 318218 164125 318454
rect 163805 318134 164125 318218
rect 163805 317898 163847 318134
rect 164083 317898 164125 318134
rect 163805 317866 164125 317898
rect 184874 318454 185194 318486
rect 184874 318218 184916 318454
rect 185152 318218 185194 318454
rect 184874 318134 185194 318218
rect 184874 317898 184916 318134
rect 185152 317898 185194 318134
rect 184874 317866 185194 317898
rect 190805 318454 191125 318486
rect 190805 318218 190847 318454
rect 191083 318218 191125 318454
rect 190805 318134 191125 318218
rect 190805 317898 190847 318134
rect 191083 317898 191125 318134
rect 190805 317866 191125 317898
rect 211874 318454 212194 318486
rect 211874 318218 211916 318454
rect 212152 318218 212194 318454
rect 211874 318134 212194 318218
rect 211874 317898 211916 318134
rect 212152 317898 212194 318134
rect 211874 317866 212194 317898
rect 217805 318454 218125 318486
rect 217805 318218 217847 318454
rect 218083 318218 218125 318454
rect 217805 318134 218125 318218
rect 217805 317898 217847 318134
rect 218083 317898 218125 318134
rect 217805 317866 218125 317898
rect 238874 318454 239194 318486
rect 238874 318218 238916 318454
rect 239152 318218 239194 318454
rect 238874 318134 239194 318218
rect 238874 317898 238916 318134
rect 239152 317898 239194 318134
rect 238874 317866 239194 317898
rect 244805 318454 245125 318486
rect 244805 318218 244847 318454
rect 245083 318218 245125 318454
rect 244805 318134 245125 318218
rect 244805 317898 244847 318134
rect 245083 317898 245125 318134
rect 244805 317866 245125 317898
rect 265874 318454 266194 318486
rect 265874 318218 265916 318454
rect 266152 318218 266194 318454
rect 265874 318134 266194 318218
rect 265874 317898 265916 318134
rect 266152 317898 266194 318134
rect 265874 317866 266194 317898
rect 271805 318454 272125 318486
rect 271805 318218 271847 318454
rect 272083 318218 272125 318454
rect 271805 318134 272125 318218
rect 271805 317898 271847 318134
rect 272083 317898 272125 318134
rect 271805 317866 272125 317898
rect 292874 318454 293194 318486
rect 292874 318218 292916 318454
rect 293152 318218 293194 318454
rect 292874 318134 293194 318218
rect 292874 317898 292916 318134
rect 293152 317898 293194 318134
rect 292874 317866 293194 317898
rect 298805 318454 299125 318486
rect 298805 318218 298847 318454
rect 299083 318218 299125 318454
rect 298805 318134 299125 318218
rect 298805 317898 298847 318134
rect 299083 317898 299125 318134
rect 298805 317866 299125 317898
rect 319874 318454 320194 318486
rect 319874 318218 319916 318454
rect 320152 318218 320194 318454
rect 319874 318134 320194 318218
rect 319874 317898 319916 318134
rect 320152 317898 320194 318134
rect 319874 317866 320194 317898
rect 325805 318454 326125 318486
rect 325805 318218 325847 318454
rect 326083 318218 326125 318454
rect 325805 318134 326125 318218
rect 325805 317898 325847 318134
rect 326083 317898 326125 318134
rect 325805 317866 326125 317898
rect 346874 318454 347194 318486
rect 346874 318218 346916 318454
rect 347152 318218 347194 318454
rect 346874 318134 347194 318218
rect 346874 317898 346916 318134
rect 347152 317898 347194 318134
rect 346874 317866 347194 317898
rect 352805 318454 353125 318486
rect 352805 318218 352847 318454
rect 353083 318218 353125 318454
rect 352805 318134 353125 318218
rect 352805 317898 352847 318134
rect 353083 317898 353125 318134
rect 352805 317866 353125 317898
rect 373874 318454 374194 318486
rect 373874 318218 373916 318454
rect 374152 318218 374194 318454
rect 373874 318134 374194 318218
rect 373874 317898 373916 318134
rect 374152 317898 374194 318134
rect 373874 317866 374194 317898
rect 379805 318454 380125 318486
rect 379805 318218 379847 318454
rect 380083 318218 380125 318454
rect 379805 318134 380125 318218
rect 379805 317898 379847 318134
rect 380083 317898 380125 318134
rect 379805 317866 380125 317898
rect 400874 318454 401194 318486
rect 400874 318218 400916 318454
rect 401152 318218 401194 318454
rect 400874 318134 401194 318218
rect 400874 317898 400916 318134
rect 401152 317898 401194 318134
rect 400874 317866 401194 317898
rect 406805 318454 407125 318486
rect 406805 318218 406847 318454
rect 407083 318218 407125 318454
rect 406805 318134 407125 318218
rect 406805 317898 406847 318134
rect 407083 317898 407125 318134
rect 406805 317866 407125 317898
rect 427874 318454 428194 318486
rect 427874 318218 427916 318454
rect 428152 318218 428194 318454
rect 427874 318134 428194 318218
rect 427874 317898 427916 318134
rect 428152 317898 428194 318134
rect 427874 317866 428194 317898
rect 433805 318454 434125 318486
rect 433805 318218 433847 318454
rect 434083 318218 434125 318454
rect 433805 318134 434125 318218
rect 433805 317898 433847 318134
rect 434083 317898 434125 318134
rect 433805 317866 434125 317898
rect 454874 318454 455194 318486
rect 454874 318218 454916 318454
rect 455152 318218 455194 318454
rect 454874 318134 455194 318218
rect 454874 317898 454916 318134
rect 455152 317898 455194 318134
rect 454874 317866 455194 317898
rect 460805 318454 461125 318486
rect 460805 318218 460847 318454
rect 461083 318218 461125 318454
rect 460805 318134 461125 318218
rect 460805 317898 460847 318134
rect 461083 317898 461125 318134
rect 460805 317866 461125 317898
rect 481874 318454 482194 318486
rect 481874 318218 481916 318454
rect 482152 318218 482194 318454
rect 481874 318134 482194 318218
rect 481874 317898 481916 318134
rect 482152 317898 482194 318134
rect 481874 317866 482194 317898
rect 487805 318454 488125 318486
rect 487805 318218 487847 318454
rect 488083 318218 488125 318454
rect 487805 318134 488125 318218
rect 487805 317898 487847 318134
rect 488083 317898 488125 318134
rect 487805 317866 488125 317898
rect 508874 318454 509194 318486
rect 508874 318218 508916 318454
rect 509152 318218 509194 318454
rect 508874 318134 509194 318218
rect 508874 317898 508916 318134
rect 509152 317898 509194 318134
rect 508874 317866 509194 317898
rect 514805 318454 515125 318486
rect 514805 318218 514847 318454
rect 515083 318218 515125 318454
rect 514805 318134 515125 318218
rect 514805 317898 514847 318134
rect 515083 317898 515125 318134
rect 514805 317866 515125 317898
rect 535874 318454 536194 318486
rect 535874 318218 535916 318454
rect 536152 318218 536194 318454
rect 535874 318134 536194 318218
rect 535874 317898 535916 318134
rect 536152 317898 536194 318134
rect 535874 317866 536194 317898
rect 541805 318454 542125 318486
rect 541805 318218 541847 318454
rect 542083 318218 542125 318454
rect 541805 318134 542125 318218
rect 541805 317898 541847 318134
rect 542083 317898 542125 318134
rect 541805 317866 542125 317898
rect 19794 309454 20414 311000
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 308000 20414 308898
rect 28794 310394 29414 311000
rect 28794 310158 28826 310394
rect 29062 310158 29146 310394
rect 29382 310158 29414 310394
rect 28794 310074 29414 310158
rect 28794 309838 28826 310074
rect 29062 309838 29146 310074
rect 29382 309838 29414 310074
rect 28794 308000 29414 309838
rect 37794 309454 38414 311000
rect 37794 309218 37826 309454
rect 38062 309218 38146 309454
rect 38382 309218 38414 309454
rect 37794 309134 38414 309218
rect 37794 308898 37826 309134
rect 38062 308898 38146 309134
rect 38382 308898 38414 309134
rect 37794 308000 38414 308898
rect 46794 310394 47414 311000
rect 46794 310158 46826 310394
rect 47062 310158 47146 310394
rect 47382 310158 47414 310394
rect 46794 310074 47414 310158
rect 46794 309838 46826 310074
rect 47062 309838 47146 310074
rect 47382 309838 47414 310074
rect 46794 308000 47414 309838
rect 55794 309454 56414 311000
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 308000 56414 308898
rect 64794 310394 65414 311000
rect 64794 310158 64826 310394
rect 65062 310158 65146 310394
rect 65382 310158 65414 310394
rect 64794 310074 65414 310158
rect 64794 309838 64826 310074
rect 65062 309838 65146 310074
rect 65382 309838 65414 310074
rect 64794 308000 65414 309838
rect 73794 309454 74414 311000
rect 73794 309218 73826 309454
rect 74062 309218 74146 309454
rect 74382 309218 74414 309454
rect 73794 309134 74414 309218
rect 73794 308898 73826 309134
rect 74062 308898 74146 309134
rect 74382 308898 74414 309134
rect 73794 308000 74414 308898
rect 82794 310394 83414 311000
rect 82794 310158 82826 310394
rect 83062 310158 83146 310394
rect 83382 310158 83414 310394
rect 82794 310074 83414 310158
rect 82794 309838 82826 310074
rect 83062 309838 83146 310074
rect 83382 309838 83414 310074
rect 82794 308000 83414 309838
rect 91794 309454 92414 311000
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 308000 92414 308898
rect 100794 310394 101414 311000
rect 100794 310158 100826 310394
rect 101062 310158 101146 310394
rect 101382 310158 101414 310394
rect 100794 310074 101414 310158
rect 100794 309838 100826 310074
rect 101062 309838 101146 310074
rect 101382 309838 101414 310074
rect 100794 308000 101414 309838
rect 109794 309454 110414 311000
rect 109794 309218 109826 309454
rect 110062 309218 110146 309454
rect 110382 309218 110414 309454
rect 109794 309134 110414 309218
rect 109794 308898 109826 309134
rect 110062 308898 110146 309134
rect 110382 308898 110414 309134
rect 109794 308000 110414 308898
rect 118794 310394 119414 311000
rect 118794 310158 118826 310394
rect 119062 310158 119146 310394
rect 119382 310158 119414 310394
rect 118794 310074 119414 310158
rect 118794 309838 118826 310074
rect 119062 309838 119146 310074
rect 119382 309838 119414 310074
rect 118794 308000 119414 309838
rect 127794 309454 128414 311000
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 308000 128414 308898
rect 136794 310394 137414 311000
rect 136794 310158 136826 310394
rect 137062 310158 137146 310394
rect 137382 310158 137414 310394
rect 136794 310074 137414 310158
rect 136794 309838 136826 310074
rect 137062 309838 137146 310074
rect 137382 309838 137414 310074
rect 136794 308000 137414 309838
rect 145794 309454 146414 311000
rect 145794 309218 145826 309454
rect 146062 309218 146146 309454
rect 146382 309218 146414 309454
rect 145794 309134 146414 309218
rect 145794 308898 145826 309134
rect 146062 308898 146146 309134
rect 146382 308898 146414 309134
rect 145794 308000 146414 308898
rect 154794 310394 155414 311000
rect 154794 310158 154826 310394
rect 155062 310158 155146 310394
rect 155382 310158 155414 310394
rect 154794 310074 155414 310158
rect 154794 309838 154826 310074
rect 155062 309838 155146 310074
rect 155382 309838 155414 310074
rect 154794 308000 155414 309838
rect 163794 309454 164414 311000
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 308000 164414 308898
rect 172794 310394 173414 311000
rect 172794 310158 172826 310394
rect 173062 310158 173146 310394
rect 173382 310158 173414 310394
rect 172794 310074 173414 310158
rect 172794 309838 172826 310074
rect 173062 309838 173146 310074
rect 173382 309838 173414 310074
rect 172794 308000 173414 309838
rect 181794 309454 182414 311000
rect 181794 309218 181826 309454
rect 182062 309218 182146 309454
rect 182382 309218 182414 309454
rect 181794 309134 182414 309218
rect 181794 308898 181826 309134
rect 182062 308898 182146 309134
rect 182382 308898 182414 309134
rect 181794 308000 182414 308898
rect 190794 310394 191414 311000
rect 190794 310158 190826 310394
rect 191062 310158 191146 310394
rect 191382 310158 191414 310394
rect 190794 310074 191414 310158
rect 190794 309838 190826 310074
rect 191062 309838 191146 310074
rect 191382 309838 191414 310074
rect 190794 308000 191414 309838
rect 199794 309454 200414 311000
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 308000 200414 308898
rect 208794 310394 209414 311000
rect 208794 310158 208826 310394
rect 209062 310158 209146 310394
rect 209382 310158 209414 310394
rect 208794 310074 209414 310158
rect 208794 309838 208826 310074
rect 209062 309838 209146 310074
rect 209382 309838 209414 310074
rect 208794 308000 209414 309838
rect 217794 309454 218414 311000
rect 217794 309218 217826 309454
rect 218062 309218 218146 309454
rect 218382 309218 218414 309454
rect 217794 309134 218414 309218
rect 217794 308898 217826 309134
rect 218062 308898 218146 309134
rect 218382 308898 218414 309134
rect 217794 308000 218414 308898
rect 226794 310394 227414 311000
rect 226794 310158 226826 310394
rect 227062 310158 227146 310394
rect 227382 310158 227414 310394
rect 226794 310074 227414 310158
rect 226794 309838 226826 310074
rect 227062 309838 227146 310074
rect 227382 309838 227414 310074
rect 226794 308000 227414 309838
rect 235794 309454 236414 311000
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 308000 236414 308898
rect 244794 310394 245414 311000
rect 244794 310158 244826 310394
rect 245062 310158 245146 310394
rect 245382 310158 245414 310394
rect 244794 310074 245414 310158
rect 244794 309838 244826 310074
rect 245062 309838 245146 310074
rect 245382 309838 245414 310074
rect 244794 308000 245414 309838
rect 253794 309454 254414 311000
rect 253794 309218 253826 309454
rect 254062 309218 254146 309454
rect 254382 309218 254414 309454
rect 253794 309134 254414 309218
rect 253794 308898 253826 309134
rect 254062 308898 254146 309134
rect 254382 308898 254414 309134
rect 253794 308000 254414 308898
rect 262794 310394 263414 311000
rect 262794 310158 262826 310394
rect 263062 310158 263146 310394
rect 263382 310158 263414 310394
rect 262794 310074 263414 310158
rect 262794 309838 262826 310074
rect 263062 309838 263146 310074
rect 263382 309838 263414 310074
rect 262794 308000 263414 309838
rect 271794 309454 272414 311000
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 308000 272414 308898
rect 280794 310394 281414 311000
rect 280794 310158 280826 310394
rect 281062 310158 281146 310394
rect 281382 310158 281414 310394
rect 280794 310074 281414 310158
rect 280794 309838 280826 310074
rect 281062 309838 281146 310074
rect 281382 309838 281414 310074
rect 280794 308000 281414 309838
rect 289794 309454 290414 311000
rect 289794 309218 289826 309454
rect 290062 309218 290146 309454
rect 290382 309218 290414 309454
rect 289794 309134 290414 309218
rect 289794 308898 289826 309134
rect 290062 308898 290146 309134
rect 290382 308898 290414 309134
rect 289794 308000 290414 308898
rect 298794 310394 299414 311000
rect 298794 310158 298826 310394
rect 299062 310158 299146 310394
rect 299382 310158 299414 310394
rect 298794 310074 299414 310158
rect 298794 309838 298826 310074
rect 299062 309838 299146 310074
rect 299382 309838 299414 310074
rect 298794 308000 299414 309838
rect 307794 309454 308414 311000
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 308000 308414 308898
rect 316794 310394 317414 311000
rect 316794 310158 316826 310394
rect 317062 310158 317146 310394
rect 317382 310158 317414 310394
rect 316794 310074 317414 310158
rect 316794 309838 316826 310074
rect 317062 309838 317146 310074
rect 317382 309838 317414 310074
rect 316794 308000 317414 309838
rect 325794 309454 326414 311000
rect 325794 309218 325826 309454
rect 326062 309218 326146 309454
rect 326382 309218 326414 309454
rect 325794 309134 326414 309218
rect 325794 308898 325826 309134
rect 326062 308898 326146 309134
rect 326382 308898 326414 309134
rect 325794 308000 326414 308898
rect 334794 310394 335414 311000
rect 334794 310158 334826 310394
rect 335062 310158 335146 310394
rect 335382 310158 335414 310394
rect 334794 310074 335414 310158
rect 334794 309838 334826 310074
rect 335062 309838 335146 310074
rect 335382 309838 335414 310074
rect 334794 308000 335414 309838
rect 343794 309454 344414 311000
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 308000 344414 308898
rect 352794 310394 353414 311000
rect 352794 310158 352826 310394
rect 353062 310158 353146 310394
rect 353382 310158 353414 310394
rect 352794 310074 353414 310158
rect 352794 309838 352826 310074
rect 353062 309838 353146 310074
rect 353382 309838 353414 310074
rect 352794 308000 353414 309838
rect 361794 309454 362414 311000
rect 361794 309218 361826 309454
rect 362062 309218 362146 309454
rect 362382 309218 362414 309454
rect 361794 309134 362414 309218
rect 361794 308898 361826 309134
rect 362062 308898 362146 309134
rect 362382 308898 362414 309134
rect 361794 308000 362414 308898
rect 370794 310394 371414 311000
rect 370794 310158 370826 310394
rect 371062 310158 371146 310394
rect 371382 310158 371414 310394
rect 370794 310074 371414 310158
rect 370794 309838 370826 310074
rect 371062 309838 371146 310074
rect 371382 309838 371414 310074
rect 370794 308000 371414 309838
rect 379794 309454 380414 311000
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 308000 380414 308898
rect 388794 310394 389414 311000
rect 388794 310158 388826 310394
rect 389062 310158 389146 310394
rect 389382 310158 389414 310394
rect 388794 310074 389414 310158
rect 388794 309838 388826 310074
rect 389062 309838 389146 310074
rect 389382 309838 389414 310074
rect 388794 308000 389414 309838
rect 397794 309454 398414 311000
rect 397794 309218 397826 309454
rect 398062 309218 398146 309454
rect 398382 309218 398414 309454
rect 397794 309134 398414 309218
rect 397794 308898 397826 309134
rect 398062 308898 398146 309134
rect 398382 308898 398414 309134
rect 397794 308000 398414 308898
rect 406794 310394 407414 311000
rect 406794 310158 406826 310394
rect 407062 310158 407146 310394
rect 407382 310158 407414 310394
rect 406794 310074 407414 310158
rect 406794 309838 406826 310074
rect 407062 309838 407146 310074
rect 407382 309838 407414 310074
rect 406794 308000 407414 309838
rect 415794 309454 416414 311000
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 308000 416414 308898
rect 424794 310394 425414 311000
rect 424794 310158 424826 310394
rect 425062 310158 425146 310394
rect 425382 310158 425414 310394
rect 424794 310074 425414 310158
rect 424794 309838 424826 310074
rect 425062 309838 425146 310074
rect 425382 309838 425414 310074
rect 424794 308000 425414 309838
rect 433794 309454 434414 311000
rect 433794 309218 433826 309454
rect 434062 309218 434146 309454
rect 434382 309218 434414 309454
rect 433794 309134 434414 309218
rect 433794 308898 433826 309134
rect 434062 308898 434146 309134
rect 434382 308898 434414 309134
rect 433794 308000 434414 308898
rect 442794 310394 443414 311000
rect 442794 310158 442826 310394
rect 443062 310158 443146 310394
rect 443382 310158 443414 310394
rect 442794 310074 443414 310158
rect 442794 309838 442826 310074
rect 443062 309838 443146 310074
rect 443382 309838 443414 310074
rect 442794 308000 443414 309838
rect 451794 309454 452414 311000
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 308000 452414 308898
rect 460794 310394 461414 311000
rect 460794 310158 460826 310394
rect 461062 310158 461146 310394
rect 461382 310158 461414 310394
rect 460794 310074 461414 310158
rect 460794 309838 460826 310074
rect 461062 309838 461146 310074
rect 461382 309838 461414 310074
rect 460794 308000 461414 309838
rect 469794 309454 470414 311000
rect 469794 309218 469826 309454
rect 470062 309218 470146 309454
rect 470382 309218 470414 309454
rect 469794 309134 470414 309218
rect 469794 308898 469826 309134
rect 470062 308898 470146 309134
rect 470382 308898 470414 309134
rect 469794 308000 470414 308898
rect 478794 310394 479414 311000
rect 478794 310158 478826 310394
rect 479062 310158 479146 310394
rect 479382 310158 479414 310394
rect 478794 310074 479414 310158
rect 478794 309838 478826 310074
rect 479062 309838 479146 310074
rect 479382 309838 479414 310074
rect 478794 308000 479414 309838
rect 487794 309454 488414 311000
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 308000 488414 308898
rect 496794 310394 497414 311000
rect 496794 310158 496826 310394
rect 497062 310158 497146 310394
rect 497382 310158 497414 310394
rect 496794 310074 497414 310158
rect 496794 309838 496826 310074
rect 497062 309838 497146 310074
rect 497382 309838 497414 310074
rect 496794 308000 497414 309838
rect 505794 309454 506414 311000
rect 505794 309218 505826 309454
rect 506062 309218 506146 309454
rect 506382 309218 506414 309454
rect 505794 309134 506414 309218
rect 505794 308898 505826 309134
rect 506062 308898 506146 309134
rect 506382 308898 506414 309134
rect 505794 308000 506414 308898
rect 514794 310394 515414 311000
rect 514794 310158 514826 310394
rect 515062 310158 515146 310394
rect 515382 310158 515414 310394
rect 514794 310074 515414 310158
rect 514794 309838 514826 310074
rect 515062 309838 515146 310074
rect 515382 309838 515414 310074
rect 514794 308000 515414 309838
rect 523794 309454 524414 311000
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 308000 524414 308898
rect 532794 310394 533414 311000
rect 532794 310158 532826 310394
rect 533062 310158 533146 310394
rect 533382 310158 533414 310394
rect 532794 310074 533414 310158
rect 532794 309838 532826 310074
rect 533062 309838 533146 310074
rect 533382 309838 533414 310074
rect 532794 308000 533414 309838
rect 541794 309454 542414 311000
rect 541794 309218 541826 309454
rect 542062 309218 542146 309454
rect 542382 309218 542414 309454
rect 541794 309134 542414 309218
rect 541794 308898 541826 309134
rect 542062 308898 542146 309134
rect 542382 308898 542414 309134
rect 541794 308000 542414 308898
rect 550794 310394 551414 311000
rect 550794 310158 550826 310394
rect 551062 310158 551146 310394
rect 551382 310158 551414 310394
rect 550794 310074 551414 310158
rect 550794 309838 550826 310074
rect 551062 309838 551146 310074
rect 551382 309838 551414 310074
rect 550794 308000 551414 309838
rect 559794 309454 560414 326898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 282454 11414 299898
rect 22874 300454 23194 300486
rect 22874 300218 22916 300454
rect 23152 300218 23194 300454
rect 22874 300134 23194 300218
rect 22874 299898 22916 300134
rect 23152 299898 23194 300134
rect 22874 299866 23194 299898
rect 28805 300454 29125 300486
rect 28805 300218 28847 300454
rect 29083 300218 29125 300454
rect 28805 300134 29125 300218
rect 28805 299898 28847 300134
rect 29083 299898 29125 300134
rect 28805 299866 29125 299898
rect 49874 300454 50194 300486
rect 49874 300218 49916 300454
rect 50152 300218 50194 300454
rect 49874 300134 50194 300218
rect 49874 299898 49916 300134
rect 50152 299898 50194 300134
rect 49874 299866 50194 299898
rect 55805 300454 56125 300486
rect 55805 300218 55847 300454
rect 56083 300218 56125 300454
rect 55805 300134 56125 300218
rect 55805 299898 55847 300134
rect 56083 299898 56125 300134
rect 55805 299866 56125 299898
rect 76874 300454 77194 300486
rect 76874 300218 76916 300454
rect 77152 300218 77194 300454
rect 76874 300134 77194 300218
rect 76874 299898 76916 300134
rect 77152 299898 77194 300134
rect 76874 299866 77194 299898
rect 82805 300454 83125 300486
rect 82805 300218 82847 300454
rect 83083 300218 83125 300454
rect 82805 300134 83125 300218
rect 82805 299898 82847 300134
rect 83083 299898 83125 300134
rect 82805 299866 83125 299898
rect 103874 300454 104194 300486
rect 103874 300218 103916 300454
rect 104152 300218 104194 300454
rect 103874 300134 104194 300218
rect 103874 299898 103916 300134
rect 104152 299898 104194 300134
rect 103874 299866 104194 299898
rect 109805 300454 110125 300486
rect 109805 300218 109847 300454
rect 110083 300218 110125 300454
rect 109805 300134 110125 300218
rect 109805 299898 109847 300134
rect 110083 299898 110125 300134
rect 109805 299866 110125 299898
rect 130874 300454 131194 300486
rect 130874 300218 130916 300454
rect 131152 300218 131194 300454
rect 130874 300134 131194 300218
rect 130874 299898 130916 300134
rect 131152 299898 131194 300134
rect 130874 299866 131194 299898
rect 136805 300454 137125 300486
rect 136805 300218 136847 300454
rect 137083 300218 137125 300454
rect 136805 300134 137125 300218
rect 136805 299898 136847 300134
rect 137083 299898 137125 300134
rect 136805 299866 137125 299898
rect 157874 300454 158194 300486
rect 157874 300218 157916 300454
rect 158152 300218 158194 300454
rect 157874 300134 158194 300218
rect 157874 299898 157916 300134
rect 158152 299898 158194 300134
rect 157874 299866 158194 299898
rect 163805 300454 164125 300486
rect 163805 300218 163847 300454
rect 164083 300218 164125 300454
rect 163805 300134 164125 300218
rect 163805 299898 163847 300134
rect 164083 299898 164125 300134
rect 163805 299866 164125 299898
rect 184874 300454 185194 300486
rect 184874 300218 184916 300454
rect 185152 300218 185194 300454
rect 184874 300134 185194 300218
rect 184874 299898 184916 300134
rect 185152 299898 185194 300134
rect 184874 299866 185194 299898
rect 190805 300454 191125 300486
rect 190805 300218 190847 300454
rect 191083 300218 191125 300454
rect 190805 300134 191125 300218
rect 190805 299898 190847 300134
rect 191083 299898 191125 300134
rect 190805 299866 191125 299898
rect 211874 300454 212194 300486
rect 211874 300218 211916 300454
rect 212152 300218 212194 300454
rect 211874 300134 212194 300218
rect 211874 299898 211916 300134
rect 212152 299898 212194 300134
rect 211874 299866 212194 299898
rect 217805 300454 218125 300486
rect 217805 300218 217847 300454
rect 218083 300218 218125 300454
rect 217805 300134 218125 300218
rect 217805 299898 217847 300134
rect 218083 299898 218125 300134
rect 217805 299866 218125 299898
rect 238874 300454 239194 300486
rect 238874 300218 238916 300454
rect 239152 300218 239194 300454
rect 238874 300134 239194 300218
rect 238874 299898 238916 300134
rect 239152 299898 239194 300134
rect 238874 299866 239194 299898
rect 244805 300454 245125 300486
rect 244805 300218 244847 300454
rect 245083 300218 245125 300454
rect 244805 300134 245125 300218
rect 244805 299898 244847 300134
rect 245083 299898 245125 300134
rect 244805 299866 245125 299898
rect 265874 300454 266194 300486
rect 265874 300218 265916 300454
rect 266152 300218 266194 300454
rect 265874 300134 266194 300218
rect 265874 299898 265916 300134
rect 266152 299898 266194 300134
rect 265874 299866 266194 299898
rect 271805 300454 272125 300486
rect 271805 300218 271847 300454
rect 272083 300218 272125 300454
rect 271805 300134 272125 300218
rect 271805 299898 271847 300134
rect 272083 299898 272125 300134
rect 271805 299866 272125 299898
rect 292874 300454 293194 300486
rect 292874 300218 292916 300454
rect 293152 300218 293194 300454
rect 292874 300134 293194 300218
rect 292874 299898 292916 300134
rect 293152 299898 293194 300134
rect 292874 299866 293194 299898
rect 298805 300454 299125 300486
rect 298805 300218 298847 300454
rect 299083 300218 299125 300454
rect 298805 300134 299125 300218
rect 298805 299898 298847 300134
rect 299083 299898 299125 300134
rect 298805 299866 299125 299898
rect 319874 300454 320194 300486
rect 319874 300218 319916 300454
rect 320152 300218 320194 300454
rect 319874 300134 320194 300218
rect 319874 299898 319916 300134
rect 320152 299898 320194 300134
rect 319874 299866 320194 299898
rect 325805 300454 326125 300486
rect 325805 300218 325847 300454
rect 326083 300218 326125 300454
rect 325805 300134 326125 300218
rect 325805 299898 325847 300134
rect 326083 299898 326125 300134
rect 325805 299866 326125 299898
rect 346874 300454 347194 300486
rect 346874 300218 346916 300454
rect 347152 300218 347194 300454
rect 346874 300134 347194 300218
rect 346874 299898 346916 300134
rect 347152 299898 347194 300134
rect 346874 299866 347194 299898
rect 352805 300454 353125 300486
rect 352805 300218 352847 300454
rect 353083 300218 353125 300454
rect 352805 300134 353125 300218
rect 352805 299898 352847 300134
rect 353083 299898 353125 300134
rect 352805 299866 353125 299898
rect 373874 300454 374194 300486
rect 373874 300218 373916 300454
rect 374152 300218 374194 300454
rect 373874 300134 374194 300218
rect 373874 299898 373916 300134
rect 374152 299898 374194 300134
rect 373874 299866 374194 299898
rect 379805 300454 380125 300486
rect 379805 300218 379847 300454
rect 380083 300218 380125 300454
rect 379805 300134 380125 300218
rect 379805 299898 379847 300134
rect 380083 299898 380125 300134
rect 379805 299866 380125 299898
rect 400874 300454 401194 300486
rect 400874 300218 400916 300454
rect 401152 300218 401194 300454
rect 400874 300134 401194 300218
rect 400874 299898 400916 300134
rect 401152 299898 401194 300134
rect 400874 299866 401194 299898
rect 406805 300454 407125 300486
rect 406805 300218 406847 300454
rect 407083 300218 407125 300454
rect 406805 300134 407125 300218
rect 406805 299898 406847 300134
rect 407083 299898 407125 300134
rect 406805 299866 407125 299898
rect 427874 300454 428194 300486
rect 427874 300218 427916 300454
rect 428152 300218 428194 300454
rect 427874 300134 428194 300218
rect 427874 299898 427916 300134
rect 428152 299898 428194 300134
rect 427874 299866 428194 299898
rect 433805 300454 434125 300486
rect 433805 300218 433847 300454
rect 434083 300218 434125 300454
rect 433805 300134 434125 300218
rect 433805 299898 433847 300134
rect 434083 299898 434125 300134
rect 433805 299866 434125 299898
rect 454874 300454 455194 300486
rect 454874 300218 454916 300454
rect 455152 300218 455194 300454
rect 454874 300134 455194 300218
rect 454874 299898 454916 300134
rect 455152 299898 455194 300134
rect 454874 299866 455194 299898
rect 460805 300454 461125 300486
rect 460805 300218 460847 300454
rect 461083 300218 461125 300454
rect 460805 300134 461125 300218
rect 460805 299898 460847 300134
rect 461083 299898 461125 300134
rect 460805 299866 461125 299898
rect 481874 300454 482194 300486
rect 481874 300218 481916 300454
rect 482152 300218 482194 300454
rect 481874 300134 482194 300218
rect 481874 299898 481916 300134
rect 482152 299898 482194 300134
rect 481874 299866 482194 299898
rect 487805 300454 488125 300486
rect 487805 300218 487847 300454
rect 488083 300218 488125 300454
rect 487805 300134 488125 300218
rect 487805 299898 487847 300134
rect 488083 299898 488125 300134
rect 487805 299866 488125 299898
rect 508874 300454 509194 300486
rect 508874 300218 508916 300454
rect 509152 300218 509194 300454
rect 508874 300134 509194 300218
rect 508874 299898 508916 300134
rect 509152 299898 509194 300134
rect 508874 299866 509194 299898
rect 514805 300454 515125 300486
rect 514805 300218 514847 300454
rect 515083 300218 515125 300454
rect 514805 300134 515125 300218
rect 514805 299898 514847 300134
rect 515083 299898 515125 300134
rect 514805 299866 515125 299898
rect 535874 300454 536194 300486
rect 535874 300218 535916 300454
rect 536152 300218 536194 300454
rect 535874 300134 536194 300218
rect 535874 299898 535916 300134
rect 536152 299898 536194 300134
rect 535874 299866 536194 299898
rect 541805 300454 542125 300486
rect 541805 300218 541847 300454
rect 542083 300218 542125 300454
rect 541805 300134 542125 300218
rect 541805 299898 541847 300134
rect 542083 299898 542125 300134
rect 541805 299866 542125 299898
rect 19910 291454 20230 291486
rect 19910 291218 19952 291454
rect 20188 291218 20230 291454
rect 19910 291134 20230 291218
rect 19910 290898 19952 291134
rect 20188 290898 20230 291134
rect 19910 290866 20230 290898
rect 25840 291454 26160 291486
rect 25840 291218 25882 291454
rect 26118 291218 26160 291454
rect 25840 291134 26160 291218
rect 25840 290898 25882 291134
rect 26118 290898 26160 291134
rect 25840 290866 26160 290898
rect 31771 291454 32091 291486
rect 31771 291218 31813 291454
rect 32049 291218 32091 291454
rect 31771 291134 32091 291218
rect 31771 290898 31813 291134
rect 32049 290898 32091 291134
rect 31771 290866 32091 290898
rect 46910 291454 47230 291486
rect 46910 291218 46952 291454
rect 47188 291218 47230 291454
rect 46910 291134 47230 291218
rect 46910 290898 46952 291134
rect 47188 290898 47230 291134
rect 46910 290866 47230 290898
rect 52840 291454 53160 291486
rect 52840 291218 52882 291454
rect 53118 291218 53160 291454
rect 52840 291134 53160 291218
rect 52840 290898 52882 291134
rect 53118 290898 53160 291134
rect 52840 290866 53160 290898
rect 58771 291454 59091 291486
rect 58771 291218 58813 291454
rect 59049 291218 59091 291454
rect 58771 291134 59091 291218
rect 58771 290898 58813 291134
rect 59049 290898 59091 291134
rect 58771 290866 59091 290898
rect 73910 291454 74230 291486
rect 73910 291218 73952 291454
rect 74188 291218 74230 291454
rect 73910 291134 74230 291218
rect 73910 290898 73952 291134
rect 74188 290898 74230 291134
rect 73910 290866 74230 290898
rect 79840 291454 80160 291486
rect 79840 291218 79882 291454
rect 80118 291218 80160 291454
rect 79840 291134 80160 291218
rect 79840 290898 79882 291134
rect 80118 290898 80160 291134
rect 79840 290866 80160 290898
rect 85771 291454 86091 291486
rect 85771 291218 85813 291454
rect 86049 291218 86091 291454
rect 85771 291134 86091 291218
rect 85771 290898 85813 291134
rect 86049 290898 86091 291134
rect 85771 290866 86091 290898
rect 100910 291454 101230 291486
rect 100910 291218 100952 291454
rect 101188 291218 101230 291454
rect 100910 291134 101230 291218
rect 100910 290898 100952 291134
rect 101188 290898 101230 291134
rect 100910 290866 101230 290898
rect 106840 291454 107160 291486
rect 106840 291218 106882 291454
rect 107118 291218 107160 291454
rect 106840 291134 107160 291218
rect 106840 290898 106882 291134
rect 107118 290898 107160 291134
rect 106840 290866 107160 290898
rect 112771 291454 113091 291486
rect 112771 291218 112813 291454
rect 113049 291218 113091 291454
rect 112771 291134 113091 291218
rect 112771 290898 112813 291134
rect 113049 290898 113091 291134
rect 112771 290866 113091 290898
rect 127910 291454 128230 291486
rect 127910 291218 127952 291454
rect 128188 291218 128230 291454
rect 127910 291134 128230 291218
rect 127910 290898 127952 291134
rect 128188 290898 128230 291134
rect 127910 290866 128230 290898
rect 133840 291454 134160 291486
rect 133840 291218 133882 291454
rect 134118 291218 134160 291454
rect 133840 291134 134160 291218
rect 133840 290898 133882 291134
rect 134118 290898 134160 291134
rect 133840 290866 134160 290898
rect 139771 291454 140091 291486
rect 139771 291218 139813 291454
rect 140049 291218 140091 291454
rect 139771 291134 140091 291218
rect 139771 290898 139813 291134
rect 140049 290898 140091 291134
rect 139771 290866 140091 290898
rect 154910 291454 155230 291486
rect 154910 291218 154952 291454
rect 155188 291218 155230 291454
rect 154910 291134 155230 291218
rect 154910 290898 154952 291134
rect 155188 290898 155230 291134
rect 154910 290866 155230 290898
rect 160840 291454 161160 291486
rect 160840 291218 160882 291454
rect 161118 291218 161160 291454
rect 160840 291134 161160 291218
rect 160840 290898 160882 291134
rect 161118 290898 161160 291134
rect 160840 290866 161160 290898
rect 166771 291454 167091 291486
rect 166771 291218 166813 291454
rect 167049 291218 167091 291454
rect 166771 291134 167091 291218
rect 166771 290898 166813 291134
rect 167049 290898 167091 291134
rect 166771 290866 167091 290898
rect 181910 291454 182230 291486
rect 181910 291218 181952 291454
rect 182188 291218 182230 291454
rect 181910 291134 182230 291218
rect 181910 290898 181952 291134
rect 182188 290898 182230 291134
rect 181910 290866 182230 290898
rect 187840 291454 188160 291486
rect 187840 291218 187882 291454
rect 188118 291218 188160 291454
rect 187840 291134 188160 291218
rect 187840 290898 187882 291134
rect 188118 290898 188160 291134
rect 187840 290866 188160 290898
rect 193771 291454 194091 291486
rect 193771 291218 193813 291454
rect 194049 291218 194091 291454
rect 193771 291134 194091 291218
rect 193771 290898 193813 291134
rect 194049 290898 194091 291134
rect 193771 290866 194091 290898
rect 208910 291454 209230 291486
rect 208910 291218 208952 291454
rect 209188 291218 209230 291454
rect 208910 291134 209230 291218
rect 208910 290898 208952 291134
rect 209188 290898 209230 291134
rect 208910 290866 209230 290898
rect 214840 291454 215160 291486
rect 214840 291218 214882 291454
rect 215118 291218 215160 291454
rect 214840 291134 215160 291218
rect 214840 290898 214882 291134
rect 215118 290898 215160 291134
rect 214840 290866 215160 290898
rect 220771 291454 221091 291486
rect 220771 291218 220813 291454
rect 221049 291218 221091 291454
rect 220771 291134 221091 291218
rect 220771 290898 220813 291134
rect 221049 290898 221091 291134
rect 220771 290866 221091 290898
rect 235910 291454 236230 291486
rect 235910 291218 235952 291454
rect 236188 291218 236230 291454
rect 235910 291134 236230 291218
rect 235910 290898 235952 291134
rect 236188 290898 236230 291134
rect 235910 290866 236230 290898
rect 241840 291454 242160 291486
rect 241840 291218 241882 291454
rect 242118 291218 242160 291454
rect 241840 291134 242160 291218
rect 241840 290898 241882 291134
rect 242118 290898 242160 291134
rect 241840 290866 242160 290898
rect 247771 291454 248091 291486
rect 247771 291218 247813 291454
rect 248049 291218 248091 291454
rect 247771 291134 248091 291218
rect 247771 290898 247813 291134
rect 248049 290898 248091 291134
rect 247771 290866 248091 290898
rect 262910 291454 263230 291486
rect 262910 291218 262952 291454
rect 263188 291218 263230 291454
rect 262910 291134 263230 291218
rect 262910 290898 262952 291134
rect 263188 290898 263230 291134
rect 262910 290866 263230 290898
rect 268840 291454 269160 291486
rect 268840 291218 268882 291454
rect 269118 291218 269160 291454
rect 268840 291134 269160 291218
rect 268840 290898 268882 291134
rect 269118 290898 269160 291134
rect 268840 290866 269160 290898
rect 274771 291454 275091 291486
rect 274771 291218 274813 291454
rect 275049 291218 275091 291454
rect 274771 291134 275091 291218
rect 274771 290898 274813 291134
rect 275049 290898 275091 291134
rect 274771 290866 275091 290898
rect 289910 291454 290230 291486
rect 289910 291218 289952 291454
rect 290188 291218 290230 291454
rect 289910 291134 290230 291218
rect 289910 290898 289952 291134
rect 290188 290898 290230 291134
rect 289910 290866 290230 290898
rect 295840 291454 296160 291486
rect 295840 291218 295882 291454
rect 296118 291218 296160 291454
rect 295840 291134 296160 291218
rect 295840 290898 295882 291134
rect 296118 290898 296160 291134
rect 295840 290866 296160 290898
rect 301771 291454 302091 291486
rect 301771 291218 301813 291454
rect 302049 291218 302091 291454
rect 301771 291134 302091 291218
rect 301771 290898 301813 291134
rect 302049 290898 302091 291134
rect 301771 290866 302091 290898
rect 316910 291454 317230 291486
rect 316910 291218 316952 291454
rect 317188 291218 317230 291454
rect 316910 291134 317230 291218
rect 316910 290898 316952 291134
rect 317188 290898 317230 291134
rect 316910 290866 317230 290898
rect 322840 291454 323160 291486
rect 322840 291218 322882 291454
rect 323118 291218 323160 291454
rect 322840 291134 323160 291218
rect 322840 290898 322882 291134
rect 323118 290898 323160 291134
rect 322840 290866 323160 290898
rect 328771 291454 329091 291486
rect 328771 291218 328813 291454
rect 329049 291218 329091 291454
rect 328771 291134 329091 291218
rect 328771 290898 328813 291134
rect 329049 290898 329091 291134
rect 328771 290866 329091 290898
rect 343910 291454 344230 291486
rect 343910 291218 343952 291454
rect 344188 291218 344230 291454
rect 343910 291134 344230 291218
rect 343910 290898 343952 291134
rect 344188 290898 344230 291134
rect 343910 290866 344230 290898
rect 349840 291454 350160 291486
rect 349840 291218 349882 291454
rect 350118 291218 350160 291454
rect 349840 291134 350160 291218
rect 349840 290898 349882 291134
rect 350118 290898 350160 291134
rect 349840 290866 350160 290898
rect 355771 291454 356091 291486
rect 355771 291218 355813 291454
rect 356049 291218 356091 291454
rect 355771 291134 356091 291218
rect 355771 290898 355813 291134
rect 356049 290898 356091 291134
rect 355771 290866 356091 290898
rect 370910 291454 371230 291486
rect 370910 291218 370952 291454
rect 371188 291218 371230 291454
rect 370910 291134 371230 291218
rect 370910 290898 370952 291134
rect 371188 290898 371230 291134
rect 370910 290866 371230 290898
rect 376840 291454 377160 291486
rect 376840 291218 376882 291454
rect 377118 291218 377160 291454
rect 376840 291134 377160 291218
rect 376840 290898 376882 291134
rect 377118 290898 377160 291134
rect 376840 290866 377160 290898
rect 382771 291454 383091 291486
rect 382771 291218 382813 291454
rect 383049 291218 383091 291454
rect 382771 291134 383091 291218
rect 382771 290898 382813 291134
rect 383049 290898 383091 291134
rect 382771 290866 383091 290898
rect 397910 291454 398230 291486
rect 397910 291218 397952 291454
rect 398188 291218 398230 291454
rect 397910 291134 398230 291218
rect 397910 290898 397952 291134
rect 398188 290898 398230 291134
rect 397910 290866 398230 290898
rect 403840 291454 404160 291486
rect 403840 291218 403882 291454
rect 404118 291218 404160 291454
rect 403840 291134 404160 291218
rect 403840 290898 403882 291134
rect 404118 290898 404160 291134
rect 403840 290866 404160 290898
rect 409771 291454 410091 291486
rect 409771 291218 409813 291454
rect 410049 291218 410091 291454
rect 409771 291134 410091 291218
rect 409771 290898 409813 291134
rect 410049 290898 410091 291134
rect 409771 290866 410091 290898
rect 424910 291454 425230 291486
rect 424910 291218 424952 291454
rect 425188 291218 425230 291454
rect 424910 291134 425230 291218
rect 424910 290898 424952 291134
rect 425188 290898 425230 291134
rect 424910 290866 425230 290898
rect 430840 291454 431160 291486
rect 430840 291218 430882 291454
rect 431118 291218 431160 291454
rect 430840 291134 431160 291218
rect 430840 290898 430882 291134
rect 431118 290898 431160 291134
rect 430840 290866 431160 290898
rect 436771 291454 437091 291486
rect 436771 291218 436813 291454
rect 437049 291218 437091 291454
rect 436771 291134 437091 291218
rect 436771 290898 436813 291134
rect 437049 290898 437091 291134
rect 436771 290866 437091 290898
rect 451910 291454 452230 291486
rect 451910 291218 451952 291454
rect 452188 291218 452230 291454
rect 451910 291134 452230 291218
rect 451910 290898 451952 291134
rect 452188 290898 452230 291134
rect 451910 290866 452230 290898
rect 457840 291454 458160 291486
rect 457840 291218 457882 291454
rect 458118 291218 458160 291454
rect 457840 291134 458160 291218
rect 457840 290898 457882 291134
rect 458118 290898 458160 291134
rect 457840 290866 458160 290898
rect 463771 291454 464091 291486
rect 463771 291218 463813 291454
rect 464049 291218 464091 291454
rect 463771 291134 464091 291218
rect 463771 290898 463813 291134
rect 464049 290898 464091 291134
rect 463771 290866 464091 290898
rect 478910 291454 479230 291486
rect 478910 291218 478952 291454
rect 479188 291218 479230 291454
rect 478910 291134 479230 291218
rect 478910 290898 478952 291134
rect 479188 290898 479230 291134
rect 478910 290866 479230 290898
rect 484840 291454 485160 291486
rect 484840 291218 484882 291454
rect 485118 291218 485160 291454
rect 484840 291134 485160 291218
rect 484840 290898 484882 291134
rect 485118 290898 485160 291134
rect 484840 290866 485160 290898
rect 490771 291454 491091 291486
rect 490771 291218 490813 291454
rect 491049 291218 491091 291454
rect 490771 291134 491091 291218
rect 490771 290898 490813 291134
rect 491049 290898 491091 291134
rect 490771 290866 491091 290898
rect 505910 291454 506230 291486
rect 505910 291218 505952 291454
rect 506188 291218 506230 291454
rect 505910 291134 506230 291218
rect 505910 290898 505952 291134
rect 506188 290898 506230 291134
rect 505910 290866 506230 290898
rect 511840 291454 512160 291486
rect 511840 291218 511882 291454
rect 512118 291218 512160 291454
rect 511840 291134 512160 291218
rect 511840 290898 511882 291134
rect 512118 290898 512160 291134
rect 511840 290866 512160 290898
rect 517771 291454 518091 291486
rect 517771 291218 517813 291454
rect 518049 291218 518091 291454
rect 517771 291134 518091 291218
rect 517771 290898 517813 291134
rect 518049 290898 518091 291134
rect 517771 290866 518091 290898
rect 532910 291454 533230 291486
rect 532910 291218 532952 291454
rect 533188 291218 533230 291454
rect 532910 291134 533230 291218
rect 532910 290898 532952 291134
rect 533188 290898 533230 291134
rect 532910 290866 533230 290898
rect 538840 291454 539160 291486
rect 538840 291218 538882 291454
rect 539118 291218 539160 291454
rect 538840 291134 539160 291218
rect 538840 290898 538882 291134
rect 539118 290898 539160 291134
rect 538840 290866 539160 290898
rect 544771 291454 545091 291486
rect 544771 291218 544813 291454
rect 545049 291218 545091 291454
rect 544771 291134 545091 291218
rect 544771 290898 544813 291134
rect 545049 290898 545091 291134
rect 544771 290866 545091 290898
rect 559794 291454 560414 308898
rect 559794 291218 559826 291454
rect 560062 291218 560146 291454
rect 560382 291218 560414 291454
rect 559794 291134 560414 291218
rect 559794 290898 559826 291134
rect 560062 290898 560146 291134
rect 560382 290898 560414 291134
rect 10794 282218 10826 282454
rect 11062 282218 11146 282454
rect 11382 282218 11414 282454
rect 10794 282134 11414 282218
rect 10794 281898 10826 282134
rect 11062 281898 11146 282134
rect 11382 281898 11414 282134
rect 10794 264454 11414 281898
rect 19794 283394 20414 284000
rect 19794 283158 19826 283394
rect 20062 283158 20146 283394
rect 20382 283158 20414 283394
rect 19794 283074 20414 283158
rect 19794 282838 19826 283074
rect 20062 282838 20146 283074
rect 20382 282838 20414 283074
rect 19794 281000 20414 282838
rect 28794 282454 29414 284000
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 281000 29414 281898
rect 37794 283394 38414 284000
rect 37794 283158 37826 283394
rect 38062 283158 38146 283394
rect 38382 283158 38414 283394
rect 37794 283074 38414 283158
rect 37794 282838 37826 283074
rect 38062 282838 38146 283074
rect 38382 282838 38414 283074
rect 37794 281000 38414 282838
rect 46794 282454 47414 284000
rect 46794 282218 46826 282454
rect 47062 282218 47146 282454
rect 47382 282218 47414 282454
rect 46794 282134 47414 282218
rect 46794 281898 46826 282134
rect 47062 281898 47146 282134
rect 47382 281898 47414 282134
rect 46794 281000 47414 281898
rect 55794 283394 56414 284000
rect 55794 283158 55826 283394
rect 56062 283158 56146 283394
rect 56382 283158 56414 283394
rect 55794 283074 56414 283158
rect 55794 282838 55826 283074
rect 56062 282838 56146 283074
rect 56382 282838 56414 283074
rect 55794 281000 56414 282838
rect 64794 282454 65414 284000
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 281000 65414 281898
rect 73794 283394 74414 284000
rect 73794 283158 73826 283394
rect 74062 283158 74146 283394
rect 74382 283158 74414 283394
rect 73794 283074 74414 283158
rect 73794 282838 73826 283074
rect 74062 282838 74146 283074
rect 74382 282838 74414 283074
rect 73794 281000 74414 282838
rect 82794 282454 83414 284000
rect 82794 282218 82826 282454
rect 83062 282218 83146 282454
rect 83382 282218 83414 282454
rect 82794 282134 83414 282218
rect 82794 281898 82826 282134
rect 83062 281898 83146 282134
rect 83382 281898 83414 282134
rect 82794 281000 83414 281898
rect 91794 283394 92414 284000
rect 91794 283158 91826 283394
rect 92062 283158 92146 283394
rect 92382 283158 92414 283394
rect 91794 283074 92414 283158
rect 91794 282838 91826 283074
rect 92062 282838 92146 283074
rect 92382 282838 92414 283074
rect 91794 281000 92414 282838
rect 100794 282454 101414 284000
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 281000 101414 281898
rect 109794 283394 110414 284000
rect 109794 283158 109826 283394
rect 110062 283158 110146 283394
rect 110382 283158 110414 283394
rect 109794 283074 110414 283158
rect 109794 282838 109826 283074
rect 110062 282838 110146 283074
rect 110382 282838 110414 283074
rect 109794 281000 110414 282838
rect 118794 282454 119414 284000
rect 118794 282218 118826 282454
rect 119062 282218 119146 282454
rect 119382 282218 119414 282454
rect 118794 282134 119414 282218
rect 118794 281898 118826 282134
rect 119062 281898 119146 282134
rect 119382 281898 119414 282134
rect 118794 281000 119414 281898
rect 127794 283394 128414 284000
rect 127794 283158 127826 283394
rect 128062 283158 128146 283394
rect 128382 283158 128414 283394
rect 127794 283074 128414 283158
rect 127794 282838 127826 283074
rect 128062 282838 128146 283074
rect 128382 282838 128414 283074
rect 127794 281000 128414 282838
rect 136794 282454 137414 284000
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 281000 137414 281898
rect 145794 283394 146414 284000
rect 145794 283158 145826 283394
rect 146062 283158 146146 283394
rect 146382 283158 146414 283394
rect 145794 283074 146414 283158
rect 145794 282838 145826 283074
rect 146062 282838 146146 283074
rect 146382 282838 146414 283074
rect 145794 281000 146414 282838
rect 154794 282454 155414 284000
rect 154794 282218 154826 282454
rect 155062 282218 155146 282454
rect 155382 282218 155414 282454
rect 154794 282134 155414 282218
rect 154794 281898 154826 282134
rect 155062 281898 155146 282134
rect 155382 281898 155414 282134
rect 154794 281000 155414 281898
rect 163794 283394 164414 284000
rect 163794 283158 163826 283394
rect 164062 283158 164146 283394
rect 164382 283158 164414 283394
rect 163794 283074 164414 283158
rect 163794 282838 163826 283074
rect 164062 282838 164146 283074
rect 164382 282838 164414 283074
rect 163794 281000 164414 282838
rect 172794 282454 173414 284000
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 281000 173414 281898
rect 181794 283394 182414 284000
rect 181794 283158 181826 283394
rect 182062 283158 182146 283394
rect 182382 283158 182414 283394
rect 181794 283074 182414 283158
rect 181794 282838 181826 283074
rect 182062 282838 182146 283074
rect 182382 282838 182414 283074
rect 181794 281000 182414 282838
rect 190794 282454 191414 284000
rect 190794 282218 190826 282454
rect 191062 282218 191146 282454
rect 191382 282218 191414 282454
rect 190794 282134 191414 282218
rect 190794 281898 190826 282134
rect 191062 281898 191146 282134
rect 191382 281898 191414 282134
rect 190794 281000 191414 281898
rect 199794 283394 200414 284000
rect 199794 283158 199826 283394
rect 200062 283158 200146 283394
rect 200382 283158 200414 283394
rect 199794 283074 200414 283158
rect 199794 282838 199826 283074
rect 200062 282838 200146 283074
rect 200382 282838 200414 283074
rect 199794 281000 200414 282838
rect 208794 282454 209414 284000
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 281000 209414 281898
rect 217794 283394 218414 284000
rect 217794 283158 217826 283394
rect 218062 283158 218146 283394
rect 218382 283158 218414 283394
rect 217794 283074 218414 283158
rect 217794 282838 217826 283074
rect 218062 282838 218146 283074
rect 218382 282838 218414 283074
rect 217794 281000 218414 282838
rect 226794 282454 227414 284000
rect 226794 282218 226826 282454
rect 227062 282218 227146 282454
rect 227382 282218 227414 282454
rect 226794 282134 227414 282218
rect 226794 281898 226826 282134
rect 227062 281898 227146 282134
rect 227382 281898 227414 282134
rect 226794 281000 227414 281898
rect 235794 283394 236414 284000
rect 235794 283158 235826 283394
rect 236062 283158 236146 283394
rect 236382 283158 236414 283394
rect 235794 283074 236414 283158
rect 235794 282838 235826 283074
rect 236062 282838 236146 283074
rect 236382 282838 236414 283074
rect 235794 281000 236414 282838
rect 244794 282454 245414 284000
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 281000 245414 281898
rect 253794 283394 254414 284000
rect 253794 283158 253826 283394
rect 254062 283158 254146 283394
rect 254382 283158 254414 283394
rect 253794 283074 254414 283158
rect 253794 282838 253826 283074
rect 254062 282838 254146 283074
rect 254382 282838 254414 283074
rect 253794 281000 254414 282838
rect 262794 282454 263414 284000
rect 262794 282218 262826 282454
rect 263062 282218 263146 282454
rect 263382 282218 263414 282454
rect 262794 282134 263414 282218
rect 262794 281898 262826 282134
rect 263062 281898 263146 282134
rect 263382 281898 263414 282134
rect 262794 281000 263414 281898
rect 271794 283394 272414 284000
rect 271794 283158 271826 283394
rect 272062 283158 272146 283394
rect 272382 283158 272414 283394
rect 271794 283074 272414 283158
rect 271794 282838 271826 283074
rect 272062 282838 272146 283074
rect 272382 282838 272414 283074
rect 271794 281000 272414 282838
rect 280794 282454 281414 284000
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 281000 281414 281898
rect 289794 283394 290414 284000
rect 289794 283158 289826 283394
rect 290062 283158 290146 283394
rect 290382 283158 290414 283394
rect 289794 283074 290414 283158
rect 289794 282838 289826 283074
rect 290062 282838 290146 283074
rect 290382 282838 290414 283074
rect 289794 281000 290414 282838
rect 298794 282454 299414 284000
rect 298794 282218 298826 282454
rect 299062 282218 299146 282454
rect 299382 282218 299414 282454
rect 298794 282134 299414 282218
rect 298794 281898 298826 282134
rect 299062 281898 299146 282134
rect 299382 281898 299414 282134
rect 298794 281000 299414 281898
rect 307794 283394 308414 284000
rect 307794 283158 307826 283394
rect 308062 283158 308146 283394
rect 308382 283158 308414 283394
rect 307794 283074 308414 283158
rect 307794 282838 307826 283074
rect 308062 282838 308146 283074
rect 308382 282838 308414 283074
rect 307794 281000 308414 282838
rect 316794 282454 317414 284000
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 281000 317414 281898
rect 325794 283394 326414 284000
rect 325794 283158 325826 283394
rect 326062 283158 326146 283394
rect 326382 283158 326414 283394
rect 325794 283074 326414 283158
rect 325794 282838 325826 283074
rect 326062 282838 326146 283074
rect 326382 282838 326414 283074
rect 325794 281000 326414 282838
rect 334794 282454 335414 284000
rect 334794 282218 334826 282454
rect 335062 282218 335146 282454
rect 335382 282218 335414 282454
rect 334794 282134 335414 282218
rect 334794 281898 334826 282134
rect 335062 281898 335146 282134
rect 335382 281898 335414 282134
rect 334794 281000 335414 281898
rect 343794 283394 344414 284000
rect 343794 283158 343826 283394
rect 344062 283158 344146 283394
rect 344382 283158 344414 283394
rect 343794 283074 344414 283158
rect 343794 282838 343826 283074
rect 344062 282838 344146 283074
rect 344382 282838 344414 283074
rect 343794 281000 344414 282838
rect 352794 282454 353414 284000
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 281000 353414 281898
rect 361794 283394 362414 284000
rect 361794 283158 361826 283394
rect 362062 283158 362146 283394
rect 362382 283158 362414 283394
rect 361794 283074 362414 283158
rect 361794 282838 361826 283074
rect 362062 282838 362146 283074
rect 362382 282838 362414 283074
rect 361794 281000 362414 282838
rect 370794 282454 371414 284000
rect 370794 282218 370826 282454
rect 371062 282218 371146 282454
rect 371382 282218 371414 282454
rect 370794 282134 371414 282218
rect 370794 281898 370826 282134
rect 371062 281898 371146 282134
rect 371382 281898 371414 282134
rect 370794 281000 371414 281898
rect 379794 283394 380414 284000
rect 379794 283158 379826 283394
rect 380062 283158 380146 283394
rect 380382 283158 380414 283394
rect 379794 283074 380414 283158
rect 379794 282838 379826 283074
rect 380062 282838 380146 283074
rect 380382 282838 380414 283074
rect 379794 281000 380414 282838
rect 388794 282454 389414 284000
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 281000 389414 281898
rect 397794 283394 398414 284000
rect 397794 283158 397826 283394
rect 398062 283158 398146 283394
rect 398382 283158 398414 283394
rect 397794 283074 398414 283158
rect 397794 282838 397826 283074
rect 398062 282838 398146 283074
rect 398382 282838 398414 283074
rect 397794 281000 398414 282838
rect 406794 282454 407414 284000
rect 406794 282218 406826 282454
rect 407062 282218 407146 282454
rect 407382 282218 407414 282454
rect 406794 282134 407414 282218
rect 406794 281898 406826 282134
rect 407062 281898 407146 282134
rect 407382 281898 407414 282134
rect 406794 281000 407414 281898
rect 415794 283394 416414 284000
rect 415794 283158 415826 283394
rect 416062 283158 416146 283394
rect 416382 283158 416414 283394
rect 415794 283074 416414 283158
rect 415794 282838 415826 283074
rect 416062 282838 416146 283074
rect 416382 282838 416414 283074
rect 415794 281000 416414 282838
rect 424794 282454 425414 284000
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 281000 425414 281898
rect 433794 283394 434414 284000
rect 433794 283158 433826 283394
rect 434062 283158 434146 283394
rect 434382 283158 434414 283394
rect 433794 283074 434414 283158
rect 433794 282838 433826 283074
rect 434062 282838 434146 283074
rect 434382 282838 434414 283074
rect 433794 281000 434414 282838
rect 442794 282454 443414 284000
rect 442794 282218 442826 282454
rect 443062 282218 443146 282454
rect 443382 282218 443414 282454
rect 442794 282134 443414 282218
rect 442794 281898 442826 282134
rect 443062 281898 443146 282134
rect 443382 281898 443414 282134
rect 442794 281000 443414 281898
rect 451794 283394 452414 284000
rect 451794 283158 451826 283394
rect 452062 283158 452146 283394
rect 452382 283158 452414 283394
rect 451794 283074 452414 283158
rect 451794 282838 451826 283074
rect 452062 282838 452146 283074
rect 452382 282838 452414 283074
rect 451794 281000 452414 282838
rect 460794 282454 461414 284000
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 281000 461414 281898
rect 469794 283394 470414 284000
rect 469794 283158 469826 283394
rect 470062 283158 470146 283394
rect 470382 283158 470414 283394
rect 469794 283074 470414 283158
rect 469794 282838 469826 283074
rect 470062 282838 470146 283074
rect 470382 282838 470414 283074
rect 469794 281000 470414 282838
rect 478794 282454 479414 284000
rect 478794 282218 478826 282454
rect 479062 282218 479146 282454
rect 479382 282218 479414 282454
rect 478794 282134 479414 282218
rect 478794 281898 478826 282134
rect 479062 281898 479146 282134
rect 479382 281898 479414 282134
rect 478794 281000 479414 281898
rect 487794 283394 488414 284000
rect 487794 283158 487826 283394
rect 488062 283158 488146 283394
rect 488382 283158 488414 283394
rect 487794 283074 488414 283158
rect 487794 282838 487826 283074
rect 488062 282838 488146 283074
rect 488382 282838 488414 283074
rect 487794 281000 488414 282838
rect 496794 282454 497414 284000
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 281000 497414 281898
rect 505794 283394 506414 284000
rect 505794 283158 505826 283394
rect 506062 283158 506146 283394
rect 506382 283158 506414 283394
rect 505794 283074 506414 283158
rect 505794 282838 505826 283074
rect 506062 282838 506146 283074
rect 506382 282838 506414 283074
rect 505794 281000 506414 282838
rect 514794 282454 515414 284000
rect 514794 282218 514826 282454
rect 515062 282218 515146 282454
rect 515382 282218 515414 282454
rect 514794 282134 515414 282218
rect 514794 281898 514826 282134
rect 515062 281898 515146 282134
rect 515382 281898 515414 282134
rect 514794 281000 515414 281898
rect 523794 283394 524414 284000
rect 523794 283158 523826 283394
rect 524062 283158 524146 283394
rect 524382 283158 524414 283394
rect 523794 283074 524414 283158
rect 523794 282838 523826 283074
rect 524062 282838 524146 283074
rect 524382 282838 524414 283074
rect 523794 281000 524414 282838
rect 532794 282454 533414 284000
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 281000 533414 281898
rect 541794 283394 542414 284000
rect 541794 283158 541826 283394
rect 542062 283158 542146 283394
rect 542382 283158 542414 283394
rect 541794 283074 542414 283158
rect 541794 282838 541826 283074
rect 542062 282838 542146 283074
rect 542382 282838 542414 283074
rect 541794 281000 542414 282838
rect 550794 282454 551414 284000
rect 550794 282218 550826 282454
rect 551062 282218 551146 282454
rect 551382 282218 551414 282454
rect 550794 282134 551414 282218
rect 550794 281898 550826 282134
rect 551062 281898 551146 282134
rect 551382 281898 551414 282134
rect 550794 281000 551414 281898
rect 19910 273454 20230 273486
rect 19910 273218 19952 273454
rect 20188 273218 20230 273454
rect 19910 273134 20230 273218
rect 19910 272898 19952 273134
rect 20188 272898 20230 273134
rect 19910 272866 20230 272898
rect 25840 273454 26160 273486
rect 25840 273218 25882 273454
rect 26118 273218 26160 273454
rect 25840 273134 26160 273218
rect 25840 272898 25882 273134
rect 26118 272898 26160 273134
rect 25840 272866 26160 272898
rect 31771 273454 32091 273486
rect 31771 273218 31813 273454
rect 32049 273218 32091 273454
rect 31771 273134 32091 273218
rect 31771 272898 31813 273134
rect 32049 272898 32091 273134
rect 31771 272866 32091 272898
rect 46910 273454 47230 273486
rect 46910 273218 46952 273454
rect 47188 273218 47230 273454
rect 46910 273134 47230 273218
rect 46910 272898 46952 273134
rect 47188 272898 47230 273134
rect 46910 272866 47230 272898
rect 52840 273454 53160 273486
rect 52840 273218 52882 273454
rect 53118 273218 53160 273454
rect 52840 273134 53160 273218
rect 52840 272898 52882 273134
rect 53118 272898 53160 273134
rect 52840 272866 53160 272898
rect 58771 273454 59091 273486
rect 58771 273218 58813 273454
rect 59049 273218 59091 273454
rect 58771 273134 59091 273218
rect 58771 272898 58813 273134
rect 59049 272898 59091 273134
rect 58771 272866 59091 272898
rect 73910 273454 74230 273486
rect 73910 273218 73952 273454
rect 74188 273218 74230 273454
rect 73910 273134 74230 273218
rect 73910 272898 73952 273134
rect 74188 272898 74230 273134
rect 73910 272866 74230 272898
rect 79840 273454 80160 273486
rect 79840 273218 79882 273454
rect 80118 273218 80160 273454
rect 79840 273134 80160 273218
rect 79840 272898 79882 273134
rect 80118 272898 80160 273134
rect 79840 272866 80160 272898
rect 85771 273454 86091 273486
rect 85771 273218 85813 273454
rect 86049 273218 86091 273454
rect 85771 273134 86091 273218
rect 85771 272898 85813 273134
rect 86049 272898 86091 273134
rect 85771 272866 86091 272898
rect 100910 273454 101230 273486
rect 100910 273218 100952 273454
rect 101188 273218 101230 273454
rect 100910 273134 101230 273218
rect 100910 272898 100952 273134
rect 101188 272898 101230 273134
rect 100910 272866 101230 272898
rect 106840 273454 107160 273486
rect 106840 273218 106882 273454
rect 107118 273218 107160 273454
rect 106840 273134 107160 273218
rect 106840 272898 106882 273134
rect 107118 272898 107160 273134
rect 106840 272866 107160 272898
rect 112771 273454 113091 273486
rect 112771 273218 112813 273454
rect 113049 273218 113091 273454
rect 112771 273134 113091 273218
rect 112771 272898 112813 273134
rect 113049 272898 113091 273134
rect 112771 272866 113091 272898
rect 127910 273454 128230 273486
rect 127910 273218 127952 273454
rect 128188 273218 128230 273454
rect 127910 273134 128230 273218
rect 127910 272898 127952 273134
rect 128188 272898 128230 273134
rect 127910 272866 128230 272898
rect 133840 273454 134160 273486
rect 133840 273218 133882 273454
rect 134118 273218 134160 273454
rect 133840 273134 134160 273218
rect 133840 272898 133882 273134
rect 134118 272898 134160 273134
rect 133840 272866 134160 272898
rect 139771 273454 140091 273486
rect 139771 273218 139813 273454
rect 140049 273218 140091 273454
rect 139771 273134 140091 273218
rect 139771 272898 139813 273134
rect 140049 272898 140091 273134
rect 139771 272866 140091 272898
rect 154910 273454 155230 273486
rect 154910 273218 154952 273454
rect 155188 273218 155230 273454
rect 154910 273134 155230 273218
rect 154910 272898 154952 273134
rect 155188 272898 155230 273134
rect 154910 272866 155230 272898
rect 160840 273454 161160 273486
rect 160840 273218 160882 273454
rect 161118 273218 161160 273454
rect 160840 273134 161160 273218
rect 160840 272898 160882 273134
rect 161118 272898 161160 273134
rect 160840 272866 161160 272898
rect 166771 273454 167091 273486
rect 166771 273218 166813 273454
rect 167049 273218 167091 273454
rect 166771 273134 167091 273218
rect 166771 272898 166813 273134
rect 167049 272898 167091 273134
rect 166771 272866 167091 272898
rect 181910 273454 182230 273486
rect 181910 273218 181952 273454
rect 182188 273218 182230 273454
rect 181910 273134 182230 273218
rect 181910 272898 181952 273134
rect 182188 272898 182230 273134
rect 181910 272866 182230 272898
rect 187840 273454 188160 273486
rect 187840 273218 187882 273454
rect 188118 273218 188160 273454
rect 187840 273134 188160 273218
rect 187840 272898 187882 273134
rect 188118 272898 188160 273134
rect 187840 272866 188160 272898
rect 193771 273454 194091 273486
rect 193771 273218 193813 273454
rect 194049 273218 194091 273454
rect 193771 273134 194091 273218
rect 193771 272898 193813 273134
rect 194049 272898 194091 273134
rect 193771 272866 194091 272898
rect 208910 273454 209230 273486
rect 208910 273218 208952 273454
rect 209188 273218 209230 273454
rect 208910 273134 209230 273218
rect 208910 272898 208952 273134
rect 209188 272898 209230 273134
rect 208910 272866 209230 272898
rect 214840 273454 215160 273486
rect 214840 273218 214882 273454
rect 215118 273218 215160 273454
rect 214840 273134 215160 273218
rect 214840 272898 214882 273134
rect 215118 272898 215160 273134
rect 214840 272866 215160 272898
rect 220771 273454 221091 273486
rect 220771 273218 220813 273454
rect 221049 273218 221091 273454
rect 220771 273134 221091 273218
rect 220771 272898 220813 273134
rect 221049 272898 221091 273134
rect 220771 272866 221091 272898
rect 235910 273454 236230 273486
rect 235910 273218 235952 273454
rect 236188 273218 236230 273454
rect 235910 273134 236230 273218
rect 235910 272898 235952 273134
rect 236188 272898 236230 273134
rect 235910 272866 236230 272898
rect 241840 273454 242160 273486
rect 241840 273218 241882 273454
rect 242118 273218 242160 273454
rect 241840 273134 242160 273218
rect 241840 272898 241882 273134
rect 242118 272898 242160 273134
rect 241840 272866 242160 272898
rect 247771 273454 248091 273486
rect 247771 273218 247813 273454
rect 248049 273218 248091 273454
rect 247771 273134 248091 273218
rect 247771 272898 247813 273134
rect 248049 272898 248091 273134
rect 247771 272866 248091 272898
rect 262910 273454 263230 273486
rect 262910 273218 262952 273454
rect 263188 273218 263230 273454
rect 262910 273134 263230 273218
rect 262910 272898 262952 273134
rect 263188 272898 263230 273134
rect 262910 272866 263230 272898
rect 268840 273454 269160 273486
rect 268840 273218 268882 273454
rect 269118 273218 269160 273454
rect 268840 273134 269160 273218
rect 268840 272898 268882 273134
rect 269118 272898 269160 273134
rect 268840 272866 269160 272898
rect 274771 273454 275091 273486
rect 274771 273218 274813 273454
rect 275049 273218 275091 273454
rect 274771 273134 275091 273218
rect 274771 272898 274813 273134
rect 275049 272898 275091 273134
rect 274771 272866 275091 272898
rect 289910 273454 290230 273486
rect 289910 273218 289952 273454
rect 290188 273218 290230 273454
rect 289910 273134 290230 273218
rect 289910 272898 289952 273134
rect 290188 272898 290230 273134
rect 289910 272866 290230 272898
rect 295840 273454 296160 273486
rect 295840 273218 295882 273454
rect 296118 273218 296160 273454
rect 295840 273134 296160 273218
rect 295840 272898 295882 273134
rect 296118 272898 296160 273134
rect 295840 272866 296160 272898
rect 301771 273454 302091 273486
rect 301771 273218 301813 273454
rect 302049 273218 302091 273454
rect 301771 273134 302091 273218
rect 301771 272898 301813 273134
rect 302049 272898 302091 273134
rect 301771 272866 302091 272898
rect 316910 273454 317230 273486
rect 316910 273218 316952 273454
rect 317188 273218 317230 273454
rect 316910 273134 317230 273218
rect 316910 272898 316952 273134
rect 317188 272898 317230 273134
rect 316910 272866 317230 272898
rect 322840 273454 323160 273486
rect 322840 273218 322882 273454
rect 323118 273218 323160 273454
rect 322840 273134 323160 273218
rect 322840 272898 322882 273134
rect 323118 272898 323160 273134
rect 322840 272866 323160 272898
rect 328771 273454 329091 273486
rect 328771 273218 328813 273454
rect 329049 273218 329091 273454
rect 328771 273134 329091 273218
rect 328771 272898 328813 273134
rect 329049 272898 329091 273134
rect 328771 272866 329091 272898
rect 343910 273454 344230 273486
rect 343910 273218 343952 273454
rect 344188 273218 344230 273454
rect 343910 273134 344230 273218
rect 343910 272898 343952 273134
rect 344188 272898 344230 273134
rect 343910 272866 344230 272898
rect 349840 273454 350160 273486
rect 349840 273218 349882 273454
rect 350118 273218 350160 273454
rect 349840 273134 350160 273218
rect 349840 272898 349882 273134
rect 350118 272898 350160 273134
rect 349840 272866 350160 272898
rect 355771 273454 356091 273486
rect 355771 273218 355813 273454
rect 356049 273218 356091 273454
rect 355771 273134 356091 273218
rect 355771 272898 355813 273134
rect 356049 272898 356091 273134
rect 355771 272866 356091 272898
rect 370910 273454 371230 273486
rect 370910 273218 370952 273454
rect 371188 273218 371230 273454
rect 370910 273134 371230 273218
rect 370910 272898 370952 273134
rect 371188 272898 371230 273134
rect 370910 272866 371230 272898
rect 376840 273454 377160 273486
rect 376840 273218 376882 273454
rect 377118 273218 377160 273454
rect 376840 273134 377160 273218
rect 376840 272898 376882 273134
rect 377118 272898 377160 273134
rect 376840 272866 377160 272898
rect 382771 273454 383091 273486
rect 382771 273218 382813 273454
rect 383049 273218 383091 273454
rect 382771 273134 383091 273218
rect 382771 272898 382813 273134
rect 383049 272898 383091 273134
rect 382771 272866 383091 272898
rect 397910 273454 398230 273486
rect 397910 273218 397952 273454
rect 398188 273218 398230 273454
rect 397910 273134 398230 273218
rect 397910 272898 397952 273134
rect 398188 272898 398230 273134
rect 397910 272866 398230 272898
rect 403840 273454 404160 273486
rect 403840 273218 403882 273454
rect 404118 273218 404160 273454
rect 403840 273134 404160 273218
rect 403840 272898 403882 273134
rect 404118 272898 404160 273134
rect 403840 272866 404160 272898
rect 409771 273454 410091 273486
rect 409771 273218 409813 273454
rect 410049 273218 410091 273454
rect 409771 273134 410091 273218
rect 409771 272898 409813 273134
rect 410049 272898 410091 273134
rect 409771 272866 410091 272898
rect 424910 273454 425230 273486
rect 424910 273218 424952 273454
rect 425188 273218 425230 273454
rect 424910 273134 425230 273218
rect 424910 272898 424952 273134
rect 425188 272898 425230 273134
rect 424910 272866 425230 272898
rect 430840 273454 431160 273486
rect 430840 273218 430882 273454
rect 431118 273218 431160 273454
rect 430840 273134 431160 273218
rect 430840 272898 430882 273134
rect 431118 272898 431160 273134
rect 430840 272866 431160 272898
rect 436771 273454 437091 273486
rect 436771 273218 436813 273454
rect 437049 273218 437091 273454
rect 436771 273134 437091 273218
rect 436771 272898 436813 273134
rect 437049 272898 437091 273134
rect 436771 272866 437091 272898
rect 451910 273454 452230 273486
rect 451910 273218 451952 273454
rect 452188 273218 452230 273454
rect 451910 273134 452230 273218
rect 451910 272898 451952 273134
rect 452188 272898 452230 273134
rect 451910 272866 452230 272898
rect 457840 273454 458160 273486
rect 457840 273218 457882 273454
rect 458118 273218 458160 273454
rect 457840 273134 458160 273218
rect 457840 272898 457882 273134
rect 458118 272898 458160 273134
rect 457840 272866 458160 272898
rect 463771 273454 464091 273486
rect 463771 273218 463813 273454
rect 464049 273218 464091 273454
rect 463771 273134 464091 273218
rect 463771 272898 463813 273134
rect 464049 272898 464091 273134
rect 463771 272866 464091 272898
rect 478910 273454 479230 273486
rect 478910 273218 478952 273454
rect 479188 273218 479230 273454
rect 478910 273134 479230 273218
rect 478910 272898 478952 273134
rect 479188 272898 479230 273134
rect 478910 272866 479230 272898
rect 484840 273454 485160 273486
rect 484840 273218 484882 273454
rect 485118 273218 485160 273454
rect 484840 273134 485160 273218
rect 484840 272898 484882 273134
rect 485118 272898 485160 273134
rect 484840 272866 485160 272898
rect 490771 273454 491091 273486
rect 490771 273218 490813 273454
rect 491049 273218 491091 273454
rect 490771 273134 491091 273218
rect 490771 272898 490813 273134
rect 491049 272898 491091 273134
rect 490771 272866 491091 272898
rect 505910 273454 506230 273486
rect 505910 273218 505952 273454
rect 506188 273218 506230 273454
rect 505910 273134 506230 273218
rect 505910 272898 505952 273134
rect 506188 272898 506230 273134
rect 505910 272866 506230 272898
rect 511840 273454 512160 273486
rect 511840 273218 511882 273454
rect 512118 273218 512160 273454
rect 511840 273134 512160 273218
rect 511840 272898 511882 273134
rect 512118 272898 512160 273134
rect 511840 272866 512160 272898
rect 517771 273454 518091 273486
rect 517771 273218 517813 273454
rect 518049 273218 518091 273454
rect 517771 273134 518091 273218
rect 517771 272898 517813 273134
rect 518049 272898 518091 273134
rect 517771 272866 518091 272898
rect 532910 273454 533230 273486
rect 532910 273218 532952 273454
rect 533188 273218 533230 273454
rect 532910 273134 533230 273218
rect 532910 272898 532952 273134
rect 533188 272898 533230 273134
rect 532910 272866 533230 272898
rect 538840 273454 539160 273486
rect 538840 273218 538882 273454
rect 539118 273218 539160 273454
rect 538840 273134 539160 273218
rect 538840 272898 538882 273134
rect 539118 272898 539160 273134
rect 538840 272866 539160 272898
rect 544771 273454 545091 273486
rect 544771 273218 544813 273454
rect 545049 273218 545091 273454
rect 544771 273134 545091 273218
rect 544771 272898 544813 273134
rect 545049 272898 545091 273134
rect 544771 272866 545091 272898
rect 559794 273454 560414 290898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 246454 11414 263898
rect 22874 264454 23194 264486
rect 22874 264218 22916 264454
rect 23152 264218 23194 264454
rect 22874 264134 23194 264218
rect 22874 263898 22916 264134
rect 23152 263898 23194 264134
rect 22874 263866 23194 263898
rect 28805 264454 29125 264486
rect 28805 264218 28847 264454
rect 29083 264218 29125 264454
rect 28805 264134 29125 264218
rect 28805 263898 28847 264134
rect 29083 263898 29125 264134
rect 28805 263866 29125 263898
rect 49874 264454 50194 264486
rect 49874 264218 49916 264454
rect 50152 264218 50194 264454
rect 49874 264134 50194 264218
rect 49874 263898 49916 264134
rect 50152 263898 50194 264134
rect 49874 263866 50194 263898
rect 55805 264454 56125 264486
rect 55805 264218 55847 264454
rect 56083 264218 56125 264454
rect 55805 264134 56125 264218
rect 55805 263898 55847 264134
rect 56083 263898 56125 264134
rect 55805 263866 56125 263898
rect 76874 264454 77194 264486
rect 76874 264218 76916 264454
rect 77152 264218 77194 264454
rect 76874 264134 77194 264218
rect 76874 263898 76916 264134
rect 77152 263898 77194 264134
rect 76874 263866 77194 263898
rect 82805 264454 83125 264486
rect 82805 264218 82847 264454
rect 83083 264218 83125 264454
rect 82805 264134 83125 264218
rect 82805 263898 82847 264134
rect 83083 263898 83125 264134
rect 82805 263866 83125 263898
rect 103874 264454 104194 264486
rect 103874 264218 103916 264454
rect 104152 264218 104194 264454
rect 103874 264134 104194 264218
rect 103874 263898 103916 264134
rect 104152 263898 104194 264134
rect 103874 263866 104194 263898
rect 109805 264454 110125 264486
rect 109805 264218 109847 264454
rect 110083 264218 110125 264454
rect 109805 264134 110125 264218
rect 109805 263898 109847 264134
rect 110083 263898 110125 264134
rect 109805 263866 110125 263898
rect 130874 264454 131194 264486
rect 130874 264218 130916 264454
rect 131152 264218 131194 264454
rect 130874 264134 131194 264218
rect 130874 263898 130916 264134
rect 131152 263898 131194 264134
rect 130874 263866 131194 263898
rect 136805 264454 137125 264486
rect 136805 264218 136847 264454
rect 137083 264218 137125 264454
rect 136805 264134 137125 264218
rect 136805 263898 136847 264134
rect 137083 263898 137125 264134
rect 136805 263866 137125 263898
rect 157874 264454 158194 264486
rect 157874 264218 157916 264454
rect 158152 264218 158194 264454
rect 157874 264134 158194 264218
rect 157874 263898 157916 264134
rect 158152 263898 158194 264134
rect 157874 263866 158194 263898
rect 163805 264454 164125 264486
rect 163805 264218 163847 264454
rect 164083 264218 164125 264454
rect 163805 264134 164125 264218
rect 163805 263898 163847 264134
rect 164083 263898 164125 264134
rect 163805 263866 164125 263898
rect 184874 264454 185194 264486
rect 184874 264218 184916 264454
rect 185152 264218 185194 264454
rect 184874 264134 185194 264218
rect 184874 263898 184916 264134
rect 185152 263898 185194 264134
rect 184874 263866 185194 263898
rect 190805 264454 191125 264486
rect 190805 264218 190847 264454
rect 191083 264218 191125 264454
rect 190805 264134 191125 264218
rect 190805 263898 190847 264134
rect 191083 263898 191125 264134
rect 190805 263866 191125 263898
rect 211874 264454 212194 264486
rect 211874 264218 211916 264454
rect 212152 264218 212194 264454
rect 211874 264134 212194 264218
rect 211874 263898 211916 264134
rect 212152 263898 212194 264134
rect 211874 263866 212194 263898
rect 217805 264454 218125 264486
rect 217805 264218 217847 264454
rect 218083 264218 218125 264454
rect 217805 264134 218125 264218
rect 217805 263898 217847 264134
rect 218083 263898 218125 264134
rect 217805 263866 218125 263898
rect 238874 264454 239194 264486
rect 238874 264218 238916 264454
rect 239152 264218 239194 264454
rect 238874 264134 239194 264218
rect 238874 263898 238916 264134
rect 239152 263898 239194 264134
rect 238874 263866 239194 263898
rect 244805 264454 245125 264486
rect 244805 264218 244847 264454
rect 245083 264218 245125 264454
rect 244805 264134 245125 264218
rect 244805 263898 244847 264134
rect 245083 263898 245125 264134
rect 244805 263866 245125 263898
rect 265874 264454 266194 264486
rect 265874 264218 265916 264454
rect 266152 264218 266194 264454
rect 265874 264134 266194 264218
rect 265874 263898 265916 264134
rect 266152 263898 266194 264134
rect 265874 263866 266194 263898
rect 271805 264454 272125 264486
rect 271805 264218 271847 264454
rect 272083 264218 272125 264454
rect 271805 264134 272125 264218
rect 271805 263898 271847 264134
rect 272083 263898 272125 264134
rect 271805 263866 272125 263898
rect 292874 264454 293194 264486
rect 292874 264218 292916 264454
rect 293152 264218 293194 264454
rect 292874 264134 293194 264218
rect 292874 263898 292916 264134
rect 293152 263898 293194 264134
rect 292874 263866 293194 263898
rect 298805 264454 299125 264486
rect 298805 264218 298847 264454
rect 299083 264218 299125 264454
rect 298805 264134 299125 264218
rect 298805 263898 298847 264134
rect 299083 263898 299125 264134
rect 298805 263866 299125 263898
rect 319874 264454 320194 264486
rect 319874 264218 319916 264454
rect 320152 264218 320194 264454
rect 319874 264134 320194 264218
rect 319874 263898 319916 264134
rect 320152 263898 320194 264134
rect 319874 263866 320194 263898
rect 325805 264454 326125 264486
rect 325805 264218 325847 264454
rect 326083 264218 326125 264454
rect 325805 264134 326125 264218
rect 325805 263898 325847 264134
rect 326083 263898 326125 264134
rect 325805 263866 326125 263898
rect 346874 264454 347194 264486
rect 346874 264218 346916 264454
rect 347152 264218 347194 264454
rect 346874 264134 347194 264218
rect 346874 263898 346916 264134
rect 347152 263898 347194 264134
rect 346874 263866 347194 263898
rect 352805 264454 353125 264486
rect 352805 264218 352847 264454
rect 353083 264218 353125 264454
rect 352805 264134 353125 264218
rect 352805 263898 352847 264134
rect 353083 263898 353125 264134
rect 352805 263866 353125 263898
rect 373874 264454 374194 264486
rect 373874 264218 373916 264454
rect 374152 264218 374194 264454
rect 373874 264134 374194 264218
rect 373874 263898 373916 264134
rect 374152 263898 374194 264134
rect 373874 263866 374194 263898
rect 379805 264454 380125 264486
rect 379805 264218 379847 264454
rect 380083 264218 380125 264454
rect 379805 264134 380125 264218
rect 379805 263898 379847 264134
rect 380083 263898 380125 264134
rect 379805 263866 380125 263898
rect 400874 264454 401194 264486
rect 400874 264218 400916 264454
rect 401152 264218 401194 264454
rect 400874 264134 401194 264218
rect 400874 263898 400916 264134
rect 401152 263898 401194 264134
rect 400874 263866 401194 263898
rect 406805 264454 407125 264486
rect 406805 264218 406847 264454
rect 407083 264218 407125 264454
rect 406805 264134 407125 264218
rect 406805 263898 406847 264134
rect 407083 263898 407125 264134
rect 406805 263866 407125 263898
rect 427874 264454 428194 264486
rect 427874 264218 427916 264454
rect 428152 264218 428194 264454
rect 427874 264134 428194 264218
rect 427874 263898 427916 264134
rect 428152 263898 428194 264134
rect 427874 263866 428194 263898
rect 433805 264454 434125 264486
rect 433805 264218 433847 264454
rect 434083 264218 434125 264454
rect 433805 264134 434125 264218
rect 433805 263898 433847 264134
rect 434083 263898 434125 264134
rect 433805 263866 434125 263898
rect 454874 264454 455194 264486
rect 454874 264218 454916 264454
rect 455152 264218 455194 264454
rect 454874 264134 455194 264218
rect 454874 263898 454916 264134
rect 455152 263898 455194 264134
rect 454874 263866 455194 263898
rect 460805 264454 461125 264486
rect 460805 264218 460847 264454
rect 461083 264218 461125 264454
rect 460805 264134 461125 264218
rect 460805 263898 460847 264134
rect 461083 263898 461125 264134
rect 460805 263866 461125 263898
rect 481874 264454 482194 264486
rect 481874 264218 481916 264454
rect 482152 264218 482194 264454
rect 481874 264134 482194 264218
rect 481874 263898 481916 264134
rect 482152 263898 482194 264134
rect 481874 263866 482194 263898
rect 487805 264454 488125 264486
rect 487805 264218 487847 264454
rect 488083 264218 488125 264454
rect 487805 264134 488125 264218
rect 487805 263898 487847 264134
rect 488083 263898 488125 264134
rect 487805 263866 488125 263898
rect 508874 264454 509194 264486
rect 508874 264218 508916 264454
rect 509152 264218 509194 264454
rect 508874 264134 509194 264218
rect 508874 263898 508916 264134
rect 509152 263898 509194 264134
rect 508874 263866 509194 263898
rect 514805 264454 515125 264486
rect 514805 264218 514847 264454
rect 515083 264218 515125 264454
rect 514805 264134 515125 264218
rect 514805 263898 514847 264134
rect 515083 263898 515125 264134
rect 514805 263866 515125 263898
rect 535874 264454 536194 264486
rect 535874 264218 535916 264454
rect 536152 264218 536194 264454
rect 535874 264134 536194 264218
rect 535874 263898 535916 264134
rect 536152 263898 536194 264134
rect 535874 263866 536194 263898
rect 541805 264454 542125 264486
rect 541805 264218 541847 264454
rect 542083 264218 542125 264454
rect 541805 264134 542125 264218
rect 541805 263898 541847 264134
rect 542083 263898 542125 264134
rect 541805 263866 542125 263898
rect 19794 255454 20414 257000
rect 19794 255218 19826 255454
rect 20062 255218 20146 255454
rect 20382 255218 20414 255454
rect 19794 255134 20414 255218
rect 19794 254898 19826 255134
rect 20062 254898 20146 255134
rect 20382 254898 20414 255134
rect 19794 254000 20414 254898
rect 28794 256394 29414 257000
rect 28794 256158 28826 256394
rect 29062 256158 29146 256394
rect 29382 256158 29414 256394
rect 28794 256074 29414 256158
rect 28794 255838 28826 256074
rect 29062 255838 29146 256074
rect 29382 255838 29414 256074
rect 28794 254000 29414 255838
rect 37794 255454 38414 257000
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 254000 38414 254898
rect 46794 256394 47414 257000
rect 46794 256158 46826 256394
rect 47062 256158 47146 256394
rect 47382 256158 47414 256394
rect 46794 256074 47414 256158
rect 46794 255838 46826 256074
rect 47062 255838 47146 256074
rect 47382 255838 47414 256074
rect 46794 254000 47414 255838
rect 55794 255454 56414 257000
rect 55794 255218 55826 255454
rect 56062 255218 56146 255454
rect 56382 255218 56414 255454
rect 55794 255134 56414 255218
rect 55794 254898 55826 255134
rect 56062 254898 56146 255134
rect 56382 254898 56414 255134
rect 55794 254000 56414 254898
rect 64794 256394 65414 257000
rect 64794 256158 64826 256394
rect 65062 256158 65146 256394
rect 65382 256158 65414 256394
rect 64794 256074 65414 256158
rect 64794 255838 64826 256074
rect 65062 255838 65146 256074
rect 65382 255838 65414 256074
rect 64794 254000 65414 255838
rect 73794 255454 74414 257000
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 254000 74414 254898
rect 82794 256394 83414 257000
rect 82794 256158 82826 256394
rect 83062 256158 83146 256394
rect 83382 256158 83414 256394
rect 82794 256074 83414 256158
rect 82794 255838 82826 256074
rect 83062 255838 83146 256074
rect 83382 255838 83414 256074
rect 82794 254000 83414 255838
rect 91794 255454 92414 257000
rect 91794 255218 91826 255454
rect 92062 255218 92146 255454
rect 92382 255218 92414 255454
rect 91794 255134 92414 255218
rect 91794 254898 91826 255134
rect 92062 254898 92146 255134
rect 92382 254898 92414 255134
rect 91794 254000 92414 254898
rect 100794 256394 101414 257000
rect 100794 256158 100826 256394
rect 101062 256158 101146 256394
rect 101382 256158 101414 256394
rect 100794 256074 101414 256158
rect 100794 255838 100826 256074
rect 101062 255838 101146 256074
rect 101382 255838 101414 256074
rect 100794 254000 101414 255838
rect 109794 255454 110414 257000
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 254000 110414 254898
rect 118794 256394 119414 257000
rect 118794 256158 118826 256394
rect 119062 256158 119146 256394
rect 119382 256158 119414 256394
rect 118794 256074 119414 256158
rect 118794 255838 118826 256074
rect 119062 255838 119146 256074
rect 119382 255838 119414 256074
rect 118794 254000 119414 255838
rect 127794 255454 128414 257000
rect 127794 255218 127826 255454
rect 128062 255218 128146 255454
rect 128382 255218 128414 255454
rect 127794 255134 128414 255218
rect 127794 254898 127826 255134
rect 128062 254898 128146 255134
rect 128382 254898 128414 255134
rect 127794 254000 128414 254898
rect 136794 256394 137414 257000
rect 136794 256158 136826 256394
rect 137062 256158 137146 256394
rect 137382 256158 137414 256394
rect 136794 256074 137414 256158
rect 136794 255838 136826 256074
rect 137062 255838 137146 256074
rect 137382 255838 137414 256074
rect 136794 254000 137414 255838
rect 145794 255454 146414 257000
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 254000 146414 254898
rect 154794 256394 155414 257000
rect 154794 256158 154826 256394
rect 155062 256158 155146 256394
rect 155382 256158 155414 256394
rect 154794 256074 155414 256158
rect 154794 255838 154826 256074
rect 155062 255838 155146 256074
rect 155382 255838 155414 256074
rect 154794 254000 155414 255838
rect 163794 255454 164414 257000
rect 163794 255218 163826 255454
rect 164062 255218 164146 255454
rect 164382 255218 164414 255454
rect 163794 255134 164414 255218
rect 163794 254898 163826 255134
rect 164062 254898 164146 255134
rect 164382 254898 164414 255134
rect 163794 254000 164414 254898
rect 172794 256394 173414 257000
rect 172794 256158 172826 256394
rect 173062 256158 173146 256394
rect 173382 256158 173414 256394
rect 172794 256074 173414 256158
rect 172794 255838 172826 256074
rect 173062 255838 173146 256074
rect 173382 255838 173414 256074
rect 172794 254000 173414 255838
rect 181794 255454 182414 257000
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 254000 182414 254898
rect 190794 256394 191414 257000
rect 190794 256158 190826 256394
rect 191062 256158 191146 256394
rect 191382 256158 191414 256394
rect 190794 256074 191414 256158
rect 190794 255838 190826 256074
rect 191062 255838 191146 256074
rect 191382 255838 191414 256074
rect 190794 254000 191414 255838
rect 199794 255454 200414 257000
rect 199794 255218 199826 255454
rect 200062 255218 200146 255454
rect 200382 255218 200414 255454
rect 199794 255134 200414 255218
rect 199794 254898 199826 255134
rect 200062 254898 200146 255134
rect 200382 254898 200414 255134
rect 199794 254000 200414 254898
rect 208794 256394 209414 257000
rect 208794 256158 208826 256394
rect 209062 256158 209146 256394
rect 209382 256158 209414 256394
rect 208794 256074 209414 256158
rect 208794 255838 208826 256074
rect 209062 255838 209146 256074
rect 209382 255838 209414 256074
rect 208794 254000 209414 255838
rect 217794 255454 218414 257000
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 254000 218414 254898
rect 226794 256394 227414 257000
rect 226794 256158 226826 256394
rect 227062 256158 227146 256394
rect 227382 256158 227414 256394
rect 226794 256074 227414 256158
rect 226794 255838 226826 256074
rect 227062 255838 227146 256074
rect 227382 255838 227414 256074
rect 226794 254000 227414 255838
rect 235794 255454 236414 257000
rect 235794 255218 235826 255454
rect 236062 255218 236146 255454
rect 236382 255218 236414 255454
rect 235794 255134 236414 255218
rect 235794 254898 235826 255134
rect 236062 254898 236146 255134
rect 236382 254898 236414 255134
rect 235794 254000 236414 254898
rect 244794 256394 245414 257000
rect 244794 256158 244826 256394
rect 245062 256158 245146 256394
rect 245382 256158 245414 256394
rect 244794 256074 245414 256158
rect 244794 255838 244826 256074
rect 245062 255838 245146 256074
rect 245382 255838 245414 256074
rect 244794 254000 245414 255838
rect 253794 255454 254414 257000
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 254000 254414 254898
rect 262794 256394 263414 257000
rect 262794 256158 262826 256394
rect 263062 256158 263146 256394
rect 263382 256158 263414 256394
rect 262794 256074 263414 256158
rect 262794 255838 262826 256074
rect 263062 255838 263146 256074
rect 263382 255838 263414 256074
rect 262794 254000 263414 255838
rect 271794 255454 272414 257000
rect 271794 255218 271826 255454
rect 272062 255218 272146 255454
rect 272382 255218 272414 255454
rect 271794 255134 272414 255218
rect 271794 254898 271826 255134
rect 272062 254898 272146 255134
rect 272382 254898 272414 255134
rect 271794 254000 272414 254898
rect 280794 256394 281414 257000
rect 280794 256158 280826 256394
rect 281062 256158 281146 256394
rect 281382 256158 281414 256394
rect 280794 256074 281414 256158
rect 280794 255838 280826 256074
rect 281062 255838 281146 256074
rect 281382 255838 281414 256074
rect 280794 254000 281414 255838
rect 289794 255454 290414 257000
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 254000 290414 254898
rect 298794 256394 299414 257000
rect 298794 256158 298826 256394
rect 299062 256158 299146 256394
rect 299382 256158 299414 256394
rect 298794 256074 299414 256158
rect 298794 255838 298826 256074
rect 299062 255838 299146 256074
rect 299382 255838 299414 256074
rect 298794 254000 299414 255838
rect 307794 255454 308414 257000
rect 307794 255218 307826 255454
rect 308062 255218 308146 255454
rect 308382 255218 308414 255454
rect 307794 255134 308414 255218
rect 307794 254898 307826 255134
rect 308062 254898 308146 255134
rect 308382 254898 308414 255134
rect 307794 254000 308414 254898
rect 316794 256394 317414 257000
rect 316794 256158 316826 256394
rect 317062 256158 317146 256394
rect 317382 256158 317414 256394
rect 316794 256074 317414 256158
rect 316794 255838 316826 256074
rect 317062 255838 317146 256074
rect 317382 255838 317414 256074
rect 316794 254000 317414 255838
rect 325794 255454 326414 257000
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 254000 326414 254898
rect 334794 256394 335414 257000
rect 334794 256158 334826 256394
rect 335062 256158 335146 256394
rect 335382 256158 335414 256394
rect 334794 256074 335414 256158
rect 334794 255838 334826 256074
rect 335062 255838 335146 256074
rect 335382 255838 335414 256074
rect 334794 254000 335414 255838
rect 343794 255454 344414 257000
rect 343794 255218 343826 255454
rect 344062 255218 344146 255454
rect 344382 255218 344414 255454
rect 343794 255134 344414 255218
rect 343794 254898 343826 255134
rect 344062 254898 344146 255134
rect 344382 254898 344414 255134
rect 343794 254000 344414 254898
rect 352794 256394 353414 257000
rect 352794 256158 352826 256394
rect 353062 256158 353146 256394
rect 353382 256158 353414 256394
rect 352794 256074 353414 256158
rect 352794 255838 352826 256074
rect 353062 255838 353146 256074
rect 353382 255838 353414 256074
rect 352794 254000 353414 255838
rect 361794 255454 362414 257000
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 254000 362414 254898
rect 370794 256394 371414 257000
rect 370794 256158 370826 256394
rect 371062 256158 371146 256394
rect 371382 256158 371414 256394
rect 370794 256074 371414 256158
rect 370794 255838 370826 256074
rect 371062 255838 371146 256074
rect 371382 255838 371414 256074
rect 370794 254000 371414 255838
rect 379794 255454 380414 257000
rect 379794 255218 379826 255454
rect 380062 255218 380146 255454
rect 380382 255218 380414 255454
rect 379794 255134 380414 255218
rect 379794 254898 379826 255134
rect 380062 254898 380146 255134
rect 380382 254898 380414 255134
rect 379794 254000 380414 254898
rect 388794 256394 389414 257000
rect 388794 256158 388826 256394
rect 389062 256158 389146 256394
rect 389382 256158 389414 256394
rect 388794 256074 389414 256158
rect 388794 255838 388826 256074
rect 389062 255838 389146 256074
rect 389382 255838 389414 256074
rect 388794 254000 389414 255838
rect 397794 255454 398414 257000
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 254000 398414 254898
rect 406794 256394 407414 257000
rect 406794 256158 406826 256394
rect 407062 256158 407146 256394
rect 407382 256158 407414 256394
rect 406794 256074 407414 256158
rect 406794 255838 406826 256074
rect 407062 255838 407146 256074
rect 407382 255838 407414 256074
rect 406794 254000 407414 255838
rect 415794 255454 416414 257000
rect 415794 255218 415826 255454
rect 416062 255218 416146 255454
rect 416382 255218 416414 255454
rect 415794 255134 416414 255218
rect 415794 254898 415826 255134
rect 416062 254898 416146 255134
rect 416382 254898 416414 255134
rect 415794 254000 416414 254898
rect 424794 256394 425414 257000
rect 424794 256158 424826 256394
rect 425062 256158 425146 256394
rect 425382 256158 425414 256394
rect 424794 256074 425414 256158
rect 424794 255838 424826 256074
rect 425062 255838 425146 256074
rect 425382 255838 425414 256074
rect 424794 254000 425414 255838
rect 433794 255454 434414 257000
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 254000 434414 254898
rect 442794 256394 443414 257000
rect 442794 256158 442826 256394
rect 443062 256158 443146 256394
rect 443382 256158 443414 256394
rect 442794 256074 443414 256158
rect 442794 255838 442826 256074
rect 443062 255838 443146 256074
rect 443382 255838 443414 256074
rect 442794 254000 443414 255838
rect 451794 255454 452414 257000
rect 451794 255218 451826 255454
rect 452062 255218 452146 255454
rect 452382 255218 452414 255454
rect 451794 255134 452414 255218
rect 451794 254898 451826 255134
rect 452062 254898 452146 255134
rect 452382 254898 452414 255134
rect 451794 254000 452414 254898
rect 460794 256394 461414 257000
rect 460794 256158 460826 256394
rect 461062 256158 461146 256394
rect 461382 256158 461414 256394
rect 460794 256074 461414 256158
rect 460794 255838 460826 256074
rect 461062 255838 461146 256074
rect 461382 255838 461414 256074
rect 460794 254000 461414 255838
rect 469794 255454 470414 257000
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 254000 470414 254898
rect 478794 256394 479414 257000
rect 478794 256158 478826 256394
rect 479062 256158 479146 256394
rect 479382 256158 479414 256394
rect 478794 256074 479414 256158
rect 478794 255838 478826 256074
rect 479062 255838 479146 256074
rect 479382 255838 479414 256074
rect 478794 254000 479414 255838
rect 487794 255454 488414 257000
rect 487794 255218 487826 255454
rect 488062 255218 488146 255454
rect 488382 255218 488414 255454
rect 487794 255134 488414 255218
rect 487794 254898 487826 255134
rect 488062 254898 488146 255134
rect 488382 254898 488414 255134
rect 487794 254000 488414 254898
rect 496794 256394 497414 257000
rect 496794 256158 496826 256394
rect 497062 256158 497146 256394
rect 497382 256158 497414 256394
rect 496794 256074 497414 256158
rect 496794 255838 496826 256074
rect 497062 255838 497146 256074
rect 497382 255838 497414 256074
rect 496794 254000 497414 255838
rect 505794 255454 506414 257000
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 254000 506414 254898
rect 514794 256394 515414 257000
rect 514794 256158 514826 256394
rect 515062 256158 515146 256394
rect 515382 256158 515414 256394
rect 514794 256074 515414 256158
rect 514794 255838 514826 256074
rect 515062 255838 515146 256074
rect 515382 255838 515414 256074
rect 514794 254000 515414 255838
rect 523794 255454 524414 257000
rect 523794 255218 523826 255454
rect 524062 255218 524146 255454
rect 524382 255218 524414 255454
rect 523794 255134 524414 255218
rect 523794 254898 523826 255134
rect 524062 254898 524146 255134
rect 524382 254898 524414 255134
rect 523794 254000 524414 254898
rect 532794 256394 533414 257000
rect 532794 256158 532826 256394
rect 533062 256158 533146 256394
rect 533382 256158 533414 256394
rect 532794 256074 533414 256158
rect 532794 255838 532826 256074
rect 533062 255838 533146 256074
rect 533382 255838 533414 256074
rect 532794 254000 533414 255838
rect 541794 255454 542414 257000
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 254000 542414 254898
rect 550794 256394 551414 257000
rect 550794 256158 550826 256394
rect 551062 256158 551146 256394
rect 551382 256158 551414 256394
rect 550794 256074 551414 256158
rect 550794 255838 550826 256074
rect 551062 255838 551146 256074
rect 551382 255838 551414 256074
rect 550794 254000 551414 255838
rect 559794 255454 560414 272898
rect 559794 255218 559826 255454
rect 560062 255218 560146 255454
rect 560382 255218 560414 255454
rect 559794 255134 560414 255218
rect 559794 254898 559826 255134
rect 560062 254898 560146 255134
rect 560382 254898 560414 255134
rect 10794 246218 10826 246454
rect 11062 246218 11146 246454
rect 11382 246218 11414 246454
rect 10794 246134 11414 246218
rect 10794 245898 10826 246134
rect 11062 245898 11146 246134
rect 11382 245898 11414 246134
rect 10794 228454 11414 245898
rect 22874 246454 23194 246486
rect 22874 246218 22916 246454
rect 23152 246218 23194 246454
rect 22874 246134 23194 246218
rect 22874 245898 22916 246134
rect 23152 245898 23194 246134
rect 22874 245866 23194 245898
rect 28805 246454 29125 246486
rect 28805 246218 28847 246454
rect 29083 246218 29125 246454
rect 28805 246134 29125 246218
rect 28805 245898 28847 246134
rect 29083 245898 29125 246134
rect 28805 245866 29125 245898
rect 49874 246454 50194 246486
rect 49874 246218 49916 246454
rect 50152 246218 50194 246454
rect 49874 246134 50194 246218
rect 49874 245898 49916 246134
rect 50152 245898 50194 246134
rect 49874 245866 50194 245898
rect 55805 246454 56125 246486
rect 55805 246218 55847 246454
rect 56083 246218 56125 246454
rect 55805 246134 56125 246218
rect 55805 245898 55847 246134
rect 56083 245898 56125 246134
rect 55805 245866 56125 245898
rect 76874 246454 77194 246486
rect 76874 246218 76916 246454
rect 77152 246218 77194 246454
rect 76874 246134 77194 246218
rect 76874 245898 76916 246134
rect 77152 245898 77194 246134
rect 76874 245866 77194 245898
rect 82805 246454 83125 246486
rect 82805 246218 82847 246454
rect 83083 246218 83125 246454
rect 82805 246134 83125 246218
rect 82805 245898 82847 246134
rect 83083 245898 83125 246134
rect 82805 245866 83125 245898
rect 103874 246454 104194 246486
rect 103874 246218 103916 246454
rect 104152 246218 104194 246454
rect 103874 246134 104194 246218
rect 103874 245898 103916 246134
rect 104152 245898 104194 246134
rect 103874 245866 104194 245898
rect 109805 246454 110125 246486
rect 109805 246218 109847 246454
rect 110083 246218 110125 246454
rect 109805 246134 110125 246218
rect 109805 245898 109847 246134
rect 110083 245898 110125 246134
rect 109805 245866 110125 245898
rect 130874 246454 131194 246486
rect 130874 246218 130916 246454
rect 131152 246218 131194 246454
rect 130874 246134 131194 246218
rect 130874 245898 130916 246134
rect 131152 245898 131194 246134
rect 130874 245866 131194 245898
rect 136805 246454 137125 246486
rect 136805 246218 136847 246454
rect 137083 246218 137125 246454
rect 136805 246134 137125 246218
rect 136805 245898 136847 246134
rect 137083 245898 137125 246134
rect 136805 245866 137125 245898
rect 157874 246454 158194 246486
rect 157874 246218 157916 246454
rect 158152 246218 158194 246454
rect 157874 246134 158194 246218
rect 157874 245898 157916 246134
rect 158152 245898 158194 246134
rect 157874 245866 158194 245898
rect 163805 246454 164125 246486
rect 163805 246218 163847 246454
rect 164083 246218 164125 246454
rect 163805 246134 164125 246218
rect 163805 245898 163847 246134
rect 164083 245898 164125 246134
rect 163805 245866 164125 245898
rect 184874 246454 185194 246486
rect 184874 246218 184916 246454
rect 185152 246218 185194 246454
rect 184874 246134 185194 246218
rect 184874 245898 184916 246134
rect 185152 245898 185194 246134
rect 184874 245866 185194 245898
rect 190805 246454 191125 246486
rect 190805 246218 190847 246454
rect 191083 246218 191125 246454
rect 190805 246134 191125 246218
rect 190805 245898 190847 246134
rect 191083 245898 191125 246134
rect 190805 245866 191125 245898
rect 211874 246454 212194 246486
rect 211874 246218 211916 246454
rect 212152 246218 212194 246454
rect 211874 246134 212194 246218
rect 211874 245898 211916 246134
rect 212152 245898 212194 246134
rect 211874 245866 212194 245898
rect 217805 246454 218125 246486
rect 217805 246218 217847 246454
rect 218083 246218 218125 246454
rect 217805 246134 218125 246218
rect 217805 245898 217847 246134
rect 218083 245898 218125 246134
rect 217805 245866 218125 245898
rect 238874 246454 239194 246486
rect 238874 246218 238916 246454
rect 239152 246218 239194 246454
rect 238874 246134 239194 246218
rect 238874 245898 238916 246134
rect 239152 245898 239194 246134
rect 238874 245866 239194 245898
rect 244805 246454 245125 246486
rect 244805 246218 244847 246454
rect 245083 246218 245125 246454
rect 244805 246134 245125 246218
rect 244805 245898 244847 246134
rect 245083 245898 245125 246134
rect 244805 245866 245125 245898
rect 265874 246454 266194 246486
rect 265874 246218 265916 246454
rect 266152 246218 266194 246454
rect 265874 246134 266194 246218
rect 265874 245898 265916 246134
rect 266152 245898 266194 246134
rect 265874 245866 266194 245898
rect 271805 246454 272125 246486
rect 271805 246218 271847 246454
rect 272083 246218 272125 246454
rect 271805 246134 272125 246218
rect 271805 245898 271847 246134
rect 272083 245898 272125 246134
rect 271805 245866 272125 245898
rect 292874 246454 293194 246486
rect 292874 246218 292916 246454
rect 293152 246218 293194 246454
rect 292874 246134 293194 246218
rect 292874 245898 292916 246134
rect 293152 245898 293194 246134
rect 292874 245866 293194 245898
rect 298805 246454 299125 246486
rect 298805 246218 298847 246454
rect 299083 246218 299125 246454
rect 298805 246134 299125 246218
rect 298805 245898 298847 246134
rect 299083 245898 299125 246134
rect 298805 245866 299125 245898
rect 319874 246454 320194 246486
rect 319874 246218 319916 246454
rect 320152 246218 320194 246454
rect 319874 246134 320194 246218
rect 319874 245898 319916 246134
rect 320152 245898 320194 246134
rect 319874 245866 320194 245898
rect 325805 246454 326125 246486
rect 325805 246218 325847 246454
rect 326083 246218 326125 246454
rect 325805 246134 326125 246218
rect 325805 245898 325847 246134
rect 326083 245898 326125 246134
rect 325805 245866 326125 245898
rect 346874 246454 347194 246486
rect 346874 246218 346916 246454
rect 347152 246218 347194 246454
rect 346874 246134 347194 246218
rect 346874 245898 346916 246134
rect 347152 245898 347194 246134
rect 346874 245866 347194 245898
rect 352805 246454 353125 246486
rect 352805 246218 352847 246454
rect 353083 246218 353125 246454
rect 352805 246134 353125 246218
rect 352805 245898 352847 246134
rect 353083 245898 353125 246134
rect 352805 245866 353125 245898
rect 373874 246454 374194 246486
rect 373874 246218 373916 246454
rect 374152 246218 374194 246454
rect 373874 246134 374194 246218
rect 373874 245898 373916 246134
rect 374152 245898 374194 246134
rect 373874 245866 374194 245898
rect 379805 246454 380125 246486
rect 379805 246218 379847 246454
rect 380083 246218 380125 246454
rect 379805 246134 380125 246218
rect 379805 245898 379847 246134
rect 380083 245898 380125 246134
rect 379805 245866 380125 245898
rect 400874 246454 401194 246486
rect 400874 246218 400916 246454
rect 401152 246218 401194 246454
rect 400874 246134 401194 246218
rect 400874 245898 400916 246134
rect 401152 245898 401194 246134
rect 400874 245866 401194 245898
rect 406805 246454 407125 246486
rect 406805 246218 406847 246454
rect 407083 246218 407125 246454
rect 406805 246134 407125 246218
rect 406805 245898 406847 246134
rect 407083 245898 407125 246134
rect 406805 245866 407125 245898
rect 427874 246454 428194 246486
rect 427874 246218 427916 246454
rect 428152 246218 428194 246454
rect 427874 246134 428194 246218
rect 427874 245898 427916 246134
rect 428152 245898 428194 246134
rect 427874 245866 428194 245898
rect 433805 246454 434125 246486
rect 433805 246218 433847 246454
rect 434083 246218 434125 246454
rect 433805 246134 434125 246218
rect 433805 245898 433847 246134
rect 434083 245898 434125 246134
rect 433805 245866 434125 245898
rect 454874 246454 455194 246486
rect 454874 246218 454916 246454
rect 455152 246218 455194 246454
rect 454874 246134 455194 246218
rect 454874 245898 454916 246134
rect 455152 245898 455194 246134
rect 454874 245866 455194 245898
rect 460805 246454 461125 246486
rect 460805 246218 460847 246454
rect 461083 246218 461125 246454
rect 460805 246134 461125 246218
rect 460805 245898 460847 246134
rect 461083 245898 461125 246134
rect 460805 245866 461125 245898
rect 481874 246454 482194 246486
rect 481874 246218 481916 246454
rect 482152 246218 482194 246454
rect 481874 246134 482194 246218
rect 481874 245898 481916 246134
rect 482152 245898 482194 246134
rect 481874 245866 482194 245898
rect 487805 246454 488125 246486
rect 487805 246218 487847 246454
rect 488083 246218 488125 246454
rect 487805 246134 488125 246218
rect 487805 245898 487847 246134
rect 488083 245898 488125 246134
rect 487805 245866 488125 245898
rect 508874 246454 509194 246486
rect 508874 246218 508916 246454
rect 509152 246218 509194 246454
rect 508874 246134 509194 246218
rect 508874 245898 508916 246134
rect 509152 245898 509194 246134
rect 508874 245866 509194 245898
rect 514805 246454 515125 246486
rect 514805 246218 514847 246454
rect 515083 246218 515125 246454
rect 514805 246134 515125 246218
rect 514805 245898 514847 246134
rect 515083 245898 515125 246134
rect 514805 245866 515125 245898
rect 535874 246454 536194 246486
rect 535874 246218 535916 246454
rect 536152 246218 536194 246454
rect 535874 246134 536194 246218
rect 535874 245898 535916 246134
rect 536152 245898 536194 246134
rect 535874 245866 536194 245898
rect 541805 246454 542125 246486
rect 541805 246218 541847 246454
rect 542083 246218 542125 246454
rect 541805 246134 542125 246218
rect 541805 245898 541847 246134
rect 542083 245898 542125 246134
rect 541805 245866 542125 245898
rect 19910 237454 20230 237486
rect 19910 237218 19952 237454
rect 20188 237218 20230 237454
rect 19910 237134 20230 237218
rect 19910 236898 19952 237134
rect 20188 236898 20230 237134
rect 19910 236866 20230 236898
rect 25840 237454 26160 237486
rect 25840 237218 25882 237454
rect 26118 237218 26160 237454
rect 25840 237134 26160 237218
rect 25840 236898 25882 237134
rect 26118 236898 26160 237134
rect 25840 236866 26160 236898
rect 31771 237454 32091 237486
rect 31771 237218 31813 237454
rect 32049 237218 32091 237454
rect 31771 237134 32091 237218
rect 31771 236898 31813 237134
rect 32049 236898 32091 237134
rect 31771 236866 32091 236898
rect 46910 237454 47230 237486
rect 46910 237218 46952 237454
rect 47188 237218 47230 237454
rect 46910 237134 47230 237218
rect 46910 236898 46952 237134
rect 47188 236898 47230 237134
rect 46910 236866 47230 236898
rect 52840 237454 53160 237486
rect 52840 237218 52882 237454
rect 53118 237218 53160 237454
rect 52840 237134 53160 237218
rect 52840 236898 52882 237134
rect 53118 236898 53160 237134
rect 52840 236866 53160 236898
rect 58771 237454 59091 237486
rect 58771 237218 58813 237454
rect 59049 237218 59091 237454
rect 58771 237134 59091 237218
rect 58771 236898 58813 237134
rect 59049 236898 59091 237134
rect 58771 236866 59091 236898
rect 73910 237454 74230 237486
rect 73910 237218 73952 237454
rect 74188 237218 74230 237454
rect 73910 237134 74230 237218
rect 73910 236898 73952 237134
rect 74188 236898 74230 237134
rect 73910 236866 74230 236898
rect 79840 237454 80160 237486
rect 79840 237218 79882 237454
rect 80118 237218 80160 237454
rect 79840 237134 80160 237218
rect 79840 236898 79882 237134
rect 80118 236898 80160 237134
rect 79840 236866 80160 236898
rect 85771 237454 86091 237486
rect 85771 237218 85813 237454
rect 86049 237218 86091 237454
rect 85771 237134 86091 237218
rect 85771 236898 85813 237134
rect 86049 236898 86091 237134
rect 85771 236866 86091 236898
rect 100910 237454 101230 237486
rect 100910 237218 100952 237454
rect 101188 237218 101230 237454
rect 100910 237134 101230 237218
rect 100910 236898 100952 237134
rect 101188 236898 101230 237134
rect 100910 236866 101230 236898
rect 106840 237454 107160 237486
rect 106840 237218 106882 237454
rect 107118 237218 107160 237454
rect 106840 237134 107160 237218
rect 106840 236898 106882 237134
rect 107118 236898 107160 237134
rect 106840 236866 107160 236898
rect 112771 237454 113091 237486
rect 112771 237218 112813 237454
rect 113049 237218 113091 237454
rect 112771 237134 113091 237218
rect 112771 236898 112813 237134
rect 113049 236898 113091 237134
rect 112771 236866 113091 236898
rect 127910 237454 128230 237486
rect 127910 237218 127952 237454
rect 128188 237218 128230 237454
rect 127910 237134 128230 237218
rect 127910 236898 127952 237134
rect 128188 236898 128230 237134
rect 127910 236866 128230 236898
rect 133840 237454 134160 237486
rect 133840 237218 133882 237454
rect 134118 237218 134160 237454
rect 133840 237134 134160 237218
rect 133840 236898 133882 237134
rect 134118 236898 134160 237134
rect 133840 236866 134160 236898
rect 139771 237454 140091 237486
rect 139771 237218 139813 237454
rect 140049 237218 140091 237454
rect 139771 237134 140091 237218
rect 139771 236898 139813 237134
rect 140049 236898 140091 237134
rect 139771 236866 140091 236898
rect 154910 237454 155230 237486
rect 154910 237218 154952 237454
rect 155188 237218 155230 237454
rect 154910 237134 155230 237218
rect 154910 236898 154952 237134
rect 155188 236898 155230 237134
rect 154910 236866 155230 236898
rect 160840 237454 161160 237486
rect 160840 237218 160882 237454
rect 161118 237218 161160 237454
rect 160840 237134 161160 237218
rect 160840 236898 160882 237134
rect 161118 236898 161160 237134
rect 160840 236866 161160 236898
rect 166771 237454 167091 237486
rect 166771 237218 166813 237454
rect 167049 237218 167091 237454
rect 166771 237134 167091 237218
rect 166771 236898 166813 237134
rect 167049 236898 167091 237134
rect 166771 236866 167091 236898
rect 181910 237454 182230 237486
rect 181910 237218 181952 237454
rect 182188 237218 182230 237454
rect 181910 237134 182230 237218
rect 181910 236898 181952 237134
rect 182188 236898 182230 237134
rect 181910 236866 182230 236898
rect 187840 237454 188160 237486
rect 187840 237218 187882 237454
rect 188118 237218 188160 237454
rect 187840 237134 188160 237218
rect 187840 236898 187882 237134
rect 188118 236898 188160 237134
rect 187840 236866 188160 236898
rect 193771 237454 194091 237486
rect 193771 237218 193813 237454
rect 194049 237218 194091 237454
rect 193771 237134 194091 237218
rect 193771 236898 193813 237134
rect 194049 236898 194091 237134
rect 193771 236866 194091 236898
rect 208910 237454 209230 237486
rect 208910 237218 208952 237454
rect 209188 237218 209230 237454
rect 208910 237134 209230 237218
rect 208910 236898 208952 237134
rect 209188 236898 209230 237134
rect 208910 236866 209230 236898
rect 214840 237454 215160 237486
rect 214840 237218 214882 237454
rect 215118 237218 215160 237454
rect 214840 237134 215160 237218
rect 214840 236898 214882 237134
rect 215118 236898 215160 237134
rect 214840 236866 215160 236898
rect 220771 237454 221091 237486
rect 220771 237218 220813 237454
rect 221049 237218 221091 237454
rect 220771 237134 221091 237218
rect 220771 236898 220813 237134
rect 221049 236898 221091 237134
rect 220771 236866 221091 236898
rect 235910 237454 236230 237486
rect 235910 237218 235952 237454
rect 236188 237218 236230 237454
rect 235910 237134 236230 237218
rect 235910 236898 235952 237134
rect 236188 236898 236230 237134
rect 235910 236866 236230 236898
rect 241840 237454 242160 237486
rect 241840 237218 241882 237454
rect 242118 237218 242160 237454
rect 241840 237134 242160 237218
rect 241840 236898 241882 237134
rect 242118 236898 242160 237134
rect 241840 236866 242160 236898
rect 247771 237454 248091 237486
rect 247771 237218 247813 237454
rect 248049 237218 248091 237454
rect 247771 237134 248091 237218
rect 247771 236898 247813 237134
rect 248049 236898 248091 237134
rect 247771 236866 248091 236898
rect 262910 237454 263230 237486
rect 262910 237218 262952 237454
rect 263188 237218 263230 237454
rect 262910 237134 263230 237218
rect 262910 236898 262952 237134
rect 263188 236898 263230 237134
rect 262910 236866 263230 236898
rect 268840 237454 269160 237486
rect 268840 237218 268882 237454
rect 269118 237218 269160 237454
rect 268840 237134 269160 237218
rect 268840 236898 268882 237134
rect 269118 236898 269160 237134
rect 268840 236866 269160 236898
rect 274771 237454 275091 237486
rect 274771 237218 274813 237454
rect 275049 237218 275091 237454
rect 274771 237134 275091 237218
rect 274771 236898 274813 237134
rect 275049 236898 275091 237134
rect 274771 236866 275091 236898
rect 289910 237454 290230 237486
rect 289910 237218 289952 237454
rect 290188 237218 290230 237454
rect 289910 237134 290230 237218
rect 289910 236898 289952 237134
rect 290188 236898 290230 237134
rect 289910 236866 290230 236898
rect 295840 237454 296160 237486
rect 295840 237218 295882 237454
rect 296118 237218 296160 237454
rect 295840 237134 296160 237218
rect 295840 236898 295882 237134
rect 296118 236898 296160 237134
rect 295840 236866 296160 236898
rect 301771 237454 302091 237486
rect 301771 237218 301813 237454
rect 302049 237218 302091 237454
rect 301771 237134 302091 237218
rect 301771 236898 301813 237134
rect 302049 236898 302091 237134
rect 301771 236866 302091 236898
rect 316910 237454 317230 237486
rect 316910 237218 316952 237454
rect 317188 237218 317230 237454
rect 316910 237134 317230 237218
rect 316910 236898 316952 237134
rect 317188 236898 317230 237134
rect 316910 236866 317230 236898
rect 322840 237454 323160 237486
rect 322840 237218 322882 237454
rect 323118 237218 323160 237454
rect 322840 237134 323160 237218
rect 322840 236898 322882 237134
rect 323118 236898 323160 237134
rect 322840 236866 323160 236898
rect 328771 237454 329091 237486
rect 328771 237218 328813 237454
rect 329049 237218 329091 237454
rect 328771 237134 329091 237218
rect 328771 236898 328813 237134
rect 329049 236898 329091 237134
rect 328771 236866 329091 236898
rect 343910 237454 344230 237486
rect 343910 237218 343952 237454
rect 344188 237218 344230 237454
rect 343910 237134 344230 237218
rect 343910 236898 343952 237134
rect 344188 236898 344230 237134
rect 343910 236866 344230 236898
rect 349840 237454 350160 237486
rect 349840 237218 349882 237454
rect 350118 237218 350160 237454
rect 349840 237134 350160 237218
rect 349840 236898 349882 237134
rect 350118 236898 350160 237134
rect 349840 236866 350160 236898
rect 355771 237454 356091 237486
rect 355771 237218 355813 237454
rect 356049 237218 356091 237454
rect 355771 237134 356091 237218
rect 355771 236898 355813 237134
rect 356049 236898 356091 237134
rect 355771 236866 356091 236898
rect 370910 237454 371230 237486
rect 370910 237218 370952 237454
rect 371188 237218 371230 237454
rect 370910 237134 371230 237218
rect 370910 236898 370952 237134
rect 371188 236898 371230 237134
rect 370910 236866 371230 236898
rect 376840 237454 377160 237486
rect 376840 237218 376882 237454
rect 377118 237218 377160 237454
rect 376840 237134 377160 237218
rect 376840 236898 376882 237134
rect 377118 236898 377160 237134
rect 376840 236866 377160 236898
rect 382771 237454 383091 237486
rect 382771 237218 382813 237454
rect 383049 237218 383091 237454
rect 382771 237134 383091 237218
rect 382771 236898 382813 237134
rect 383049 236898 383091 237134
rect 382771 236866 383091 236898
rect 397910 237454 398230 237486
rect 397910 237218 397952 237454
rect 398188 237218 398230 237454
rect 397910 237134 398230 237218
rect 397910 236898 397952 237134
rect 398188 236898 398230 237134
rect 397910 236866 398230 236898
rect 403840 237454 404160 237486
rect 403840 237218 403882 237454
rect 404118 237218 404160 237454
rect 403840 237134 404160 237218
rect 403840 236898 403882 237134
rect 404118 236898 404160 237134
rect 403840 236866 404160 236898
rect 409771 237454 410091 237486
rect 409771 237218 409813 237454
rect 410049 237218 410091 237454
rect 409771 237134 410091 237218
rect 409771 236898 409813 237134
rect 410049 236898 410091 237134
rect 409771 236866 410091 236898
rect 424910 237454 425230 237486
rect 424910 237218 424952 237454
rect 425188 237218 425230 237454
rect 424910 237134 425230 237218
rect 424910 236898 424952 237134
rect 425188 236898 425230 237134
rect 424910 236866 425230 236898
rect 430840 237454 431160 237486
rect 430840 237218 430882 237454
rect 431118 237218 431160 237454
rect 430840 237134 431160 237218
rect 430840 236898 430882 237134
rect 431118 236898 431160 237134
rect 430840 236866 431160 236898
rect 436771 237454 437091 237486
rect 436771 237218 436813 237454
rect 437049 237218 437091 237454
rect 436771 237134 437091 237218
rect 436771 236898 436813 237134
rect 437049 236898 437091 237134
rect 436771 236866 437091 236898
rect 451910 237454 452230 237486
rect 451910 237218 451952 237454
rect 452188 237218 452230 237454
rect 451910 237134 452230 237218
rect 451910 236898 451952 237134
rect 452188 236898 452230 237134
rect 451910 236866 452230 236898
rect 457840 237454 458160 237486
rect 457840 237218 457882 237454
rect 458118 237218 458160 237454
rect 457840 237134 458160 237218
rect 457840 236898 457882 237134
rect 458118 236898 458160 237134
rect 457840 236866 458160 236898
rect 463771 237454 464091 237486
rect 463771 237218 463813 237454
rect 464049 237218 464091 237454
rect 463771 237134 464091 237218
rect 463771 236898 463813 237134
rect 464049 236898 464091 237134
rect 463771 236866 464091 236898
rect 478910 237454 479230 237486
rect 478910 237218 478952 237454
rect 479188 237218 479230 237454
rect 478910 237134 479230 237218
rect 478910 236898 478952 237134
rect 479188 236898 479230 237134
rect 478910 236866 479230 236898
rect 484840 237454 485160 237486
rect 484840 237218 484882 237454
rect 485118 237218 485160 237454
rect 484840 237134 485160 237218
rect 484840 236898 484882 237134
rect 485118 236898 485160 237134
rect 484840 236866 485160 236898
rect 490771 237454 491091 237486
rect 490771 237218 490813 237454
rect 491049 237218 491091 237454
rect 490771 237134 491091 237218
rect 490771 236898 490813 237134
rect 491049 236898 491091 237134
rect 490771 236866 491091 236898
rect 505910 237454 506230 237486
rect 505910 237218 505952 237454
rect 506188 237218 506230 237454
rect 505910 237134 506230 237218
rect 505910 236898 505952 237134
rect 506188 236898 506230 237134
rect 505910 236866 506230 236898
rect 511840 237454 512160 237486
rect 511840 237218 511882 237454
rect 512118 237218 512160 237454
rect 511840 237134 512160 237218
rect 511840 236898 511882 237134
rect 512118 236898 512160 237134
rect 511840 236866 512160 236898
rect 517771 237454 518091 237486
rect 517771 237218 517813 237454
rect 518049 237218 518091 237454
rect 517771 237134 518091 237218
rect 517771 236898 517813 237134
rect 518049 236898 518091 237134
rect 517771 236866 518091 236898
rect 532910 237454 533230 237486
rect 532910 237218 532952 237454
rect 533188 237218 533230 237454
rect 532910 237134 533230 237218
rect 532910 236898 532952 237134
rect 533188 236898 533230 237134
rect 532910 236866 533230 236898
rect 538840 237454 539160 237486
rect 538840 237218 538882 237454
rect 539118 237218 539160 237454
rect 538840 237134 539160 237218
rect 538840 236898 538882 237134
rect 539118 236898 539160 237134
rect 538840 236866 539160 236898
rect 544771 237454 545091 237486
rect 544771 237218 544813 237454
rect 545049 237218 545091 237454
rect 544771 237134 545091 237218
rect 544771 236898 544813 237134
rect 545049 236898 545091 237134
rect 544771 236866 545091 236898
rect 559794 237454 560414 254898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 210454 11414 227898
rect 19794 229394 20414 230000
rect 19794 229158 19826 229394
rect 20062 229158 20146 229394
rect 20382 229158 20414 229394
rect 19794 229074 20414 229158
rect 19794 228838 19826 229074
rect 20062 228838 20146 229074
rect 20382 228838 20414 229074
rect 19794 227000 20414 228838
rect 28794 228454 29414 230000
rect 28794 228218 28826 228454
rect 29062 228218 29146 228454
rect 29382 228218 29414 228454
rect 28794 228134 29414 228218
rect 28794 227898 28826 228134
rect 29062 227898 29146 228134
rect 29382 227898 29414 228134
rect 28794 227000 29414 227898
rect 37794 229394 38414 230000
rect 37794 229158 37826 229394
rect 38062 229158 38146 229394
rect 38382 229158 38414 229394
rect 37794 229074 38414 229158
rect 37794 228838 37826 229074
rect 38062 228838 38146 229074
rect 38382 228838 38414 229074
rect 37794 227000 38414 228838
rect 46794 228454 47414 230000
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 227000 47414 227898
rect 55794 229394 56414 230000
rect 55794 229158 55826 229394
rect 56062 229158 56146 229394
rect 56382 229158 56414 229394
rect 55794 229074 56414 229158
rect 55794 228838 55826 229074
rect 56062 228838 56146 229074
rect 56382 228838 56414 229074
rect 55794 227000 56414 228838
rect 64794 228454 65414 230000
rect 64794 228218 64826 228454
rect 65062 228218 65146 228454
rect 65382 228218 65414 228454
rect 64794 228134 65414 228218
rect 64794 227898 64826 228134
rect 65062 227898 65146 228134
rect 65382 227898 65414 228134
rect 64794 227000 65414 227898
rect 73794 229394 74414 230000
rect 73794 229158 73826 229394
rect 74062 229158 74146 229394
rect 74382 229158 74414 229394
rect 73794 229074 74414 229158
rect 73794 228838 73826 229074
rect 74062 228838 74146 229074
rect 74382 228838 74414 229074
rect 73794 227000 74414 228838
rect 82794 228454 83414 230000
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 227000 83414 227898
rect 91794 229394 92414 230000
rect 91794 229158 91826 229394
rect 92062 229158 92146 229394
rect 92382 229158 92414 229394
rect 91794 229074 92414 229158
rect 91794 228838 91826 229074
rect 92062 228838 92146 229074
rect 92382 228838 92414 229074
rect 91794 227000 92414 228838
rect 100794 228454 101414 230000
rect 100794 228218 100826 228454
rect 101062 228218 101146 228454
rect 101382 228218 101414 228454
rect 100794 228134 101414 228218
rect 100794 227898 100826 228134
rect 101062 227898 101146 228134
rect 101382 227898 101414 228134
rect 100794 227000 101414 227898
rect 109794 229394 110414 230000
rect 109794 229158 109826 229394
rect 110062 229158 110146 229394
rect 110382 229158 110414 229394
rect 109794 229074 110414 229158
rect 109794 228838 109826 229074
rect 110062 228838 110146 229074
rect 110382 228838 110414 229074
rect 109794 227000 110414 228838
rect 118794 228454 119414 230000
rect 118794 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 119414 228454
rect 118794 228134 119414 228218
rect 118794 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 119414 228134
rect 118794 227000 119414 227898
rect 127794 229394 128414 230000
rect 127794 229158 127826 229394
rect 128062 229158 128146 229394
rect 128382 229158 128414 229394
rect 127794 229074 128414 229158
rect 127794 228838 127826 229074
rect 128062 228838 128146 229074
rect 128382 228838 128414 229074
rect 127794 227000 128414 228838
rect 136794 228454 137414 230000
rect 136794 228218 136826 228454
rect 137062 228218 137146 228454
rect 137382 228218 137414 228454
rect 136794 228134 137414 228218
rect 136794 227898 136826 228134
rect 137062 227898 137146 228134
rect 137382 227898 137414 228134
rect 136794 227000 137414 227898
rect 145794 229394 146414 230000
rect 145794 229158 145826 229394
rect 146062 229158 146146 229394
rect 146382 229158 146414 229394
rect 145794 229074 146414 229158
rect 145794 228838 145826 229074
rect 146062 228838 146146 229074
rect 146382 228838 146414 229074
rect 145794 227000 146414 228838
rect 154794 228454 155414 230000
rect 154794 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 155414 228454
rect 154794 228134 155414 228218
rect 154794 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 155414 228134
rect 154794 227000 155414 227898
rect 163794 229394 164414 230000
rect 163794 229158 163826 229394
rect 164062 229158 164146 229394
rect 164382 229158 164414 229394
rect 163794 229074 164414 229158
rect 163794 228838 163826 229074
rect 164062 228838 164146 229074
rect 164382 228838 164414 229074
rect 163794 227000 164414 228838
rect 172794 228454 173414 230000
rect 172794 228218 172826 228454
rect 173062 228218 173146 228454
rect 173382 228218 173414 228454
rect 172794 228134 173414 228218
rect 172794 227898 172826 228134
rect 173062 227898 173146 228134
rect 173382 227898 173414 228134
rect 172794 227000 173414 227898
rect 181794 229394 182414 230000
rect 181794 229158 181826 229394
rect 182062 229158 182146 229394
rect 182382 229158 182414 229394
rect 181794 229074 182414 229158
rect 181794 228838 181826 229074
rect 182062 228838 182146 229074
rect 182382 228838 182414 229074
rect 181794 227000 182414 228838
rect 190794 228454 191414 230000
rect 190794 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 191414 228454
rect 190794 228134 191414 228218
rect 190794 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 191414 228134
rect 190794 227000 191414 227898
rect 199794 229394 200414 230000
rect 199794 229158 199826 229394
rect 200062 229158 200146 229394
rect 200382 229158 200414 229394
rect 199794 229074 200414 229158
rect 199794 228838 199826 229074
rect 200062 228838 200146 229074
rect 200382 228838 200414 229074
rect 199794 227000 200414 228838
rect 208794 228454 209414 230000
rect 208794 228218 208826 228454
rect 209062 228218 209146 228454
rect 209382 228218 209414 228454
rect 208794 228134 209414 228218
rect 208794 227898 208826 228134
rect 209062 227898 209146 228134
rect 209382 227898 209414 228134
rect 208794 227000 209414 227898
rect 217794 229394 218414 230000
rect 217794 229158 217826 229394
rect 218062 229158 218146 229394
rect 218382 229158 218414 229394
rect 217794 229074 218414 229158
rect 217794 228838 217826 229074
rect 218062 228838 218146 229074
rect 218382 228838 218414 229074
rect 217794 227000 218414 228838
rect 226794 228454 227414 230000
rect 226794 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 227414 228454
rect 226794 228134 227414 228218
rect 226794 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 227414 228134
rect 226794 227000 227414 227898
rect 235794 229394 236414 230000
rect 235794 229158 235826 229394
rect 236062 229158 236146 229394
rect 236382 229158 236414 229394
rect 235794 229074 236414 229158
rect 235794 228838 235826 229074
rect 236062 228838 236146 229074
rect 236382 228838 236414 229074
rect 235794 227000 236414 228838
rect 244794 228454 245414 230000
rect 244794 228218 244826 228454
rect 245062 228218 245146 228454
rect 245382 228218 245414 228454
rect 244794 228134 245414 228218
rect 244794 227898 244826 228134
rect 245062 227898 245146 228134
rect 245382 227898 245414 228134
rect 244794 227000 245414 227898
rect 253794 229394 254414 230000
rect 253794 229158 253826 229394
rect 254062 229158 254146 229394
rect 254382 229158 254414 229394
rect 253794 229074 254414 229158
rect 253794 228838 253826 229074
rect 254062 228838 254146 229074
rect 254382 228838 254414 229074
rect 253794 227000 254414 228838
rect 262794 228454 263414 230000
rect 262794 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 263414 228454
rect 262794 228134 263414 228218
rect 262794 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 263414 228134
rect 262794 227000 263414 227898
rect 271794 229394 272414 230000
rect 271794 229158 271826 229394
rect 272062 229158 272146 229394
rect 272382 229158 272414 229394
rect 271794 229074 272414 229158
rect 271794 228838 271826 229074
rect 272062 228838 272146 229074
rect 272382 228838 272414 229074
rect 271794 227000 272414 228838
rect 280794 228454 281414 230000
rect 280794 228218 280826 228454
rect 281062 228218 281146 228454
rect 281382 228218 281414 228454
rect 280794 228134 281414 228218
rect 280794 227898 280826 228134
rect 281062 227898 281146 228134
rect 281382 227898 281414 228134
rect 280794 227000 281414 227898
rect 289794 229394 290414 230000
rect 289794 229158 289826 229394
rect 290062 229158 290146 229394
rect 290382 229158 290414 229394
rect 289794 229074 290414 229158
rect 289794 228838 289826 229074
rect 290062 228838 290146 229074
rect 290382 228838 290414 229074
rect 289794 227000 290414 228838
rect 298794 228454 299414 230000
rect 298794 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 299414 228454
rect 298794 228134 299414 228218
rect 298794 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 299414 228134
rect 298794 227000 299414 227898
rect 307794 229394 308414 230000
rect 307794 229158 307826 229394
rect 308062 229158 308146 229394
rect 308382 229158 308414 229394
rect 307794 229074 308414 229158
rect 307794 228838 307826 229074
rect 308062 228838 308146 229074
rect 308382 228838 308414 229074
rect 307794 227000 308414 228838
rect 316794 228454 317414 230000
rect 316794 228218 316826 228454
rect 317062 228218 317146 228454
rect 317382 228218 317414 228454
rect 316794 228134 317414 228218
rect 316794 227898 316826 228134
rect 317062 227898 317146 228134
rect 317382 227898 317414 228134
rect 316794 227000 317414 227898
rect 325794 229394 326414 230000
rect 325794 229158 325826 229394
rect 326062 229158 326146 229394
rect 326382 229158 326414 229394
rect 325794 229074 326414 229158
rect 325794 228838 325826 229074
rect 326062 228838 326146 229074
rect 326382 228838 326414 229074
rect 325794 227000 326414 228838
rect 334794 228454 335414 230000
rect 334794 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 335414 228454
rect 334794 228134 335414 228218
rect 334794 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 335414 228134
rect 334794 227000 335414 227898
rect 343794 229394 344414 230000
rect 343794 229158 343826 229394
rect 344062 229158 344146 229394
rect 344382 229158 344414 229394
rect 343794 229074 344414 229158
rect 343794 228838 343826 229074
rect 344062 228838 344146 229074
rect 344382 228838 344414 229074
rect 343794 227000 344414 228838
rect 352794 228454 353414 230000
rect 352794 228218 352826 228454
rect 353062 228218 353146 228454
rect 353382 228218 353414 228454
rect 352794 228134 353414 228218
rect 352794 227898 352826 228134
rect 353062 227898 353146 228134
rect 353382 227898 353414 228134
rect 352794 227000 353414 227898
rect 361794 229394 362414 230000
rect 361794 229158 361826 229394
rect 362062 229158 362146 229394
rect 362382 229158 362414 229394
rect 361794 229074 362414 229158
rect 361794 228838 361826 229074
rect 362062 228838 362146 229074
rect 362382 228838 362414 229074
rect 361794 227000 362414 228838
rect 370794 228454 371414 230000
rect 370794 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 371414 228454
rect 370794 228134 371414 228218
rect 370794 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 371414 228134
rect 370794 227000 371414 227898
rect 379794 229394 380414 230000
rect 379794 229158 379826 229394
rect 380062 229158 380146 229394
rect 380382 229158 380414 229394
rect 379794 229074 380414 229158
rect 379794 228838 379826 229074
rect 380062 228838 380146 229074
rect 380382 228838 380414 229074
rect 379794 227000 380414 228838
rect 388794 228454 389414 230000
rect 388794 228218 388826 228454
rect 389062 228218 389146 228454
rect 389382 228218 389414 228454
rect 388794 228134 389414 228218
rect 388794 227898 388826 228134
rect 389062 227898 389146 228134
rect 389382 227898 389414 228134
rect 388794 227000 389414 227898
rect 397794 229394 398414 230000
rect 397794 229158 397826 229394
rect 398062 229158 398146 229394
rect 398382 229158 398414 229394
rect 397794 229074 398414 229158
rect 397794 228838 397826 229074
rect 398062 228838 398146 229074
rect 398382 228838 398414 229074
rect 397794 227000 398414 228838
rect 406794 228454 407414 230000
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 227000 407414 227898
rect 415794 229394 416414 230000
rect 415794 229158 415826 229394
rect 416062 229158 416146 229394
rect 416382 229158 416414 229394
rect 415794 229074 416414 229158
rect 415794 228838 415826 229074
rect 416062 228838 416146 229074
rect 416382 228838 416414 229074
rect 415794 227000 416414 228838
rect 424794 228454 425414 230000
rect 424794 228218 424826 228454
rect 425062 228218 425146 228454
rect 425382 228218 425414 228454
rect 424794 228134 425414 228218
rect 424794 227898 424826 228134
rect 425062 227898 425146 228134
rect 425382 227898 425414 228134
rect 424794 227000 425414 227898
rect 433794 229394 434414 230000
rect 433794 229158 433826 229394
rect 434062 229158 434146 229394
rect 434382 229158 434414 229394
rect 433794 229074 434414 229158
rect 433794 228838 433826 229074
rect 434062 228838 434146 229074
rect 434382 228838 434414 229074
rect 433794 227000 434414 228838
rect 442794 228454 443414 230000
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 227000 443414 227898
rect 451794 229394 452414 230000
rect 451794 229158 451826 229394
rect 452062 229158 452146 229394
rect 452382 229158 452414 229394
rect 451794 229074 452414 229158
rect 451794 228838 451826 229074
rect 452062 228838 452146 229074
rect 452382 228838 452414 229074
rect 451794 227000 452414 228838
rect 460794 228454 461414 230000
rect 460794 228218 460826 228454
rect 461062 228218 461146 228454
rect 461382 228218 461414 228454
rect 460794 228134 461414 228218
rect 460794 227898 460826 228134
rect 461062 227898 461146 228134
rect 461382 227898 461414 228134
rect 460794 227000 461414 227898
rect 469794 229394 470414 230000
rect 469794 229158 469826 229394
rect 470062 229158 470146 229394
rect 470382 229158 470414 229394
rect 469794 229074 470414 229158
rect 469794 228838 469826 229074
rect 470062 228838 470146 229074
rect 470382 228838 470414 229074
rect 469794 227000 470414 228838
rect 478794 228454 479414 230000
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 227000 479414 227898
rect 487794 229394 488414 230000
rect 487794 229158 487826 229394
rect 488062 229158 488146 229394
rect 488382 229158 488414 229394
rect 487794 229074 488414 229158
rect 487794 228838 487826 229074
rect 488062 228838 488146 229074
rect 488382 228838 488414 229074
rect 487794 227000 488414 228838
rect 496794 228454 497414 230000
rect 496794 228218 496826 228454
rect 497062 228218 497146 228454
rect 497382 228218 497414 228454
rect 496794 228134 497414 228218
rect 496794 227898 496826 228134
rect 497062 227898 497146 228134
rect 497382 227898 497414 228134
rect 496794 227000 497414 227898
rect 505794 229394 506414 230000
rect 505794 229158 505826 229394
rect 506062 229158 506146 229394
rect 506382 229158 506414 229394
rect 505794 229074 506414 229158
rect 505794 228838 505826 229074
rect 506062 228838 506146 229074
rect 506382 228838 506414 229074
rect 505794 227000 506414 228838
rect 514794 228454 515414 230000
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 227000 515414 227898
rect 523794 229394 524414 230000
rect 523794 229158 523826 229394
rect 524062 229158 524146 229394
rect 524382 229158 524414 229394
rect 523794 229074 524414 229158
rect 523794 228838 523826 229074
rect 524062 228838 524146 229074
rect 524382 228838 524414 229074
rect 523794 227000 524414 228838
rect 532794 228454 533414 230000
rect 532794 228218 532826 228454
rect 533062 228218 533146 228454
rect 533382 228218 533414 228454
rect 532794 228134 533414 228218
rect 532794 227898 532826 228134
rect 533062 227898 533146 228134
rect 533382 227898 533414 228134
rect 532794 227000 533414 227898
rect 541794 229394 542414 230000
rect 541794 229158 541826 229394
rect 542062 229158 542146 229394
rect 542382 229158 542414 229394
rect 541794 229074 542414 229158
rect 541794 228838 541826 229074
rect 542062 228838 542146 229074
rect 542382 228838 542414 229074
rect 541794 227000 542414 228838
rect 550794 228454 551414 230000
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 227000 551414 227898
rect 19910 219454 20230 219486
rect 19910 219218 19952 219454
rect 20188 219218 20230 219454
rect 19910 219134 20230 219218
rect 19910 218898 19952 219134
rect 20188 218898 20230 219134
rect 19910 218866 20230 218898
rect 25840 219454 26160 219486
rect 25840 219218 25882 219454
rect 26118 219218 26160 219454
rect 25840 219134 26160 219218
rect 25840 218898 25882 219134
rect 26118 218898 26160 219134
rect 25840 218866 26160 218898
rect 31771 219454 32091 219486
rect 31771 219218 31813 219454
rect 32049 219218 32091 219454
rect 31771 219134 32091 219218
rect 31771 218898 31813 219134
rect 32049 218898 32091 219134
rect 31771 218866 32091 218898
rect 46910 219454 47230 219486
rect 46910 219218 46952 219454
rect 47188 219218 47230 219454
rect 46910 219134 47230 219218
rect 46910 218898 46952 219134
rect 47188 218898 47230 219134
rect 46910 218866 47230 218898
rect 52840 219454 53160 219486
rect 52840 219218 52882 219454
rect 53118 219218 53160 219454
rect 52840 219134 53160 219218
rect 52840 218898 52882 219134
rect 53118 218898 53160 219134
rect 52840 218866 53160 218898
rect 58771 219454 59091 219486
rect 58771 219218 58813 219454
rect 59049 219218 59091 219454
rect 58771 219134 59091 219218
rect 58771 218898 58813 219134
rect 59049 218898 59091 219134
rect 58771 218866 59091 218898
rect 73910 219454 74230 219486
rect 73910 219218 73952 219454
rect 74188 219218 74230 219454
rect 73910 219134 74230 219218
rect 73910 218898 73952 219134
rect 74188 218898 74230 219134
rect 73910 218866 74230 218898
rect 79840 219454 80160 219486
rect 79840 219218 79882 219454
rect 80118 219218 80160 219454
rect 79840 219134 80160 219218
rect 79840 218898 79882 219134
rect 80118 218898 80160 219134
rect 79840 218866 80160 218898
rect 85771 219454 86091 219486
rect 85771 219218 85813 219454
rect 86049 219218 86091 219454
rect 85771 219134 86091 219218
rect 85771 218898 85813 219134
rect 86049 218898 86091 219134
rect 85771 218866 86091 218898
rect 100910 219454 101230 219486
rect 100910 219218 100952 219454
rect 101188 219218 101230 219454
rect 100910 219134 101230 219218
rect 100910 218898 100952 219134
rect 101188 218898 101230 219134
rect 100910 218866 101230 218898
rect 106840 219454 107160 219486
rect 106840 219218 106882 219454
rect 107118 219218 107160 219454
rect 106840 219134 107160 219218
rect 106840 218898 106882 219134
rect 107118 218898 107160 219134
rect 106840 218866 107160 218898
rect 112771 219454 113091 219486
rect 112771 219218 112813 219454
rect 113049 219218 113091 219454
rect 112771 219134 113091 219218
rect 112771 218898 112813 219134
rect 113049 218898 113091 219134
rect 112771 218866 113091 218898
rect 127910 219454 128230 219486
rect 127910 219218 127952 219454
rect 128188 219218 128230 219454
rect 127910 219134 128230 219218
rect 127910 218898 127952 219134
rect 128188 218898 128230 219134
rect 127910 218866 128230 218898
rect 133840 219454 134160 219486
rect 133840 219218 133882 219454
rect 134118 219218 134160 219454
rect 133840 219134 134160 219218
rect 133840 218898 133882 219134
rect 134118 218898 134160 219134
rect 133840 218866 134160 218898
rect 139771 219454 140091 219486
rect 139771 219218 139813 219454
rect 140049 219218 140091 219454
rect 139771 219134 140091 219218
rect 139771 218898 139813 219134
rect 140049 218898 140091 219134
rect 139771 218866 140091 218898
rect 154910 219454 155230 219486
rect 154910 219218 154952 219454
rect 155188 219218 155230 219454
rect 154910 219134 155230 219218
rect 154910 218898 154952 219134
rect 155188 218898 155230 219134
rect 154910 218866 155230 218898
rect 160840 219454 161160 219486
rect 160840 219218 160882 219454
rect 161118 219218 161160 219454
rect 160840 219134 161160 219218
rect 160840 218898 160882 219134
rect 161118 218898 161160 219134
rect 160840 218866 161160 218898
rect 166771 219454 167091 219486
rect 166771 219218 166813 219454
rect 167049 219218 167091 219454
rect 166771 219134 167091 219218
rect 166771 218898 166813 219134
rect 167049 218898 167091 219134
rect 166771 218866 167091 218898
rect 181910 219454 182230 219486
rect 181910 219218 181952 219454
rect 182188 219218 182230 219454
rect 181910 219134 182230 219218
rect 181910 218898 181952 219134
rect 182188 218898 182230 219134
rect 181910 218866 182230 218898
rect 187840 219454 188160 219486
rect 187840 219218 187882 219454
rect 188118 219218 188160 219454
rect 187840 219134 188160 219218
rect 187840 218898 187882 219134
rect 188118 218898 188160 219134
rect 187840 218866 188160 218898
rect 193771 219454 194091 219486
rect 193771 219218 193813 219454
rect 194049 219218 194091 219454
rect 193771 219134 194091 219218
rect 193771 218898 193813 219134
rect 194049 218898 194091 219134
rect 193771 218866 194091 218898
rect 208910 219454 209230 219486
rect 208910 219218 208952 219454
rect 209188 219218 209230 219454
rect 208910 219134 209230 219218
rect 208910 218898 208952 219134
rect 209188 218898 209230 219134
rect 208910 218866 209230 218898
rect 214840 219454 215160 219486
rect 214840 219218 214882 219454
rect 215118 219218 215160 219454
rect 214840 219134 215160 219218
rect 214840 218898 214882 219134
rect 215118 218898 215160 219134
rect 214840 218866 215160 218898
rect 220771 219454 221091 219486
rect 220771 219218 220813 219454
rect 221049 219218 221091 219454
rect 220771 219134 221091 219218
rect 220771 218898 220813 219134
rect 221049 218898 221091 219134
rect 220771 218866 221091 218898
rect 235910 219454 236230 219486
rect 235910 219218 235952 219454
rect 236188 219218 236230 219454
rect 235910 219134 236230 219218
rect 235910 218898 235952 219134
rect 236188 218898 236230 219134
rect 235910 218866 236230 218898
rect 241840 219454 242160 219486
rect 241840 219218 241882 219454
rect 242118 219218 242160 219454
rect 241840 219134 242160 219218
rect 241840 218898 241882 219134
rect 242118 218898 242160 219134
rect 241840 218866 242160 218898
rect 247771 219454 248091 219486
rect 247771 219218 247813 219454
rect 248049 219218 248091 219454
rect 247771 219134 248091 219218
rect 247771 218898 247813 219134
rect 248049 218898 248091 219134
rect 247771 218866 248091 218898
rect 262910 219454 263230 219486
rect 262910 219218 262952 219454
rect 263188 219218 263230 219454
rect 262910 219134 263230 219218
rect 262910 218898 262952 219134
rect 263188 218898 263230 219134
rect 262910 218866 263230 218898
rect 268840 219454 269160 219486
rect 268840 219218 268882 219454
rect 269118 219218 269160 219454
rect 268840 219134 269160 219218
rect 268840 218898 268882 219134
rect 269118 218898 269160 219134
rect 268840 218866 269160 218898
rect 274771 219454 275091 219486
rect 274771 219218 274813 219454
rect 275049 219218 275091 219454
rect 274771 219134 275091 219218
rect 274771 218898 274813 219134
rect 275049 218898 275091 219134
rect 274771 218866 275091 218898
rect 289910 219454 290230 219486
rect 289910 219218 289952 219454
rect 290188 219218 290230 219454
rect 289910 219134 290230 219218
rect 289910 218898 289952 219134
rect 290188 218898 290230 219134
rect 289910 218866 290230 218898
rect 295840 219454 296160 219486
rect 295840 219218 295882 219454
rect 296118 219218 296160 219454
rect 295840 219134 296160 219218
rect 295840 218898 295882 219134
rect 296118 218898 296160 219134
rect 295840 218866 296160 218898
rect 301771 219454 302091 219486
rect 301771 219218 301813 219454
rect 302049 219218 302091 219454
rect 301771 219134 302091 219218
rect 301771 218898 301813 219134
rect 302049 218898 302091 219134
rect 301771 218866 302091 218898
rect 316910 219454 317230 219486
rect 316910 219218 316952 219454
rect 317188 219218 317230 219454
rect 316910 219134 317230 219218
rect 316910 218898 316952 219134
rect 317188 218898 317230 219134
rect 316910 218866 317230 218898
rect 322840 219454 323160 219486
rect 322840 219218 322882 219454
rect 323118 219218 323160 219454
rect 322840 219134 323160 219218
rect 322840 218898 322882 219134
rect 323118 218898 323160 219134
rect 322840 218866 323160 218898
rect 328771 219454 329091 219486
rect 328771 219218 328813 219454
rect 329049 219218 329091 219454
rect 328771 219134 329091 219218
rect 328771 218898 328813 219134
rect 329049 218898 329091 219134
rect 328771 218866 329091 218898
rect 343910 219454 344230 219486
rect 343910 219218 343952 219454
rect 344188 219218 344230 219454
rect 343910 219134 344230 219218
rect 343910 218898 343952 219134
rect 344188 218898 344230 219134
rect 343910 218866 344230 218898
rect 349840 219454 350160 219486
rect 349840 219218 349882 219454
rect 350118 219218 350160 219454
rect 349840 219134 350160 219218
rect 349840 218898 349882 219134
rect 350118 218898 350160 219134
rect 349840 218866 350160 218898
rect 355771 219454 356091 219486
rect 355771 219218 355813 219454
rect 356049 219218 356091 219454
rect 355771 219134 356091 219218
rect 355771 218898 355813 219134
rect 356049 218898 356091 219134
rect 355771 218866 356091 218898
rect 370910 219454 371230 219486
rect 370910 219218 370952 219454
rect 371188 219218 371230 219454
rect 370910 219134 371230 219218
rect 370910 218898 370952 219134
rect 371188 218898 371230 219134
rect 370910 218866 371230 218898
rect 376840 219454 377160 219486
rect 376840 219218 376882 219454
rect 377118 219218 377160 219454
rect 376840 219134 377160 219218
rect 376840 218898 376882 219134
rect 377118 218898 377160 219134
rect 376840 218866 377160 218898
rect 382771 219454 383091 219486
rect 382771 219218 382813 219454
rect 383049 219218 383091 219454
rect 382771 219134 383091 219218
rect 382771 218898 382813 219134
rect 383049 218898 383091 219134
rect 382771 218866 383091 218898
rect 397910 219454 398230 219486
rect 397910 219218 397952 219454
rect 398188 219218 398230 219454
rect 397910 219134 398230 219218
rect 397910 218898 397952 219134
rect 398188 218898 398230 219134
rect 397910 218866 398230 218898
rect 403840 219454 404160 219486
rect 403840 219218 403882 219454
rect 404118 219218 404160 219454
rect 403840 219134 404160 219218
rect 403840 218898 403882 219134
rect 404118 218898 404160 219134
rect 403840 218866 404160 218898
rect 409771 219454 410091 219486
rect 409771 219218 409813 219454
rect 410049 219218 410091 219454
rect 409771 219134 410091 219218
rect 409771 218898 409813 219134
rect 410049 218898 410091 219134
rect 409771 218866 410091 218898
rect 424910 219454 425230 219486
rect 424910 219218 424952 219454
rect 425188 219218 425230 219454
rect 424910 219134 425230 219218
rect 424910 218898 424952 219134
rect 425188 218898 425230 219134
rect 424910 218866 425230 218898
rect 430840 219454 431160 219486
rect 430840 219218 430882 219454
rect 431118 219218 431160 219454
rect 430840 219134 431160 219218
rect 430840 218898 430882 219134
rect 431118 218898 431160 219134
rect 430840 218866 431160 218898
rect 436771 219454 437091 219486
rect 436771 219218 436813 219454
rect 437049 219218 437091 219454
rect 436771 219134 437091 219218
rect 436771 218898 436813 219134
rect 437049 218898 437091 219134
rect 436771 218866 437091 218898
rect 451910 219454 452230 219486
rect 451910 219218 451952 219454
rect 452188 219218 452230 219454
rect 451910 219134 452230 219218
rect 451910 218898 451952 219134
rect 452188 218898 452230 219134
rect 451910 218866 452230 218898
rect 457840 219454 458160 219486
rect 457840 219218 457882 219454
rect 458118 219218 458160 219454
rect 457840 219134 458160 219218
rect 457840 218898 457882 219134
rect 458118 218898 458160 219134
rect 457840 218866 458160 218898
rect 463771 219454 464091 219486
rect 463771 219218 463813 219454
rect 464049 219218 464091 219454
rect 463771 219134 464091 219218
rect 463771 218898 463813 219134
rect 464049 218898 464091 219134
rect 463771 218866 464091 218898
rect 478910 219454 479230 219486
rect 478910 219218 478952 219454
rect 479188 219218 479230 219454
rect 478910 219134 479230 219218
rect 478910 218898 478952 219134
rect 479188 218898 479230 219134
rect 478910 218866 479230 218898
rect 484840 219454 485160 219486
rect 484840 219218 484882 219454
rect 485118 219218 485160 219454
rect 484840 219134 485160 219218
rect 484840 218898 484882 219134
rect 485118 218898 485160 219134
rect 484840 218866 485160 218898
rect 490771 219454 491091 219486
rect 490771 219218 490813 219454
rect 491049 219218 491091 219454
rect 490771 219134 491091 219218
rect 490771 218898 490813 219134
rect 491049 218898 491091 219134
rect 490771 218866 491091 218898
rect 505910 219454 506230 219486
rect 505910 219218 505952 219454
rect 506188 219218 506230 219454
rect 505910 219134 506230 219218
rect 505910 218898 505952 219134
rect 506188 218898 506230 219134
rect 505910 218866 506230 218898
rect 511840 219454 512160 219486
rect 511840 219218 511882 219454
rect 512118 219218 512160 219454
rect 511840 219134 512160 219218
rect 511840 218898 511882 219134
rect 512118 218898 512160 219134
rect 511840 218866 512160 218898
rect 517771 219454 518091 219486
rect 517771 219218 517813 219454
rect 518049 219218 518091 219454
rect 517771 219134 518091 219218
rect 517771 218898 517813 219134
rect 518049 218898 518091 219134
rect 517771 218866 518091 218898
rect 532910 219454 533230 219486
rect 532910 219218 532952 219454
rect 533188 219218 533230 219454
rect 532910 219134 533230 219218
rect 532910 218898 532952 219134
rect 533188 218898 533230 219134
rect 532910 218866 533230 218898
rect 538840 219454 539160 219486
rect 538840 219218 538882 219454
rect 539118 219218 539160 219454
rect 538840 219134 539160 219218
rect 538840 218898 538882 219134
rect 539118 218898 539160 219134
rect 538840 218866 539160 218898
rect 544771 219454 545091 219486
rect 544771 219218 544813 219454
rect 545049 219218 545091 219454
rect 544771 219134 545091 219218
rect 544771 218898 544813 219134
rect 545049 218898 545091 219134
rect 544771 218866 545091 218898
rect 559794 219454 560414 236898
rect 559794 219218 559826 219454
rect 560062 219218 560146 219454
rect 560382 219218 560414 219454
rect 559794 219134 560414 219218
rect 559794 218898 559826 219134
rect 560062 218898 560146 219134
rect 560382 218898 560414 219134
rect 10794 210218 10826 210454
rect 11062 210218 11146 210454
rect 11382 210218 11414 210454
rect 10794 210134 11414 210218
rect 10794 209898 10826 210134
rect 11062 209898 11146 210134
rect 11382 209898 11414 210134
rect 10794 192454 11414 209898
rect 22874 210454 23194 210486
rect 22874 210218 22916 210454
rect 23152 210218 23194 210454
rect 22874 210134 23194 210218
rect 22874 209898 22916 210134
rect 23152 209898 23194 210134
rect 22874 209866 23194 209898
rect 28805 210454 29125 210486
rect 28805 210218 28847 210454
rect 29083 210218 29125 210454
rect 28805 210134 29125 210218
rect 28805 209898 28847 210134
rect 29083 209898 29125 210134
rect 28805 209866 29125 209898
rect 49874 210454 50194 210486
rect 49874 210218 49916 210454
rect 50152 210218 50194 210454
rect 49874 210134 50194 210218
rect 49874 209898 49916 210134
rect 50152 209898 50194 210134
rect 49874 209866 50194 209898
rect 55805 210454 56125 210486
rect 55805 210218 55847 210454
rect 56083 210218 56125 210454
rect 55805 210134 56125 210218
rect 55805 209898 55847 210134
rect 56083 209898 56125 210134
rect 55805 209866 56125 209898
rect 76874 210454 77194 210486
rect 76874 210218 76916 210454
rect 77152 210218 77194 210454
rect 76874 210134 77194 210218
rect 76874 209898 76916 210134
rect 77152 209898 77194 210134
rect 76874 209866 77194 209898
rect 82805 210454 83125 210486
rect 82805 210218 82847 210454
rect 83083 210218 83125 210454
rect 82805 210134 83125 210218
rect 82805 209898 82847 210134
rect 83083 209898 83125 210134
rect 82805 209866 83125 209898
rect 103874 210454 104194 210486
rect 103874 210218 103916 210454
rect 104152 210218 104194 210454
rect 103874 210134 104194 210218
rect 103874 209898 103916 210134
rect 104152 209898 104194 210134
rect 103874 209866 104194 209898
rect 109805 210454 110125 210486
rect 109805 210218 109847 210454
rect 110083 210218 110125 210454
rect 109805 210134 110125 210218
rect 109805 209898 109847 210134
rect 110083 209898 110125 210134
rect 109805 209866 110125 209898
rect 130874 210454 131194 210486
rect 130874 210218 130916 210454
rect 131152 210218 131194 210454
rect 130874 210134 131194 210218
rect 130874 209898 130916 210134
rect 131152 209898 131194 210134
rect 130874 209866 131194 209898
rect 136805 210454 137125 210486
rect 136805 210218 136847 210454
rect 137083 210218 137125 210454
rect 136805 210134 137125 210218
rect 136805 209898 136847 210134
rect 137083 209898 137125 210134
rect 136805 209866 137125 209898
rect 157874 210454 158194 210486
rect 157874 210218 157916 210454
rect 158152 210218 158194 210454
rect 157874 210134 158194 210218
rect 157874 209898 157916 210134
rect 158152 209898 158194 210134
rect 157874 209866 158194 209898
rect 163805 210454 164125 210486
rect 163805 210218 163847 210454
rect 164083 210218 164125 210454
rect 163805 210134 164125 210218
rect 163805 209898 163847 210134
rect 164083 209898 164125 210134
rect 163805 209866 164125 209898
rect 184874 210454 185194 210486
rect 184874 210218 184916 210454
rect 185152 210218 185194 210454
rect 184874 210134 185194 210218
rect 184874 209898 184916 210134
rect 185152 209898 185194 210134
rect 184874 209866 185194 209898
rect 190805 210454 191125 210486
rect 190805 210218 190847 210454
rect 191083 210218 191125 210454
rect 190805 210134 191125 210218
rect 190805 209898 190847 210134
rect 191083 209898 191125 210134
rect 190805 209866 191125 209898
rect 211874 210454 212194 210486
rect 211874 210218 211916 210454
rect 212152 210218 212194 210454
rect 211874 210134 212194 210218
rect 211874 209898 211916 210134
rect 212152 209898 212194 210134
rect 211874 209866 212194 209898
rect 217805 210454 218125 210486
rect 217805 210218 217847 210454
rect 218083 210218 218125 210454
rect 217805 210134 218125 210218
rect 217805 209898 217847 210134
rect 218083 209898 218125 210134
rect 217805 209866 218125 209898
rect 238874 210454 239194 210486
rect 238874 210218 238916 210454
rect 239152 210218 239194 210454
rect 238874 210134 239194 210218
rect 238874 209898 238916 210134
rect 239152 209898 239194 210134
rect 238874 209866 239194 209898
rect 244805 210454 245125 210486
rect 244805 210218 244847 210454
rect 245083 210218 245125 210454
rect 244805 210134 245125 210218
rect 244805 209898 244847 210134
rect 245083 209898 245125 210134
rect 244805 209866 245125 209898
rect 265874 210454 266194 210486
rect 265874 210218 265916 210454
rect 266152 210218 266194 210454
rect 265874 210134 266194 210218
rect 265874 209898 265916 210134
rect 266152 209898 266194 210134
rect 265874 209866 266194 209898
rect 271805 210454 272125 210486
rect 271805 210218 271847 210454
rect 272083 210218 272125 210454
rect 271805 210134 272125 210218
rect 271805 209898 271847 210134
rect 272083 209898 272125 210134
rect 271805 209866 272125 209898
rect 292874 210454 293194 210486
rect 292874 210218 292916 210454
rect 293152 210218 293194 210454
rect 292874 210134 293194 210218
rect 292874 209898 292916 210134
rect 293152 209898 293194 210134
rect 292874 209866 293194 209898
rect 298805 210454 299125 210486
rect 298805 210218 298847 210454
rect 299083 210218 299125 210454
rect 298805 210134 299125 210218
rect 298805 209898 298847 210134
rect 299083 209898 299125 210134
rect 298805 209866 299125 209898
rect 319874 210454 320194 210486
rect 319874 210218 319916 210454
rect 320152 210218 320194 210454
rect 319874 210134 320194 210218
rect 319874 209898 319916 210134
rect 320152 209898 320194 210134
rect 319874 209866 320194 209898
rect 325805 210454 326125 210486
rect 325805 210218 325847 210454
rect 326083 210218 326125 210454
rect 325805 210134 326125 210218
rect 325805 209898 325847 210134
rect 326083 209898 326125 210134
rect 325805 209866 326125 209898
rect 346874 210454 347194 210486
rect 346874 210218 346916 210454
rect 347152 210218 347194 210454
rect 346874 210134 347194 210218
rect 346874 209898 346916 210134
rect 347152 209898 347194 210134
rect 346874 209866 347194 209898
rect 352805 210454 353125 210486
rect 352805 210218 352847 210454
rect 353083 210218 353125 210454
rect 352805 210134 353125 210218
rect 352805 209898 352847 210134
rect 353083 209898 353125 210134
rect 352805 209866 353125 209898
rect 373874 210454 374194 210486
rect 373874 210218 373916 210454
rect 374152 210218 374194 210454
rect 373874 210134 374194 210218
rect 373874 209898 373916 210134
rect 374152 209898 374194 210134
rect 373874 209866 374194 209898
rect 379805 210454 380125 210486
rect 379805 210218 379847 210454
rect 380083 210218 380125 210454
rect 379805 210134 380125 210218
rect 379805 209898 379847 210134
rect 380083 209898 380125 210134
rect 379805 209866 380125 209898
rect 400874 210454 401194 210486
rect 400874 210218 400916 210454
rect 401152 210218 401194 210454
rect 400874 210134 401194 210218
rect 400874 209898 400916 210134
rect 401152 209898 401194 210134
rect 400874 209866 401194 209898
rect 406805 210454 407125 210486
rect 406805 210218 406847 210454
rect 407083 210218 407125 210454
rect 406805 210134 407125 210218
rect 406805 209898 406847 210134
rect 407083 209898 407125 210134
rect 406805 209866 407125 209898
rect 427874 210454 428194 210486
rect 427874 210218 427916 210454
rect 428152 210218 428194 210454
rect 427874 210134 428194 210218
rect 427874 209898 427916 210134
rect 428152 209898 428194 210134
rect 427874 209866 428194 209898
rect 433805 210454 434125 210486
rect 433805 210218 433847 210454
rect 434083 210218 434125 210454
rect 433805 210134 434125 210218
rect 433805 209898 433847 210134
rect 434083 209898 434125 210134
rect 433805 209866 434125 209898
rect 454874 210454 455194 210486
rect 454874 210218 454916 210454
rect 455152 210218 455194 210454
rect 454874 210134 455194 210218
rect 454874 209898 454916 210134
rect 455152 209898 455194 210134
rect 454874 209866 455194 209898
rect 460805 210454 461125 210486
rect 460805 210218 460847 210454
rect 461083 210218 461125 210454
rect 460805 210134 461125 210218
rect 460805 209898 460847 210134
rect 461083 209898 461125 210134
rect 460805 209866 461125 209898
rect 481874 210454 482194 210486
rect 481874 210218 481916 210454
rect 482152 210218 482194 210454
rect 481874 210134 482194 210218
rect 481874 209898 481916 210134
rect 482152 209898 482194 210134
rect 481874 209866 482194 209898
rect 487805 210454 488125 210486
rect 487805 210218 487847 210454
rect 488083 210218 488125 210454
rect 487805 210134 488125 210218
rect 487805 209898 487847 210134
rect 488083 209898 488125 210134
rect 487805 209866 488125 209898
rect 508874 210454 509194 210486
rect 508874 210218 508916 210454
rect 509152 210218 509194 210454
rect 508874 210134 509194 210218
rect 508874 209898 508916 210134
rect 509152 209898 509194 210134
rect 508874 209866 509194 209898
rect 514805 210454 515125 210486
rect 514805 210218 514847 210454
rect 515083 210218 515125 210454
rect 514805 210134 515125 210218
rect 514805 209898 514847 210134
rect 515083 209898 515125 210134
rect 514805 209866 515125 209898
rect 535874 210454 536194 210486
rect 535874 210218 535916 210454
rect 536152 210218 536194 210454
rect 535874 210134 536194 210218
rect 535874 209898 535916 210134
rect 536152 209898 536194 210134
rect 535874 209866 536194 209898
rect 541805 210454 542125 210486
rect 541805 210218 541847 210454
rect 542083 210218 542125 210454
rect 541805 210134 542125 210218
rect 541805 209898 541847 210134
rect 542083 209898 542125 210134
rect 541805 209866 542125 209898
rect 19794 201454 20414 203000
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 200000 20414 200898
rect 28794 202394 29414 203000
rect 28794 202158 28826 202394
rect 29062 202158 29146 202394
rect 29382 202158 29414 202394
rect 28794 202074 29414 202158
rect 28794 201838 28826 202074
rect 29062 201838 29146 202074
rect 29382 201838 29414 202074
rect 28794 200000 29414 201838
rect 37794 201454 38414 203000
rect 37794 201218 37826 201454
rect 38062 201218 38146 201454
rect 38382 201218 38414 201454
rect 37794 201134 38414 201218
rect 37794 200898 37826 201134
rect 38062 200898 38146 201134
rect 38382 200898 38414 201134
rect 37794 200000 38414 200898
rect 46794 202394 47414 203000
rect 46794 202158 46826 202394
rect 47062 202158 47146 202394
rect 47382 202158 47414 202394
rect 46794 202074 47414 202158
rect 46794 201838 46826 202074
rect 47062 201838 47146 202074
rect 47382 201838 47414 202074
rect 46794 200000 47414 201838
rect 55794 201454 56414 203000
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 200000 56414 200898
rect 64794 202394 65414 203000
rect 64794 202158 64826 202394
rect 65062 202158 65146 202394
rect 65382 202158 65414 202394
rect 64794 202074 65414 202158
rect 64794 201838 64826 202074
rect 65062 201838 65146 202074
rect 65382 201838 65414 202074
rect 64794 200000 65414 201838
rect 73794 201454 74414 203000
rect 73794 201218 73826 201454
rect 74062 201218 74146 201454
rect 74382 201218 74414 201454
rect 73794 201134 74414 201218
rect 73794 200898 73826 201134
rect 74062 200898 74146 201134
rect 74382 200898 74414 201134
rect 73794 200000 74414 200898
rect 82794 202394 83414 203000
rect 82794 202158 82826 202394
rect 83062 202158 83146 202394
rect 83382 202158 83414 202394
rect 82794 202074 83414 202158
rect 82794 201838 82826 202074
rect 83062 201838 83146 202074
rect 83382 201838 83414 202074
rect 82794 200000 83414 201838
rect 91794 201454 92414 203000
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 200000 92414 200898
rect 100794 202394 101414 203000
rect 100794 202158 100826 202394
rect 101062 202158 101146 202394
rect 101382 202158 101414 202394
rect 100794 202074 101414 202158
rect 100794 201838 100826 202074
rect 101062 201838 101146 202074
rect 101382 201838 101414 202074
rect 100794 200000 101414 201838
rect 109794 201454 110414 203000
rect 109794 201218 109826 201454
rect 110062 201218 110146 201454
rect 110382 201218 110414 201454
rect 109794 201134 110414 201218
rect 109794 200898 109826 201134
rect 110062 200898 110146 201134
rect 110382 200898 110414 201134
rect 109794 200000 110414 200898
rect 118794 202394 119414 203000
rect 118794 202158 118826 202394
rect 119062 202158 119146 202394
rect 119382 202158 119414 202394
rect 118794 202074 119414 202158
rect 118794 201838 118826 202074
rect 119062 201838 119146 202074
rect 119382 201838 119414 202074
rect 118794 200000 119414 201838
rect 127794 201454 128414 203000
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 200000 128414 200898
rect 136794 202394 137414 203000
rect 136794 202158 136826 202394
rect 137062 202158 137146 202394
rect 137382 202158 137414 202394
rect 136794 202074 137414 202158
rect 136794 201838 136826 202074
rect 137062 201838 137146 202074
rect 137382 201838 137414 202074
rect 136794 200000 137414 201838
rect 145794 201454 146414 203000
rect 145794 201218 145826 201454
rect 146062 201218 146146 201454
rect 146382 201218 146414 201454
rect 145794 201134 146414 201218
rect 145794 200898 145826 201134
rect 146062 200898 146146 201134
rect 146382 200898 146414 201134
rect 145794 200000 146414 200898
rect 154794 202394 155414 203000
rect 154794 202158 154826 202394
rect 155062 202158 155146 202394
rect 155382 202158 155414 202394
rect 154794 202074 155414 202158
rect 154794 201838 154826 202074
rect 155062 201838 155146 202074
rect 155382 201838 155414 202074
rect 154794 200000 155414 201838
rect 163794 201454 164414 203000
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 200000 164414 200898
rect 172794 202394 173414 203000
rect 172794 202158 172826 202394
rect 173062 202158 173146 202394
rect 173382 202158 173414 202394
rect 172794 202074 173414 202158
rect 172794 201838 172826 202074
rect 173062 201838 173146 202074
rect 173382 201838 173414 202074
rect 172794 200000 173414 201838
rect 181794 201454 182414 203000
rect 181794 201218 181826 201454
rect 182062 201218 182146 201454
rect 182382 201218 182414 201454
rect 181794 201134 182414 201218
rect 181794 200898 181826 201134
rect 182062 200898 182146 201134
rect 182382 200898 182414 201134
rect 181794 200000 182414 200898
rect 190794 202394 191414 203000
rect 190794 202158 190826 202394
rect 191062 202158 191146 202394
rect 191382 202158 191414 202394
rect 190794 202074 191414 202158
rect 190794 201838 190826 202074
rect 191062 201838 191146 202074
rect 191382 201838 191414 202074
rect 190794 200000 191414 201838
rect 199794 201454 200414 203000
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 200000 200414 200898
rect 208794 202394 209414 203000
rect 208794 202158 208826 202394
rect 209062 202158 209146 202394
rect 209382 202158 209414 202394
rect 208794 202074 209414 202158
rect 208794 201838 208826 202074
rect 209062 201838 209146 202074
rect 209382 201838 209414 202074
rect 208794 200000 209414 201838
rect 217794 201454 218414 203000
rect 217794 201218 217826 201454
rect 218062 201218 218146 201454
rect 218382 201218 218414 201454
rect 217794 201134 218414 201218
rect 217794 200898 217826 201134
rect 218062 200898 218146 201134
rect 218382 200898 218414 201134
rect 217794 200000 218414 200898
rect 226794 202394 227414 203000
rect 226794 202158 226826 202394
rect 227062 202158 227146 202394
rect 227382 202158 227414 202394
rect 226794 202074 227414 202158
rect 226794 201838 226826 202074
rect 227062 201838 227146 202074
rect 227382 201838 227414 202074
rect 226794 200000 227414 201838
rect 235794 201454 236414 203000
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 200000 236414 200898
rect 244794 202394 245414 203000
rect 244794 202158 244826 202394
rect 245062 202158 245146 202394
rect 245382 202158 245414 202394
rect 244794 202074 245414 202158
rect 244794 201838 244826 202074
rect 245062 201838 245146 202074
rect 245382 201838 245414 202074
rect 244794 200000 245414 201838
rect 253794 201454 254414 203000
rect 253794 201218 253826 201454
rect 254062 201218 254146 201454
rect 254382 201218 254414 201454
rect 253794 201134 254414 201218
rect 253794 200898 253826 201134
rect 254062 200898 254146 201134
rect 254382 200898 254414 201134
rect 253794 200000 254414 200898
rect 262794 202394 263414 203000
rect 262794 202158 262826 202394
rect 263062 202158 263146 202394
rect 263382 202158 263414 202394
rect 262794 202074 263414 202158
rect 262794 201838 262826 202074
rect 263062 201838 263146 202074
rect 263382 201838 263414 202074
rect 262794 200000 263414 201838
rect 271794 201454 272414 203000
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 200000 272414 200898
rect 280794 202394 281414 203000
rect 280794 202158 280826 202394
rect 281062 202158 281146 202394
rect 281382 202158 281414 202394
rect 280794 202074 281414 202158
rect 280794 201838 280826 202074
rect 281062 201838 281146 202074
rect 281382 201838 281414 202074
rect 280794 200000 281414 201838
rect 289794 201454 290414 203000
rect 289794 201218 289826 201454
rect 290062 201218 290146 201454
rect 290382 201218 290414 201454
rect 289794 201134 290414 201218
rect 289794 200898 289826 201134
rect 290062 200898 290146 201134
rect 290382 200898 290414 201134
rect 289794 200000 290414 200898
rect 298794 202394 299414 203000
rect 298794 202158 298826 202394
rect 299062 202158 299146 202394
rect 299382 202158 299414 202394
rect 298794 202074 299414 202158
rect 298794 201838 298826 202074
rect 299062 201838 299146 202074
rect 299382 201838 299414 202074
rect 298794 200000 299414 201838
rect 307794 201454 308414 203000
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 200000 308414 200898
rect 316794 202394 317414 203000
rect 316794 202158 316826 202394
rect 317062 202158 317146 202394
rect 317382 202158 317414 202394
rect 316794 202074 317414 202158
rect 316794 201838 316826 202074
rect 317062 201838 317146 202074
rect 317382 201838 317414 202074
rect 316794 200000 317414 201838
rect 325794 201454 326414 203000
rect 325794 201218 325826 201454
rect 326062 201218 326146 201454
rect 326382 201218 326414 201454
rect 325794 201134 326414 201218
rect 325794 200898 325826 201134
rect 326062 200898 326146 201134
rect 326382 200898 326414 201134
rect 325794 200000 326414 200898
rect 334794 202394 335414 203000
rect 334794 202158 334826 202394
rect 335062 202158 335146 202394
rect 335382 202158 335414 202394
rect 334794 202074 335414 202158
rect 334794 201838 334826 202074
rect 335062 201838 335146 202074
rect 335382 201838 335414 202074
rect 334794 200000 335414 201838
rect 343794 201454 344414 203000
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 200000 344414 200898
rect 352794 202394 353414 203000
rect 352794 202158 352826 202394
rect 353062 202158 353146 202394
rect 353382 202158 353414 202394
rect 352794 202074 353414 202158
rect 352794 201838 352826 202074
rect 353062 201838 353146 202074
rect 353382 201838 353414 202074
rect 352794 200000 353414 201838
rect 361794 201454 362414 203000
rect 361794 201218 361826 201454
rect 362062 201218 362146 201454
rect 362382 201218 362414 201454
rect 361794 201134 362414 201218
rect 361794 200898 361826 201134
rect 362062 200898 362146 201134
rect 362382 200898 362414 201134
rect 361794 200000 362414 200898
rect 370794 202394 371414 203000
rect 370794 202158 370826 202394
rect 371062 202158 371146 202394
rect 371382 202158 371414 202394
rect 370794 202074 371414 202158
rect 370794 201838 370826 202074
rect 371062 201838 371146 202074
rect 371382 201838 371414 202074
rect 370794 200000 371414 201838
rect 379794 201454 380414 203000
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 200000 380414 200898
rect 388794 202394 389414 203000
rect 388794 202158 388826 202394
rect 389062 202158 389146 202394
rect 389382 202158 389414 202394
rect 388794 202074 389414 202158
rect 388794 201838 388826 202074
rect 389062 201838 389146 202074
rect 389382 201838 389414 202074
rect 388794 200000 389414 201838
rect 397794 201454 398414 203000
rect 397794 201218 397826 201454
rect 398062 201218 398146 201454
rect 398382 201218 398414 201454
rect 397794 201134 398414 201218
rect 397794 200898 397826 201134
rect 398062 200898 398146 201134
rect 398382 200898 398414 201134
rect 397794 200000 398414 200898
rect 406794 202394 407414 203000
rect 406794 202158 406826 202394
rect 407062 202158 407146 202394
rect 407382 202158 407414 202394
rect 406794 202074 407414 202158
rect 406794 201838 406826 202074
rect 407062 201838 407146 202074
rect 407382 201838 407414 202074
rect 406794 200000 407414 201838
rect 415794 201454 416414 203000
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 200000 416414 200898
rect 424794 202394 425414 203000
rect 424794 202158 424826 202394
rect 425062 202158 425146 202394
rect 425382 202158 425414 202394
rect 424794 202074 425414 202158
rect 424794 201838 424826 202074
rect 425062 201838 425146 202074
rect 425382 201838 425414 202074
rect 424794 200000 425414 201838
rect 433794 201454 434414 203000
rect 433794 201218 433826 201454
rect 434062 201218 434146 201454
rect 434382 201218 434414 201454
rect 433794 201134 434414 201218
rect 433794 200898 433826 201134
rect 434062 200898 434146 201134
rect 434382 200898 434414 201134
rect 433794 200000 434414 200898
rect 442794 202394 443414 203000
rect 442794 202158 442826 202394
rect 443062 202158 443146 202394
rect 443382 202158 443414 202394
rect 442794 202074 443414 202158
rect 442794 201838 442826 202074
rect 443062 201838 443146 202074
rect 443382 201838 443414 202074
rect 442794 200000 443414 201838
rect 451794 201454 452414 203000
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 200000 452414 200898
rect 460794 202394 461414 203000
rect 460794 202158 460826 202394
rect 461062 202158 461146 202394
rect 461382 202158 461414 202394
rect 460794 202074 461414 202158
rect 460794 201838 460826 202074
rect 461062 201838 461146 202074
rect 461382 201838 461414 202074
rect 460794 200000 461414 201838
rect 469794 201454 470414 203000
rect 469794 201218 469826 201454
rect 470062 201218 470146 201454
rect 470382 201218 470414 201454
rect 469794 201134 470414 201218
rect 469794 200898 469826 201134
rect 470062 200898 470146 201134
rect 470382 200898 470414 201134
rect 469794 200000 470414 200898
rect 478794 202394 479414 203000
rect 478794 202158 478826 202394
rect 479062 202158 479146 202394
rect 479382 202158 479414 202394
rect 478794 202074 479414 202158
rect 478794 201838 478826 202074
rect 479062 201838 479146 202074
rect 479382 201838 479414 202074
rect 478794 200000 479414 201838
rect 487794 201454 488414 203000
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 200000 488414 200898
rect 496794 202394 497414 203000
rect 496794 202158 496826 202394
rect 497062 202158 497146 202394
rect 497382 202158 497414 202394
rect 496794 202074 497414 202158
rect 496794 201838 496826 202074
rect 497062 201838 497146 202074
rect 497382 201838 497414 202074
rect 496794 200000 497414 201838
rect 505794 201454 506414 203000
rect 505794 201218 505826 201454
rect 506062 201218 506146 201454
rect 506382 201218 506414 201454
rect 505794 201134 506414 201218
rect 505794 200898 505826 201134
rect 506062 200898 506146 201134
rect 506382 200898 506414 201134
rect 505794 200000 506414 200898
rect 514794 202394 515414 203000
rect 514794 202158 514826 202394
rect 515062 202158 515146 202394
rect 515382 202158 515414 202394
rect 514794 202074 515414 202158
rect 514794 201838 514826 202074
rect 515062 201838 515146 202074
rect 515382 201838 515414 202074
rect 514794 200000 515414 201838
rect 523794 201454 524414 203000
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 200000 524414 200898
rect 532794 202394 533414 203000
rect 532794 202158 532826 202394
rect 533062 202158 533146 202394
rect 533382 202158 533414 202394
rect 532794 202074 533414 202158
rect 532794 201838 532826 202074
rect 533062 201838 533146 202074
rect 533382 201838 533414 202074
rect 532794 200000 533414 201838
rect 541794 201454 542414 203000
rect 541794 201218 541826 201454
rect 542062 201218 542146 201454
rect 542382 201218 542414 201454
rect 541794 201134 542414 201218
rect 541794 200898 541826 201134
rect 542062 200898 542146 201134
rect 542382 200898 542414 201134
rect 541794 200000 542414 200898
rect 550794 202394 551414 203000
rect 550794 202158 550826 202394
rect 551062 202158 551146 202394
rect 551382 202158 551414 202394
rect 550794 202074 551414 202158
rect 550794 201838 550826 202074
rect 551062 201838 551146 202074
rect 551382 201838 551414 202074
rect 550794 200000 551414 201838
rect 559794 201454 560414 218898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 174454 11414 191898
rect 22874 192454 23194 192486
rect 22874 192218 22916 192454
rect 23152 192218 23194 192454
rect 22874 192134 23194 192218
rect 22874 191898 22916 192134
rect 23152 191898 23194 192134
rect 22874 191866 23194 191898
rect 28805 192454 29125 192486
rect 28805 192218 28847 192454
rect 29083 192218 29125 192454
rect 28805 192134 29125 192218
rect 28805 191898 28847 192134
rect 29083 191898 29125 192134
rect 28805 191866 29125 191898
rect 49874 192454 50194 192486
rect 49874 192218 49916 192454
rect 50152 192218 50194 192454
rect 49874 192134 50194 192218
rect 49874 191898 49916 192134
rect 50152 191898 50194 192134
rect 49874 191866 50194 191898
rect 55805 192454 56125 192486
rect 55805 192218 55847 192454
rect 56083 192218 56125 192454
rect 55805 192134 56125 192218
rect 55805 191898 55847 192134
rect 56083 191898 56125 192134
rect 55805 191866 56125 191898
rect 76874 192454 77194 192486
rect 76874 192218 76916 192454
rect 77152 192218 77194 192454
rect 76874 192134 77194 192218
rect 76874 191898 76916 192134
rect 77152 191898 77194 192134
rect 76874 191866 77194 191898
rect 82805 192454 83125 192486
rect 82805 192218 82847 192454
rect 83083 192218 83125 192454
rect 82805 192134 83125 192218
rect 82805 191898 82847 192134
rect 83083 191898 83125 192134
rect 82805 191866 83125 191898
rect 103874 192454 104194 192486
rect 103874 192218 103916 192454
rect 104152 192218 104194 192454
rect 103874 192134 104194 192218
rect 103874 191898 103916 192134
rect 104152 191898 104194 192134
rect 103874 191866 104194 191898
rect 109805 192454 110125 192486
rect 109805 192218 109847 192454
rect 110083 192218 110125 192454
rect 109805 192134 110125 192218
rect 109805 191898 109847 192134
rect 110083 191898 110125 192134
rect 109805 191866 110125 191898
rect 130874 192454 131194 192486
rect 130874 192218 130916 192454
rect 131152 192218 131194 192454
rect 130874 192134 131194 192218
rect 130874 191898 130916 192134
rect 131152 191898 131194 192134
rect 130874 191866 131194 191898
rect 136805 192454 137125 192486
rect 136805 192218 136847 192454
rect 137083 192218 137125 192454
rect 136805 192134 137125 192218
rect 136805 191898 136847 192134
rect 137083 191898 137125 192134
rect 136805 191866 137125 191898
rect 157874 192454 158194 192486
rect 157874 192218 157916 192454
rect 158152 192218 158194 192454
rect 157874 192134 158194 192218
rect 157874 191898 157916 192134
rect 158152 191898 158194 192134
rect 157874 191866 158194 191898
rect 163805 192454 164125 192486
rect 163805 192218 163847 192454
rect 164083 192218 164125 192454
rect 163805 192134 164125 192218
rect 163805 191898 163847 192134
rect 164083 191898 164125 192134
rect 163805 191866 164125 191898
rect 184874 192454 185194 192486
rect 184874 192218 184916 192454
rect 185152 192218 185194 192454
rect 184874 192134 185194 192218
rect 184874 191898 184916 192134
rect 185152 191898 185194 192134
rect 184874 191866 185194 191898
rect 190805 192454 191125 192486
rect 190805 192218 190847 192454
rect 191083 192218 191125 192454
rect 190805 192134 191125 192218
rect 190805 191898 190847 192134
rect 191083 191898 191125 192134
rect 190805 191866 191125 191898
rect 211874 192454 212194 192486
rect 211874 192218 211916 192454
rect 212152 192218 212194 192454
rect 211874 192134 212194 192218
rect 211874 191898 211916 192134
rect 212152 191898 212194 192134
rect 211874 191866 212194 191898
rect 217805 192454 218125 192486
rect 217805 192218 217847 192454
rect 218083 192218 218125 192454
rect 217805 192134 218125 192218
rect 217805 191898 217847 192134
rect 218083 191898 218125 192134
rect 217805 191866 218125 191898
rect 238874 192454 239194 192486
rect 238874 192218 238916 192454
rect 239152 192218 239194 192454
rect 238874 192134 239194 192218
rect 238874 191898 238916 192134
rect 239152 191898 239194 192134
rect 238874 191866 239194 191898
rect 244805 192454 245125 192486
rect 244805 192218 244847 192454
rect 245083 192218 245125 192454
rect 244805 192134 245125 192218
rect 244805 191898 244847 192134
rect 245083 191898 245125 192134
rect 244805 191866 245125 191898
rect 265874 192454 266194 192486
rect 265874 192218 265916 192454
rect 266152 192218 266194 192454
rect 265874 192134 266194 192218
rect 265874 191898 265916 192134
rect 266152 191898 266194 192134
rect 265874 191866 266194 191898
rect 271805 192454 272125 192486
rect 271805 192218 271847 192454
rect 272083 192218 272125 192454
rect 271805 192134 272125 192218
rect 271805 191898 271847 192134
rect 272083 191898 272125 192134
rect 271805 191866 272125 191898
rect 292874 192454 293194 192486
rect 292874 192218 292916 192454
rect 293152 192218 293194 192454
rect 292874 192134 293194 192218
rect 292874 191898 292916 192134
rect 293152 191898 293194 192134
rect 292874 191866 293194 191898
rect 298805 192454 299125 192486
rect 298805 192218 298847 192454
rect 299083 192218 299125 192454
rect 298805 192134 299125 192218
rect 298805 191898 298847 192134
rect 299083 191898 299125 192134
rect 298805 191866 299125 191898
rect 319874 192454 320194 192486
rect 319874 192218 319916 192454
rect 320152 192218 320194 192454
rect 319874 192134 320194 192218
rect 319874 191898 319916 192134
rect 320152 191898 320194 192134
rect 319874 191866 320194 191898
rect 325805 192454 326125 192486
rect 325805 192218 325847 192454
rect 326083 192218 326125 192454
rect 325805 192134 326125 192218
rect 325805 191898 325847 192134
rect 326083 191898 326125 192134
rect 325805 191866 326125 191898
rect 346874 192454 347194 192486
rect 346874 192218 346916 192454
rect 347152 192218 347194 192454
rect 346874 192134 347194 192218
rect 346874 191898 346916 192134
rect 347152 191898 347194 192134
rect 346874 191866 347194 191898
rect 352805 192454 353125 192486
rect 352805 192218 352847 192454
rect 353083 192218 353125 192454
rect 352805 192134 353125 192218
rect 352805 191898 352847 192134
rect 353083 191898 353125 192134
rect 352805 191866 353125 191898
rect 373874 192454 374194 192486
rect 373874 192218 373916 192454
rect 374152 192218 374194 192454
rect 373874 192134 374194 192218
rect 373874 191898 373916 192134
rect 374152 191898 374194 192134
rect 373874 191866 374194 191898
rect 379805 192454 380125 192486
rect 379805 192218 379847 192454
rect 380083 192218 380125 192454
rect 379805 192134 380125 192218
rect 379805 191898 379847 192134
rect 380083 191898 380125 192134
rect 379805 191866 380125 191898
rect 400874 192454 401194 192486
rect 400874 192218 400916 192454
rect 401152 192218 401194 192454
rect 400874 192134 401194 192218
rect 400874 191898 400916 192134
rect 401152 191898 401194 192134
rect 400874 191866 401194 191898
rect 406805 192454 407125 192486
rect 406805 192218 406847 192454
rect 407083 192218 407125 192454
rect 406805 192134 407125 192218
rect 406805 191898 406847 192134
rect 407083 191898 407125 192134
rect 406805 191866 407125 191898
rect 427874 192454 428194 192486
rect 427874 192218 427916 192454
rect 428152 192218 428194 192454
rect 427874 192134 428194 192218
rect 427874 191898 427916 192134
rect 428152 191898 428194 192134
rect 427874 191866 428194 191898
rect 433805 192454 434125 192486
rect 433805 192218 433847 192454
rect 434083 192218 434125 192454
rect 433805 192134 434125 192218
rect 433805 191898 433847 192134
rect 434083 191898 434125 192134
rect 433805 191866 434125 191898
rect 454874 192454 455194 192486
rect 454874 192218 454916 192454
rect 455152 192218 455194 192454
rect 454874 192134 455194 192218
rect 454874 191898 454916 192134
rect 455152 191898 455194 192134
rect 454874 191866 455194 191898
rect 460805 192454 461125 192486
rect 460805 192218 460847 192454
rect 461083 192218 461125 192454
rect 460805 192134 461125 192218
rect 460805 191898 460847 192134
rect 461083 191898 461125 192134
rect 460805 191866 461125 191898
rect 481874 192454 482194 192486
rect 481874 192218 481916 192454
rect 482152 192218 482194 192454
rect 481874 192134 482194 192218
rect 481874 191898 481916 192134
rect 482152 191898 482194 192134
rect 481874 191866 482194 191898
rect 487805 192454 488125 192486
rect 487805 192218 487847 192454
rect 488083 192218 488125 192454
rect 487805 192134 488125 192218
rect 487805 191898 487847 192134
rect 488083 191898 488125 192134
rect 487805 191866 488125 191898
rect 508874 192454 509194 192486
rect 508874 192218 508916 192454
rect 509152 192218 509194 192454
rect 508874 192134 509194 192218
rect 508874 191898 508916 192134
rect 509152 191898 509194 192134
rect 508874 191866 509194 191898
rect 514805 192454 515125 192486
rect 514805 192218 514847 192454
rect 515083 192218 515125 192454
rect 514805 192134 515125 192218
rect 514805 191898 514847 192134
rect 515083 191898 515125 192134
rect 514805 191866 515125 191898
rect 535874 192454 536194 192486
rect 535874 192218 535916 192454
rect 536152 192218 536194 192454
rect 535874 192134 536194 192218
rect 535874 191898 535916 192134
rect 536152 191898 536194 192134
rect 535874 191866 536194 191898
rect 541805 192454 542125 192486
rect 541805 192218 541847 192454
rect 542083 192218 542125 192454
rect 541805 192134 542125 192218
rect 541805 191898 541847 192134
rect 542083 191898 542125 192134
rect 541805 191866 542125 191898
rect 19910 183454 20230 183486
rect 19910 183218 19952 183454
rect 20188 183218 20230 183454
rect 19910 183134 20230 183218
rect 19910 182898 19952 183134
rect 20188 182898 20230 183134
rect 19910 182866 20230 182898
rect 25840 183454 26160 183486
rect 25840 183218 25882 183454
rect 26118 183218 26160 183454
rect 25840 183134 26160 183218
rect 25840 182898 25882 183134
rect 26118 182898 26160 183134
rect 25840 182866 26160 182898
rect 31771 183454 32091 183486
rect 31771 183218 31813 183454
rect 32049 183218 32091 183454
rect 31771 183134 32091 183218
rect 31771 182898 31813 183134
rect 32049 182898 32091 183134
rect 31771 182866 32091 182898
rect 46910 183454 47230 183486
rect 46910 183218 46952 183454
rect 47188 183218 47230 183454
rect 46910 183134 47230 183218
rect 46910 182898 46952 183134
rect 47188 182898 47230 183134
rect 46910 182866 47230 182898
rect 52840 183454 53160 183486
rect 52840 183218 52882 183454
rect 53118 183218 53160 183454
rect 52840 183134 53160 183218
rect 52840 182898 52882 183134
rect 53118 182898 53160 183134
rect 52840 182866 53160 182898
rect 58771 183454 59091 183486
rect 58771 183218 58813 183454
rect 59049 183218 59091 183454
rect 58771 183134 59091 183218
rect 58771 182898 58813 183134
rect 59049 182898 59091 183134
rect 58771 182866 59091 182898
rect 73910 183454 74230 183486
rect 73910 183218 73952 183454
rect 74188 183218 74230 183454
rect 73910 183134 74230 183218
rect 73910 182898 73952 183134
rect 74188 182898 74230 183134
rect 73910 182866 74230 182898
rect 79840 183454 80160 183486
rect 79840 183218 79882 183454
rect 80118 183218 80160 183454
rect 79840 183134 80160 183218
rect 79840 182898 79882 183134
rect 80118 182898 80160 183134
rect 79840 182866 80160 182898
rect 85771 183454 86091 183486
rect 85771 183218 85813 183454
rect 86049 183218 86091 183454
rect 85771 183134 86091 183218
rect 85771 182898 85813 183134
rect 86049 182898 86091 183134
rect 85771 182866 86091 182898
rect 100910 183454 101230 183486
rect 100910 183218 100952 183454
rect 101188 183218 101230 183454
rect 100910 183134 101230 183218
rect 100910 182898 100952 183134
rect 101188 182898 101230 183134
rect 100910 182866 101230 182898
rect 106840 183454 107160 183486
rect 106840 183218 106882 183454
rect 107118 183218 107160 183454
rect 106840 183134 107160 183218
rect 106840 182898 106882 183134
rect 107118 182898 107160 183134
rect 106840 182866 107160 182898
rect 112771 183454 113091 183486
rect 112771 183218 112813 183454
rect 113049 183218 113091 183454
rect 112771 183134 113091 183218
rect 112771 182898 112813 183134
rect 113049 182898 113091 183134
rect 112771 182866 113091 182898
rect 127910 183454 128230 183486
rect 127910 183218 127952 183454
rect 128188 183218 128230 183454
rect 127910 183134 128230 183218
rect 127910 182898 127952 183134
rect 128188 182898 128230 183134
rect 127910 182866 128230 182898
rect 133840 183454 134160 183486
rect 133840 183218 133882 183454
rect 134118 183218 134160 183454
rect 133840 183134 134160 183218
rect 133840 182898 133882 183134
rect 134118 182898 134160 183134
rect 133840 182866 134160 182898
rect 139771 183454 140091 183486
rect 139771 183218 139813 183454
rect 140049 183218 140091 183454
rect 139771 183134 140091 183218
rect 139771 182898 139813 183134
rect 140049 182898 140091 183134
rect 139771 182866 140091 182898
rect 154910 183454 155230 183486
rect 154910 183218 154952 183454
rect 155188 183218 155230 183454
rect 154910 183134 155230 183218
rect 154910 182898 154952 183134
rect 155188 182898 155230 183134
rect 154910 182866 155230 182898
rect 160840 183454 161160 183486
rect 160840 183218 160882 183454
rect 161118 183218 161160 183454
rect 160840 183134 161160 183218
rect 160840 182898 160882 183134
rect 161118 182898 161160 183134
rect 160840 182866 161160 182898
rect 166771 183454 167091 183486
rect 166771 183218 166813 183454
rect 167049 183218 167091 183454
rect 166771 183134 167091 183218
rect 166771 182898 166813 183134
rect 167049 182898 167091 183134
rect 166771 182866 167091 182898
rect 181910 183454 182230 183486
rect 181910 183218 181952 183454
rect 182188 183218 182230 183454
rect 181910 183134 182230 183218
rect 181910 182898 181952 183134
rect 182188 182898 182230 183134
rect 181910 182866 182230 182898
rect 187840 183454 188160 183486
rect 187840 183218 187882 183454
rect 188118 183218 188160 183454
rect 187840 183134 188160 183218
rect 187840 182898 187882 183134
rect 188118 182898 188160 183134
rect 187840 182866 188160 182898
rect 193771 183454 194091 183486
rect 193771 183218 193813 183454
rect 194049 183218 194091 183454
rect 193771 183134 194091 183218
rect 193771 182898 193813 183134
rect 194049 182898 194091 183134
rect 193771 182866 194091 182898
rect 208910 183454 209230 183486
rect 208910 183218 208952 183454
rect 209188 183218 209230 183454
rect 208910 183134 209230 183218
rect 208910 182898 208952 183134
rect 209188 182898 209230 183134
rect 208910 182866 209230 182898
rect 214840 183454 215160 183486
rect 214840 183218 214882 183454
rect 215118 183218 215160 183454
rect 214840 183134 215160 183218
rect 214840 182898 214882 183134
rect 215118 182898 215160 183134
rect 214840 182866 215160 182898
rect 220771 183454 221091 183486
rect 220771 183218 220813 183454
rect 221049 183218 221091 183454
rect 220771 183134 221091 183218
rect 220771 182898 220813 183134
rect 221049 182898 221091 183134
rect 220771 182866 221091 182898
rect 235910 183454 236230 183486
rect 235910 183218 235952 183454
rect 236188 183218 236230 183454
rect 235910 183134 236230 183218
rect 235910 182898 235952 183134
rect 236188 182898 236230 183134
rect 235910 182866 236230 182898
rect 241840 183454 242160 183486
rect 241840 183218 241882 183454
rect 242118 183218 242160 183454
rect 241840 183134 242160 183218
rect 241840 182898 241882 183134
rect 242118 182898 242160 183134
rect 241840 182866 242160 182898
rect 247771 183454 248091 183486
rect 247771 183218 247813 183454
rect 248049 183218 248091 183454
rect 247771 183134 248091 183218
rect 247771 182898 247813 183134
rect 248049 182898 248091 183134
rect 247771 182866 248091 182898
rect 262910 183454 263230 183486
rect 262910 183218 262952 183454
rect 263188 183218 263230 183454
rect 262910 183134 263230 183218
rect 262910 182898 262952 183134
rect 263188 182898 263230 183134
rect 262910 182866 263230 182898
rect 268840 183454 269160 183486
rect 268840 183218 268882 183454
rect 269118 183218 269160 183454
rect 268840 183134 269160 183218
rect 268840 182898 268882 183134
rect 269118 182898 269160 183134
rect 268840 182866 269160 182898
rect 274771 183454 275091 183486
rect 274771 183218 274813 183454
rect 275049 183218 275091 183454
rect 274771 183134 275091 183218
rect 274771 182898 274813 183134
rect 275049 182898 275091 183134
rect 274771 182866 275091 182898
rect 289910 183454 290230 183486
rect 289910 183218 289952 183454
rect 290188 183218 290230 183454
rect 289910 183134 290230 183218
rect 289910 182898 289952 183134
rect 290188 182898 290230 183134
rect 289910 182866 290230 182898
rect 295840 183454 296160 183486
rect 295840 183218 295882 183454
rect 296118 183218 296160 183454
rect 295840 183134 296160 183218
rect 295840 182898 295882 183134
rect 296118 182898 296160 183134
rect 295840 182866 296160 182898
rect 301771 183454 302091 183486
rect 301771 183218 301813 183454
rect 302049 183218 302091 183454
rect 301771 183134 302091 183218
rect 301771 182898 301813 183134
rect 302049 182898 302091 183134
rect 301771 182866 302091 182898
rect 316910 183454 317230 183486
rect 316910 183218 316952 183454
rect 317188 183218 317230 183454
rect 316910 183134 317230 183218
rect 316910 182898 316952 183134
rect 317188 182898 317230 183134
rect 316910 182866 317230 182898
rect 322840 183454 323160 183486
rect 322840 183218 322882 183454
rect 323118 183218 323160 183454
rect 322840 183134 323160 183218
rect 322840 182898 322882 183134
rect 323118 182898 323160 183134
rect 322840 182866 323160 182898
rect 328771 183454 329091 183486
rect 328771 183218 328813 183454
rect 329049 183218 329091 183454
rect 328771 183134 329091 183218
rect 328771 182898 328813 183134
rect 329049 182898 329091 183134
rect 328771 182866 329091 182898
rect 343910 183454 344230 183486
rect 343910 183218 343952 183454
rect 344188 183218 344230 183454
rect 343910 183134 344230 183218
rect 343910 182898 343952 183134
rect 344188 182898 344230 183134
rect 343910 182866 344230 182898
rect 349840 183454 350160 183486
rect 349840 183218 349882 183454
rect 350118 183218 350160 183454
rect 349840 183134 350160 183218
rect 349840 182898 349882 183134
rect 350118 182898 350160 183134
rect 349840 182866 350160 182898
rect 355771 183454 356091 183486
rect 355771 183218 355813 183454
rect 356049 183218 356091 183454
rect 355771 183134 356091 183218
rect 355771 182898 355813 183134
rect 356049 182898 356091 183134
rect 355771 182866 356091 182898
rect 370910 183454 371230 183486
rect 370910 183218 370952 183454
rect 371188 183218 371230 183454
rect 370910 183134 371230 183218
rect 370910 182898 370952 183134
rect 371188 182898 371230 183134
rect 370910 182866 371230 182898
rect 376840 183454 377160 183486
rect 376840 183218 376882 183454
rect 377118 183218 377160 183454
rect 376840 183134 377160 183218
rect 376840 182898 376882 183134
rect 377118 182898 377160 183134
rect 376840 182866 377160 182898
rect 382771 183454 383091 183486
rect 382771 183218 382813 183454
rect 383049 183218 383091 183454
rect 382771 183134 383091 183218
rect 382771 182898 382813 183134
rect 383049 182898 383091 183134
rect 382771 182866 383091 182898
rect 397910 183454 398230 183486
rect 397910 183218 397952 183454
rect 398188 183218 398230 183454
rect 397910 183134 398230 183218
rect 397910 182898 397952 183134
rect 398188 182898 398230 183134
rect 397910 182866 398230 182898
rect 403840 183454 404160 183486
rect 403840 183218 403882 183454
rect 404118 183218 404160 183454
rect 403840 183134 404160 183218
rect 403840 182898 403882 183134
rect 404118 182898 404160 183134
rect 403840 182866 404160 182898
rect 409771 183454 410091 183486
rect 409771 183218 409813 183454
rect 410049 183218 410091 183454
rect 409771 183134 410091 183218
rect 409771 182898 409813 183134
rect 410049 182898 410091 183134
rect 409771 182866 410091 182898
rect 424910 183454 425230 183486
rect 424910 183218 424952 183454
rect 425188 183218 425230 183454
rect 424910 183134 425230 183218
rect 424910 182898 424952 183134
rect 425188 182898 425230 183134
rect 424910 182866 425230 182898
rect 430840 183454 431160 183486
rect 430840 183218 430882 183454
rect 431118 183218 431160 183454
rect 430840 183134 431160 183218
rect 430840 182898 430882 183134
rect 431118 182898 431160 183134
rect 430840 182866 431160 182898
rect 436771 183454 437091 183486
rect 436771 183218 436813 183454
rect 437049 183218 437091 183454
rect 436771 183134 437091 183218
rect 436771 182898 436813 183134
rect 437049 182898 437091 183134
rect 436771 182866 437091 182898
rect 451910 183454 452230 183486
rect 451910 183218 451952 183454
rect 452188 183218 452230 183454
rect 451910 183134 452230 183218
rect 451910 182898 451952 183134
rect 452188 182898 452230 183134
rect 451910 182866 452230 182898
rect 457840 183454 458160 183486
rect 457840 183218 457882 183454
rect 458118 183218 458160 183454
rect 457840 183134 458160 183218
rect 457840 182898 457882 183134
rect 458118 182898 458160 183134
rect 457840 182866 458160 182898
rect 463771 183454 464091 183486
rect 463771 183218 463813 183454
rect 464049 183218 464091 183454
rect 463771 183134 464091 183218
rect 463771 182898 463813 183134
rect 464049 182898 464091 183134
rect 463771 182866 464091 182898
rect 478910 183454 479230 183486
rect 478910 183218 478952 183454
rect 479188 183218 479230 183454
rect 478910 183134 479230 183218
rect 478910 182898 478952 183134
rect 479188 182898 479230 183134
rect 478910 182866 479230 182898
rect 484840 183454 485160 183486
rect 484840 183218 484882 183454
rect 485118 183218 485160 183454
rect 484840 183134 485160 183218
rect 484840 182898 484882 183134
rect 485118 182898 485160 183134
rect 484840 182866 485160 182898
rect 490771 183454 491091 183486
rect 490771 183218 490813 183454
rect 491049 183218 491091 183454
rect 490771 183134 491091 183218
rect 490771 182898 490813 183134
rect 491049 182898 491091 183134
rect 490771 182866 491091 182898
rect 505910 183454 506230 183486
rect 505910 183218 505952 183454
rect 506188 183218 506230 183454
rect 505910 183134 506230 183218
rect 505910 182898 505952 183134
rect 506188 182898 506230 183134
rect 505910 182866 506230 182898
rect 511840 183454 512160 183486
rect 511840 183218 511882 183454
rect 512118 183218 512160 183454
rect 511840 183134 512160 183218
rect 511840 182898 511882 183134
rect 512118 182898 512160 183134
rect 511840 182866 512160 182898
rect 517771 183454 518091 183486
rect 517771 183218 517813 183454
rect 518049 183218 518091 183454
rect 517771 183134 518091 183218
rect 517771 182898 517813 183134
rect 518049 182898 518091 183134
rect 517771 182866 518091 182898
rect 532910 183454 533230 183486
rect 532910 183218 532952 183454
rect 533188 183218 533230 183454
rect 532910 183134 533230 183218
rect 532910 182898 532952 183134
rect 533188 182898 533230 183134
rect 532910 182866 533230 182898
rect 538840 183454 539160 183486
rect 538840 183218 538882 183454
rect 539118 183218 539160 183454
rect 538840 183134 539160 183218
rect 538840 182898 538882 183134
rect 539118 182898 539160 183134
rect 538840 182866 539160 182898
rect 544771 183454 545091 183486
rect 544771 183218 544813 183454
rect 545049 183218 545091 183454
rect 544771 183134 545091 183218
rect 544771 182898 544813 183134
rect 545049 182898 545091 183134
rect 544771 182866 545091 182898
rect 559794 183454 560414 200898
rect 559794 183218 559826 183454
rect 560062 183218 560146 183454
rect 560382 183218 560414 183454
rect 559794 183134 560414 183218
rect 559794 182898 559826 183134
rect 560062 182898 560146 183134
rect 560382 182898 560414 183134
rect 10794 174218 10826 174454
rect 11062 174218 11146 174454
rect 11382 174218 11414 174454
rect 10794 174134 11414 174218
rect 10794 173898 10826 174134
rect 11062 173898 11146 174134
rect 11382 173898 11414 174134
rect 10794 156454 11414 173898
rect 19794 175394 20414 176000
rect 19794 175158 19826 175394
rect 20062 175158 20146 175394
rect 20382 175158 20414 175394
rect 19794 175074 20414 175158
rect 19794 174838 19826 175074
rect 20062 174838 20146 175074
rect 20382 174838 20414 175074
rect 19794 173000 20414 174838
rect 28794 174454 29414 176000
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 173000 29414 173898
rect 37794 175394 38414 176000
rect 37794 175158 37826 175394
rect 38062 175158 38146 175394
rect 38382 175158 38414 175394
rect 37794 175074 38414 175158
rect 37794 174838 37826 175074
rect 38062 174838 38146 175074
rect 38382 174838 38414 175074
rect 37794 173000 38414 174838
rect 46794 174454 47414 176000
rect 46794 174218 46826 174454
rect 47062 174218 47146 174454
rect 47382 174218 47414 174454
rect 46794 174134 47414 174218
rect 46794 173898 46826 174134
rect 47062 173898 47146 174134
rect 47382 173898 47414 174134
rect 46794 173000 47414 173898
rect 55794 175394 56414 176000
rect 55794 175158 55826 175394
rect 56062 175158 56146 175394
rect 56382 175158 56414 175394
rect 55794 175074 56414 175158
rect 55794 174838 55826 175074
rect 56062 174838 56146 175074
rect 56382 174838 56414 175074
rect 55794 173000 56414 174838
rect 64794 174454 65414 176000
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 173000 65414 173898
rect 73794 175394 74414 176000
rect 73794 175158 73826 175394
rect 74062 175158 74146 175394
rect 74382 175158 74414 175394
rect 73794 175074 74414 175158
rect 73794 174838 73826 175074
rect 74062 174838 74146 175074
rect 74382 174838 74414 175074
rect 73794 173000 74414 174838
rect 82794 174454 83414 176000
rect 82794 174218 82826 174454
rect 83062 174218 83146 174454
rect 83382 174218 83414 174454
rect 82794 174134 83414 174218
rect 82794 173898 82826 174134
rect 83062 173898 83146 174134
rect 83382 173898 83414 174134
rect 82794 173000 83414 173898
rect 91794 175394 92414 176000
rect 91794 175158 91826 175394
rect 92062 175158 92146 175394
rect 92382 175158 92414 175394
rect 91794 175074 92414 175158
rect 91794 174838 91826 175074
rect 92062 174838 92146 175074
rect 92382 174838 92414 175074
rect 91794 173000 92414 174838
rect 100794 174454 101414 176000
rect 100794 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 101414 174454
rect 100794 174134 101414 174218
rect 100794 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 101414 174134
rect 100794 173000 101414 173898
rect 109794 175394 110414 176000
rect 109794 175158 109826 175394
rect 110062 175158 110146 175394
rect 110382 175158 110414 175394
rect 109794 175074 110414 175158
rect 109794 174838 109826 175074
rect 110062 174838 110146 175074
rect 110382 174838 110414 175074
rect 109794 173000 110414 174838
rect 118794 174454 119414 176000
rect 118794 174218 118826 174454
rect 119062 174218 119146 174454
rect 119382 174218 119414 174454
rect 118794 174134 119414 174218
rect 118794 173898 118826 174134
rect 119062 173898 119146 174134
rect 119382 173898 119414 174134
rect 118794 173000 119414 173898
rect 127794 175394 128414 176000
rect 127794 175158 127826 175394
rect 128062 175158 128146 175394
rect 128382 175158 128414 175394
rect 127794 175074 128414 175158
rect 127794 174838 127826 175074
rect 128062 174838 128146 175074
rect 128382 174838 128414 175074
rect 127794 173000 128414 174838
rect 136794 174454 137414 176000
rect 136794 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 137414 174454
rect 136794 174134 137414 174218
rect 136794 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 137414 174134
rect 136794 173000 137414 173898
rect 145794 175394 146414 176000
rect 145794 175158 145826 175394
rect 146062 175158 146146 175394
rect 146382 175158 146414 175394
rect 145794 175074 146414 175158
rect 145794 174838 145826 175074
rect 146062 174838 146146 175074
rect 146382 174838 146414 175074
rect 145794 173000 146414 174838
rect 154794 174454 155414 176000
rect 154794 174218 154826 174454
rect 155062 174218 155146 174454
rect 155382 174218 155414 174454
rect 154794 174134 155414 174218
rect 154794 173898 154826 174134
rect 155062 173898 155146 174134
rect 155382 173898 155414 174134
rect 154794 173000 155414 173898
rect 163794 175394 164414 176000
rect 163794 175158 163826 175394
rect 164062 175158 164146 175394
rect 164382 175158 164414 175394
rect 163794 175074 164414 175158
rect 163794 174838 163826 175074
rect 164062 174838 164146 175074
rect 164382 174838 164414 175074
rect 163794 173000 164414 174838
rect 172794 174454 173414 176000
rect 172794 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 173414 174454
rect 172794 174134 173414 174218
rect 172794 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 173414 174134
rect 172794 173000 173414 173898
rect 181794 175394 182414 176000
rect 181794 175158 181826 175394
rect 182062 175158 182146 175394
rect 182382 175158 182414 175394
rect 181794 175074 182414 175158
rect 181794 174838 181826 175074
rect 182062 174838 182146 175074
rect 182382 174838 182414 175074
rect 181794 173000 182414 174838
rect 190794 174454 191414 176000
rect 190794 174218 190826 174454
rect 191062 174218 191146 174454
rect 191382 174218 191414 174454
rect 190794 174134 191414 174218
rect 190794 173898 190826 174134
rect 191062 173898 191146 174134
rect 191382 173898 191414 174134
rect 190794 173000 191414 173898
rect 199794 175394 200414 176000
rect 199794 175158 199826 175394
rect 200062 175158 200146 175394
rect 200382 175158 200414 175394
rect 199794 175074 200414 175158
rect 199794 174838 199826 175074
rect 200062 174838 200146 175074
rect 200382 174838 200414 175074
rect 199794 173000 200414 174838
rect 208794 174454 209414 176000
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 173000 209414 173898
rect 217794 175394 218414 176000
rect 217794 175158 217826 175394
rect 218062 175158 218146 175394
rect 218382 175158 218414 175394
rect 217794 175074 218414 175158
rect 217794 174838 217826 175074
rect 218062 174838 218146 175074
rect 218382 174838 218414 175074
rect 217794 173000 218414 174838
rect 226794 174454 227414 176000
rect 226794 174218 226826 174454
rect 227062 174218 227146 174454
rect 227382 174218 227414 174454
rect 226794 174134 227414 174218
rect 226794 173898 226826 174134
rect 227062 173898 227146 174134
rect 227382 173898 227414 174134
rect 226794 173000 227414 173898
rect 235794 175394 236414 176000
rect 235794 175158 235826 175394
rect 236062 175158 236146 175394
rect 236382 175158 236414 175394
rect 235794 175074 236414 175158
rect 235794 174838 235826 175074
rect 236062 174838 236146 175074
rect 236382 174838 236414 175074
rect 235794 173000 236414 174838
rect 244794 174454 245414 176000
rect 244794 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 245414 174454
rect 244794 174134 245414 174218
rect 244794 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 245414 174134
rect 244794 173000 245414 173898
rect 253794 175394 254414 176000
rect 253794 175158 253826 175394
rect 254062 175158 254146 175394
rect 254382 175158 254414 175394
rect 253794 175074 254414 175158
rect 253794 174838 253826 175074
rect 254062 174838 254146 175074
rect 254382 174838 254414 175074
rect 253794 173000 254414 174838
rect 262794 174454 263414 176000
rect 262794 174218 262826 174454
rect 263062 174218 263146 174454
rect 263382 174218 263414 174454
rect 262794 174134 263414 174218
rect 262794 173898 262826 174134
rect 263062 173898 263146 174134
rect 263382 173898 263414 174134
rect 262794 173000 263414 173898
rect 271794 175394 272414 176000
rect 271794 175158 271826 175394
rect 272062 175158 272146 175394
rect 272382 175158 272414 175394
rect 271794 175074 272414 175158
rect 271794 174838 271826 175074
rect 272062 174838 272146 175074
rect 272382 174838 272414 175074
rect 271794 173000 272414 174838
rect 280794 174454 281414 176000
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 173000 281414 173898
rect 289794 175394 290414 176000
rect 289794 175158 289826 175394
rect 290062 175158 290146 175394
rect 290382 175158 290414 175394
rect 289794 175074 290414 175158
rect 289794 174838 289826 175074
rect 290062 174838 290146 175074
rect 290382 174838 290414 175074
rect 289794 173000 290414 174838
rect 298794 174454 299414 176000
rect 298794 174218 298826 174454
rect 299062 174218 299146 174454
rect 299382 174218 299414 174454
rect 298794 174134 299414 174218
rect 298794 173898 298826 174134
rect 299062 173898 299146 174134
rect 299382 173898 299414 174134
rect 298794 173000 299414 173898
rect 307794 175394 308414 176000
rect 307794 175158 307826 175394
rect 308062 175158 308146 175394
rect 308382 175158 308414 175394
rect 307794 175074 308414 175158
rect 307794 174838 307826 175074
rect 308062 174838 308146 175074
rect 308382 174838 308414 175074
rect 307794 173000 308414 174838
rect 316794 174454 317414 176000
rect 316794 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 317414 174454
rect 316794 174134 317414 174218
rect 316794 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 317414 174134
rect 316794 173000 317414 173898
rect 325794 175394 326414 176000
rect 325794 175158 325826 175394
rect 326062 175158 326146 175394
rect 326382 175158 326414 175394
rect 325794 175074 326414 175158
rect 325794 174838 325826 175074
rect 326062 174838 326146 175074
rect 326382 174838 326414 175074
rect 325794 173000 326414 174838
rect 334794 174454 335414 176000
rect 334794 174218 334826 174454
rect 335062 174218 335146 174454
rect 335382 174218 335414 174454
rect 334794 174134 335414 174218
rect 334794 173898 334826 174134
rect 335062 173898 335146 174134
rect 335382 173898 335414 174134
rect 334794 173000 335414 173898
rect 343794 175394 344414 176000
rect 343794 175158 343826 175394
rect 344062 175158 344146 175394
rect 344382 175158 344414 175394
rect 343794 175074 344414 175158
rect 343794 174838 343826 175074
rect 344062 174838 344146 175074
rect 344382 174838 344414 175074
rect 343794 173000 344414 174838
rect 352794 174454 353414 176000
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 352794 173000 353414 173898
rect 361794 175394 362414 176000
rect 361794 175158 361826 175394
rect 362062 175158 362146 175394
rect 362382 175158 362414 175394
rect 361794 175074 362414 175158
rect 361794 174838 361826 175074
rect 362062 174838 362146 175074
rect 362382 174838 362414 175074
rect 361794 173000 362414 174838
rect 370794 174454 371414 176000
rect 370794 174218 370826 174454
rect 371062 174218 371146 174454
rect 371382 174218 371414 174454
rect 370794 174134 371414 174218
rect 370794 173898 370826 174134
rect 371062 173898 371146 174134
rect 371382 173898 371414 174134
rect 370794 173000 371414 173898
rect 379794 175394 380414 176000
rect 379794 175158 379826 175394
rect 380062 175158 380146 175394
rect 380382 175158 380414 175394
rect 379794 175074 380414 175158
rect 379794 174838 379826 175074
rect 380062 174838 380146 175074
rect 380382 174838 380414 175074
rect 379794 173000 380414 174838
rect 388794 174454 389414 176000
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 173000 389414 173898
rect 397794 175394 398414 176000
rect 397794 175158 397826 175394
rect 398062 175158 398146 175394
rect 398382 175158 398414 175394
rect 397794 175074 398414 175158
rect 397794 174838 397826 175074
rect 398062 174838 398146 175074
rect 398382 174838 398414 175074
rect 397794 173000 398414 174838
rect 406794 174454 407414 176000
rect 406794 174218 406826 174454
rect 407062 174218 407146 174454
rect 407382 174218 407414 174454
rect 406794 174134 407414 174218
rect 406794 173898 406826 174134
rect 407062 173898 407146 174134
rect 407382 173898 407414 174134
rect 406794 173000 407414 173898
rect 415794 175394 416414 176000
rect 415794 175158 415826 175394
rect 416062 175158 416146 175394
rect 416382 175158 416414 175394
rect 415794 175074 416414 175158
rect 415794 174838 415826 175074
rect 416062 174838 416146 175074
rect 416382 174838 416414 175074
rect 415794 173000 416414 174838
rect 424794 174454 425414 176000
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 173000 425414 173898
rect 433794 175394 434414 176000
rect 433794 175158 433826 175394
rect 434062 175158 434146 175394
rect 434382 175158 434414 175394
rect 433794 175074 434414 175158
rect 433794 174838 433826 175074
rect 434062 174838 434146 175074
rect 434382 174838 434414 175074
rect 433794 173000 434414 174838
rect 442794 174454 443414 176000
rect 442794 174218 442826 174454
rect 443062 174218 443146 174454
rect 443382 174218 443414 174454
rect 442794 174134 443414 174218
rect 442794 173898 442826 174134
rect 443062 173898 443146 174134
rect 443382 173898 443414 174134
rect 442794 173000 443414 173898
rect 451794 175394 452414 176000
rect 451794 175158 451826 175394
rect 452062 175158 452146 175394
rect 452382 175158 452414 175394
rect 451794 175074 452414 175158
rect 451794 174838 451826 175074
rect 452062 174838 452146 175074
rect 452382 174838 452414 175074
rect 451794 173000 452414 174838
rect 460794 174454 461414 176000
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 173000 461414 173898
rect 469794 175394 470414 176000
rect 469794 175158 469826 175394
rect 470062 175158 470146 175394
rect 470382 175158 470414 175394
rect 469794 175074 470414 175158
rect 469794 174838 469826 175074
rect 470062 174838 470146 175074
rect 470382 174838 470414 175074
rect 469794 173000 470414 174838
rect 478794 174454 479414 176000
rect 478794 174218 478826 174454
rect 479062 174218 479146 174454
rect 479382 174218 479414 174454
rect 478794 174134 479414 174218
rect 478794 173898 478826 174134
rect 479062 173898 479146 174134
rect 479382 173898 479414 174134
rect 478794 173000 479414 173898
rect 487794 175394 488414 176000
rect 487794 175158 487826 175394
rect 488062 175158 488146 175394
rect 488382 175158 488414 175394
rect 487794 175074 488414 175158
rect 487794 174838 487826 175074
rect 488062 174838 488146 175074
rect 488382 174838 488414 175074
rect 487794 173000 488414 174838
rect 496794 174454 497414 176000
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 173000 497414 173898
rect 505794 175394 506414 176000
rect 505794 175158 505826 175394
rect 506062 175158 506146 175394
rect 506382 175158 506414 175394
rect 505794 175074 506414 175158
rect 505794 174838 505826 175074
rect 506062 174838 506146 175074
rect 506382 174838 506414 175074
rect 505794 173000 506414 174838
rect 514794 174454 515414 176000
rect 514794 174218 514826 174454
rect 515062 174218 515146 174454
rect 515382 174218 515414 174454
rect 514794 174134 515414 174218
rect 514794 173898 514826 174134
rect 515062 173898 515146 174134
rect 515382 173898 515414 174134
rect 514794 173000 515414 173898
rect 523794 175394 524414 176000
rect 523794 175158 523826 175394
rect 524062 175158 524146 175394
rect 524382 175158 524414 175394
rect 523794 175074 524414 175158
rect 523794 174838 523826 175074
rect 524062 174838 524146 175074
rect 524382 174838 524414 175074
rect 523794 173000 524414 174838
rect 532794 174454 533414 176000
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 173000 533414 173898
rect 541794 175394 542414 176000
rect 541794 175158 541826 175394
rect 542062 175158 542146 175394
rect 542382 175158 542414 175394
rect 541794 175074 542414 175158
rect 541794 174838 541826 175074
rect 542062 174838 542146 175074
rect 542382 174838 542414 175074
rect 541794 173000 542414 174838
rect 550794 174454 551414 176000
rect 550794 174218 550826 174454
rect 551062 174218 551146 174454
rect 551382 174218 551414 174454
rect 550794 174134 551414 174218
rect 550794 173898 550826 174134
rect 551062 173898 551146 174134
rect 551382 173898 551414 174134
rect 550794 173000 551414 173898
rect 19910 165454 20230 165486
rect 19910 165218 19952 165454
rect 20188 165218 20230 165454
rect 19910 165134 20230 165218
rect 19910 164898 19952 165134
rect 20188 164898 20230 165134
rect 19910 164866 20230 164898
rect 25840 165454 26160 165486
rect 25840 165218 25882 165454
rect 26118 165218 26160 165454
rect 25840 165134 26160 165218
rect 25840 164898 25882 165134
rect 26118 164898 26160 165134
rect 25840 164866 26160 164898
rect 31771 165454 32091 165486
rect 31771 165218 31813 165454
rect 32049 165218 32091 165454
rect 31771 165134 32091 165218
rect 31771 164898 31813 165134
rect 32049 164898 32091 165134
rect 31771 164866 32091 164898
rect 46910 165454 47230 165486
rect 46910 165218 46952 165454
rect 47188 165218 47230 165454
rect 46910 165134 47230 165218
rect 46910 164898 46952 165134
rect 47188 164898 47230 165134
rect 46910 164866 47230 164898
rect 52840 165454 53160 165486
rect 52840 165218 52882 165454
rect 53118 165218 53160 165454
rect 52840 165134 53160 165218
rect 52840 164898 52882 165134
rect 53118 164898 53160 165134
rect 52840 164866 53160 164898
rect 58771 165454 59091 165486
rect 58771 165218 58813 165454
rect 59049 165218 59091 165454
rect 58771 165134 59091 165218
rect 58771 164898 58813 165134
rect 59049 164898 59091 165134
rect 58771 164866 59091 164898
rect 73910 165454 74230 165486
rect 73910 165218 73952 165454
rect 74188 165218 74230 165454
rect 73910 165134 74230 165218
rect 73910 164898 73952 165134
rect 74188 164898 74230 165134
rect 73910 164866 74230 164898
rect 79840 165454 80160 165486
rect 79840 165218 79882 165454
rect 80118 165218 80160 165454
rect 79840 165134 80160 165218
rect 79840 164898 79882 165134
rect 80118 164898 80160 165134
rect 79840 164866 80160 164898
rect 85771 165454 86091 165486
rect 85771 165218 85813 165454
rect 86049 165218 86091 165454
rect 85771 165134 86091 165218
rect 85771 164898 85813 165134
rect 86049 164898 86091 165134
rect 85771 164866 86091 164898
rect 100910 165454 101230 165486
rect 100910 165218 100952 165454
rect 101188 165218 101230 165454
rect 100910 165134 101230 165218
rect 100910 164898 100952 165134
rect 101188 164898 101230 165134
rect 100910 164866 101230 164898
rect 106840 165454 107160 165486
rect 106840 165218 106882 165454
rect 107118 165218 107160 165454
rect 106840 165134 107160 165218
rect 106840 164898 106882 165134
rect 107118 164898 107160 165134
rect 106840 164866 107160 164898
rect 112771 165454 113091 165486
rect 112771 165218 112813 165454
rect 113049 165218 113091 165454
rect 112771 165134 113091 165218
rect 112771 164898 112813 165134
rect 113049 164898 113091 165134
rect 112771 164866 113091 164898
rect 127910 165454 128230 165486
rect 127910 165218 127952 165454
rect 128188 165218 128230 165454
rect 127910 165134 128230 165218
rect 127910 164898 127952 165134
rect 128188 164898 128230 165134
rect 127910 164866 128230 164898
rect 133840 165454 134160 165486
rect 133840 165218 133882 165454
rect 134118 165218 134160 165454
rect 133840 165134 134160 165218
rect 133840 164898 133882 165134
rect 134118 164898 134160 165134
rect 133840 164866 134160 164898
rect 139771 165454 140091 165486
rect 139771 165218 139813 165454
rect 140049 165218 140091 165454
rect 139771 165134 140091 165218
rect 139771 164898 139813 165134
rect 140049 164898 140091 165134
rect 139771 164866 140091 164898
rect 154910 165454 155230 165486
rect 154910 165218 154952 165454
rect 155188 165218 155230 165454
rect 154910 165134 155230 165218
rect 154910 164898 154952 165134
rect 155188 164898 155230 165134
rect 154910 164866 155230 164898
rect 160840 165454 161160 165486
rect 160840 165218 160882 165454
rect 161118 165218 161160 165454
rect 160840 165134 161160 165218
rect 160840 164898 160882 165134
rect 161118 164898 161160 165134
rect 160840 164866 161160 164898
rect 166771 165454 167091 165486
rect 166771 165218 166813 165454
rect 167049 165218 167091 165454
rect 166771 165134 167091 165218
rect 166771 164898 166813 165134
rect 167049 164898 167091 165134
rect 166771 164866 167091 164898
rect 181910 165454 182230 165486
rect 181910 165218 181952 165454
rect 182188 165218 182230 165454
rect 181910 165134 182230 165218
rect 181910 164898 181952 165134
rect 182188 164898 182230 165134
rect 181910 164866 182230 164898
rect 187840 165454 188160 165486
rect 187840 165218 187882 165454
rect 188118 165218 188160 165454
rect 187840 165134 188160 165218
rect 187840 164898 187882 165134
rect 188118 164898 188160 165134
rect 187840 164866 188160 164898
rect 193771 165454 194091 165486
rect 193771 165218 193813 165454
rect 194049 165218 194091 165454
rect 193771 165134 194091 165218
rect 193771 164898 193813 165134
rect 194049 164898 194091 165134
rect 193771 164866 194091 164898
rect 208910 165454 209230 165486
rect 208910 165218 208952 165454
rect 209188 165218 209230 165454
rect 208910 165134 209230 165218
rect 208910 164898 208952 165134
rect 209188 164898 209230 165134
rect 208910 164866 209230 164898
rect 214840 165454 215160 165486
rect 214840 165218 214882 165454
rect 215118 165218 215160 165454
rect 214840 165134 215160 165218
rect 214840 164898 214882 165134
rect 215118 164898 215160 165134
rect 214840 164866 215160 164898
rect 220771 165454 221091 165486
rect 220771 165218 220813 165454
rect 221049 165218 221091 165454
rect 220771 165134 221091 165218
rect 220771 164898 220813 165134
rect 221049 164898 221091 165134
rect 220771 164866 221091 164898
rect 235910 165454 236230 165486
rect 235910 165218 235952 165454
rect 236188 165218 236230 165454
rect 235910 165134 236230 165218
rect 235910 164898 235952 165134
rect 236188 164898 236230 165134
rect 235910 164866 236230 164898
rect 241840 165454 242160 165486
rect 241840 165218 241882 165454
rect 242118 165218 242160 165454
rect 241840 165134 242160 165218
rect 241840 164898 241882 165134
rect 242118 164898 242160 165134
rect 241840 164866 242160 164898
rect 247771 165454 248091 165486
rect 247771 165218 247813 165454
rect 248049 165218 248091 165454
rect 247771 165134 248091 165218
rect 247771 164898 247813 165134
rect 248049 164898 248091 165134
rect 247771 164866 248091 164898
rect 262910 165454 263230 165486
rect 262910 165218 262952 165454
rect 263188 165218 263230 165454
rect 262910 165134 263230 165218
rect 262910 164898 262952 165134
rect 263188 164898 263230 165134
rect 262910 164866 263230 164898
rect 268840 165454 269160 165486
rect 268840 165218 268882 165454
rect 269118 165218 269160 165454
rect 268840 165134 269160 165218
rect 268840 164898 268882 165134
rect 269118 164898 269160 165134
rect 268840 164866 269160 164898
rect 274771 165454 275091 165486
rect 274771 165218 274813 165454
rect 275049 165218 275091 165454
rect 274771 165134 275091 165218
rect 274771 164898 274813 165134
rect 275049 164898 275091 165134
rect 274771 164866 275091 164898
rect 289910 165454 290230 165486
rect 289910 165218 289952 165454
rect 290188 165218 290230 165454
rect 289910 165134 290230 165218
rect 289910 164898 289952 165134
rect 290188 164898 290230 165134
rect 289910 164866 290230 164898
rect 295840 165454 296160 165486
rect 295840 165218 295882 165454
rect 296118 165218 296160 165454
rect 295840 165134 296160 165218
rect 295840 164898 295882 165134
rect 296118 164898 296160 165134
rect 295840 164866 296160 164898
rect 301771 165454 302091 165486
rect 301771 165218 301813 165454
rect 302049 165218 302091 165454
rect 301771 165134 302091 165218
rect 301771 164898 301813 165134
rect 302049 164898 302091 165134
rect 301771 164866 302091 164898
rect 316910 165454 317230 165486
rect 316910 165218 316952 165454
rect 317188 165218 317230 165454
rect 316910 165134 317230 165218
rect 316910 164898 316952 165134
rect 317188 164898 317230 165134
rect 316910 164866 317230 164898
rect 322840 165454 323160 165486
rect 322840 165218 322882 165454
rect 323118 165218 323160 165454
rect 322840 165134 323160 165218
rect 322840 164898 322882 165134
rect 323118 164898 323160 165134
rect 322840 164866 323160 164898
rect 328771 165454 329091 165486
rect 328771 165218 328813 165454
rect 329049 165218 329091 165454
rect 328771 165134 329091 165218
rect 328771 164898 328813 165134
rect 329049 164898 329091 165134
rect 328771 164866 329091 164898
rect 343910 165454 344230 165486
rect 343910 165218 343952 165454
rect 344188 165218 344230 165454
rect 343910 165134 344230 165218
rect 343910 164898 343952 165134
rect 344188 164898 344230 165134
rect 343910 164866 344230 164898
rect 349840 165454 350160 165486
rect 349840 165218 349882 165454
rect 350118 165218 350160 165454
rect 349840 165134 350160 165218
rect 349840 164898 349882 165134
rect 350118 164898 350160 165134
rect 349840 164866 350160 164898
rect 355771 165454 356091 165486
rect 355771 165218 355813 165454
rect 356049 165218 356091 165454
rect 355771 165134 356091 165218
rect 355771 164898 355813 165134
rect 356049 164898 356091 165134
rect 355771 164866 356091 164898
rect 370910 165454 371230 165486
rect 370910 165218 370952 165454
rect 371188 165218 371230 165454
rect 370910 165134 371230 165218
rect 370910 164898 370952 165134
rect 371188 164898 371230 165134
rect 370910 164866 371230 164898
rect 376840 165454 377160 165486
rect 376840 165218 376882 165454
rect 377118 165218 377160 165454
rect 376840 165134 377160 165218
rect 376840 164898 376882 165134
rect 377118 164898 377160 165134
rect 376840 164866 377160 164898
rect 382771 165454 383091 165486
rect 382771 165218 382813 165454
rect 383049 165218 383091 165454
rect 382771 165134 383091 165218
rect 382771 164898 382813 165134
rect 383049 164898 383091 165134
rect 382771 164866 383091 164898
rect 397910 165454 398230 165486
rect 397910 165218 397952 165454
rect 398188 165218 398230 165454
rect 397910 165134 398230 165218
rect 397910 164898 397952 165134
rect 398188 164898 398230 165134
rect 397910 164866 398230 164898
rect 403840 165454 404160 165486
rect 403840 165218 403882 165454
rect 404118 165218 404160 165454
rect 403840 165134 404160 165218
rect 403840 164898 403882 165134
rect 404118 164898 404160 165134
rect 403840 164866 404160 164898
rect 409771 165454 410091 165486
rect 409771 165218 409813 165454
rect 410049 165218 410091 165454
rect 409771 165134 410091 165218
rect 409771 164898 409813 165134
rect 410049 164898 410091 165134
rect 409771 164866 410091 164898
rect 424910 165454 425230 165486
rect 424910 165218 424952 165454
rect 425188 165218 425230 165454
rect 424910 165134 425230 165218
rect 424910 164898 424952 165134
rect 425188 164898 425230 165134
rect 424910 164866 425230 164898
rect 430840 165454 431160 165486
rect 430840 165218 430882 165454
rect 431118 165218 431160 165454
rect 430840 165134 431160 165218
rect 430840 164898 430882 165134
rect 431118 164898 431160 165134
rect 430840 164866 431160 164898
rect 436771 165454 437091 165486
rect 436771 165218 436813 165454
rect 437049 165218 437091 165454
rect 436771 165134 437091 165218
rect 436771 164898 436813 165134
rect 437049 164898 437091 165134
rect 436771 164866 437091 164898
rect 451910 165454 452230 165486
rect 451910 165218 451952 165454
rect 452188 165218 452230 165454
rect 451910 165134 452230 165218
rect 451910 164898 451952 165134
rect 452188 164898 452230 165134
rect 451910 164866 452230 164898
rect 457840 165454 458160 165486
rect 457840 165218 457882 165454
rect 458118 165218 458160 165454
rect 457840 165134 458160 165218
rect 457840 164898 457882 165134
rect 458118 164898 458160 165134
rect 457840 164866 458160 164898
rect 463771 165454 464091 165486
rect 463771 165218 463813 165454
rect 464049 165218 464091 165454
rect 463771 165134 464091 165218
rect 463771 164898 463813 165134
rect 464049 164898 464091 165134
rect 463771 164866 464091 164898
rect 478910 165454 479230 165486
rect 478910 165218 478952 165454
rect 479188 165218 479230 165454
rect 478910 165134 479230 165218
rect 478910 164898 478952 165134
rect 479188 164898 479230 165134
rect 478910 164866 479230 164898
rect 484840 165454 485160 165486
rect 484840 165218 484882 165454
rect 485118 165218 485160 165454
rect 484840 165134 485160 165218
rect 484840 164898 484882 165134
rect 485118 164898 485160 165134
rect 484840 164866 485160 164898
rect 490771 165454 491091 165486
rect 490771 165218 490813 165454
rect 491049 165218 491091 165454
rect 490771 165134 491091 165218
rect 490771 164898 490813 165134
rect 491049 164898 491091 165134
rect 490771 164866 491091 164898
rect 505910 165454 506230 165486
rect 505910 165218 505952 165454
rect 506188 165218 506230 165454
rect 505910 165134 506230 165218
rect 505910 164898 505952 165134
rect 506188 164898 506230 165134
rect 505910 164866 506230 164898
rect 511840 165454 512160 165486
rect 511840 165218 511882 165454
rect 512118 165218 512160 165454
rect 511840 165134 512160 165218
rect 511840 164898 511882 165134
rect 512118 164898 512160 165134
rect 511840 164866 512160 164898
rect 517771 165454 518091 165486
rect 517771 165218 517813 165454
rect 518049 165218 518091 165454
rect 517771 165134 518091 165218
rect 517771 164898 517813 165134
rect 518049 164898 518091 165134
rect 517771 164866 518091 164898
rect 532910 165454 533230 165486
rect 532910 165218 532952 165454
rect 533188 165218 533230 165454
rect 532910 165134 533230 165218
rect 532910 164898 532952 165134
rect 533188 164898 533230 165134
rect 532910 164866 533230 164898
rect 538840 165454 539160 165486
rect 538840 165218 538882 165454
rect 539118 165218 539160 165454
rect 538840 165134 539160 165218
rect 538840 164898 538882 165134
rect 539118 164898 539160 165134
rect 538840 164866 539160 164898
rect 544771 165454 545091 165486
rect 544771 165218 544813 165454
rect 545049 165218 545091 165454
rect 544771 165134 545091 165218
rect 544771 164898 544813 165134
rect 545049 164898 545091 165134
rect 544771 164866 545091 164898
rect 559794 165454 560414 182898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 138454 11414 155898
rect 22874 156454 23194 156486
rect 22874 156218 22916 156454
rect 23152 156218 23194 156454
rect 22874 156134 23194 156218
rect 22874 155898 22916 156134
rect 23152 155898 23194 156134
rect 22874 155866 23194 155898
rect 28805 156454 29125 156486
rect 28805 156218 28847 156454
rect 29083 156218 29125 156454
rect 28805 156134 29125 156218
rect 28805 155898 28847 156134
rect 29083 155898 29125 156134
rect 28805 155866 29125 155898
rect 49874 156454 50194 156486
rect 49874 156218 49916 156454
rect 50152 156218 50194 156454
rect 49874 156134 50194 156218
rect 49874 155898 49916 156134
rect 50152 155898 50194 156134
rect 49874 155866 50194 155898
rect 55805 156454 56125 156486
rect 55805 156218 55847 156454
rect 56083 156218 56125 156454
rect 55805 156134 56125 156218
rect 55805 155898 55847 156134
rect 56083 155898 56125 156134
rect 55805 155866 56125 155898
rect 76874 156454 77194 156486
rect 76874 156218 76916 156454
rect 77152 156218 77194 156454
rect 76874 156134 77194 156218
rect 76874 155898 76916 156134
rect 77152 155898 77194 156134
rect 76874 155866 77194 155898
rect 82805 156454 83125 156486
rect 82805 156218 82847 156454
rect 83083 156218 83125 156454
rect 82805 156134 83125 156218
rect 82805 155898 82847 156134
rect 83083 155898 83125 156134
rect 82805 155866 83125 155898
rect 103874 156454 104194 156486
rect 103874 156218 103916 156454
rect 104152 156218 104194 156454
rect 103874 156134 104194 156218
rect 103874 155898 103916 156134
rect 104152 155898 104194 156134
rect 103874 155866 104194 155898
rect 109805 156454 110125 156486
rect 109805 156218 109847 156454
rect 110083 156218 110125 156454
rect 109805 156134 110125 156218
rect 109805 155898 109847 156134
rect 110083 155898 110125 156134
rect 109805 155866 110125 155898
rect 130874 156454 131194 156486
rect 130874 156218 130916 156454
rect 131152 156218 131194 156454
rect 130874 156134 131194 156218
rect 130874 155898 130916 156134
rect 131152 155898 131194 156134
rect 130874 155866 131194 155898
rect 136805 156454 137125 156486
rect 136805 156218 136847 156454
rect 137083 156218 137125 156454
rect 136805 156134 137125 156218
rect 136805 155898 136847 156134
rect 137083 155898 137125 156134
rect 136805 155866 137125 155898
rect 157874 156454 158194 156486
rect 157874 156218 157916 156454
rect 158152 156218 158194 156454
rect 157874 156134 158194 156218
rect 157874 155898 157916 156134
rect 158152 155898 158194 156134
rect 157874 155866 158194 155898
rect 163805 156454 164125 156486
rect 163805 156218 163847 156454
rect 164083 156218 164125 156454
rect 163805 156134 164125 156218
rect 163805 155898 163847 156134
rect 164083 155898 164125 156134
rect 163805 155866 164125 155898
rect 184874 156454 185194 156486
rect 184874 156218 184916 156454
rect 185152 156218 185194 156454
rect 184874 156134 185194 156218
rect 184874 155898 184916 156134
rect 185152 155898 185194 156134
rect 184874 155866 185194 155898
rect 190805 156454 191125 156486
rect 190805 156218 190847 156454
rect 191083 156218 191125 156454
rect 190805 156134 191125 156218
rect 190805 155898 190847 156134
rect 191083 155898 191125 156134
rect 190805 155866 191125 155898
rect 211874 156454 212194 156486
rect 211874 156218 211916 156454
rect 212152 156218 212194 156454
rect 211874 156134 212194 156218
rect 211874 155898 211916 156134
rect 212152 155898 212194 156134
rect 211874 155866 212194 155898
rect 217805 156454 218125 156486
rect 217805 156218 217847 156454
rect 218083 156218 218125 156454
rect 217805 156134 218125 156218
rect 217805 155898 217847 156134
rect 218083 155898 218125 156134
rect 217805 155866 218125 155898
rect 238874 156454 239194 156486
rect 238874 156218 238916 156454
rect 239152 156218 239194 156454
rect 238874 156134 239194 156218
rect 238874 155898 238916 156134
rect 239152 155898 239194 156134
rect 238874 155866 239194 155898
rect 244805 156454 245125 156486
rect 244805 156218 244847 156454
rect 245083 156218 245125 156454
rect 244805 156134 245125 156218
rect 244805 155898 244847 156134
rect 245083 155898 245125 156134
rect 244805 155866 245125 155898
rect 265874 156454 266194 156486
rect 265874 156218 265916 156454
rect 266152 156218 266194 156454
rect 265874 156134 266194 156218
rect 265874 155898 265916 156134
rect 266152 155898 266194 156134
rect 265874 155866 266194 155898
rect 271805 156454 272125 156486
rect 271805 156218 271847 156454
rect 272083 156218 272125 156454
rect 271805 156134 272125 156218
rect 271805 155898 271847 156134
rect 272083 155898 272125 156134
rect 271805 155866 272125 155898
rect 292874 156454 293194 156486
rect 292874 156218 292916 156454
rect 293152 156218 293194 156454
rect 292874 156134 293194 156218
rect 292874 155898 292916 156134
rect 293152 155898 293194 156134
rect 292874 155866 293194 155898
rect 298805 156454 299125 156486
rect 298805 156218 298847 156454
rect 299083 156218 299125 156454
rect 298805 156134 299125 156218
rect 298805 155898 298847 156134
rect 299083 155898 299125 156134
rect 298805 155866 299125 155898
rect 319874 156454 320194 156486
rect 319874 156218 319916 156454
rect 320152 156218 320194 156454
rect 319874 156134 320194 156218
rect 319874 155898 319916 156134
rect 320152 155898 320194 156134
rect 319874 155866 320194 155898
rect 325805 156454 326125 156486
rect 325805 156218 325847 156454
rect 326083 156218 326125 156454
rect 325805 156134 326125 156218
rect 325805 155898 325847 156134
rect 326083 155898 326125 156134
rect 325805 155866 326125 155898
rect 346874 156454 347194 156486
rect 346874 156218 346916 156454
rect 347152 156218 347194 156454
rect 346874 156134 347194 156218
rect 346874 155898 346916 156134
rect 347152 155898 347194 156134
rect 346874 155866 347194 155898
rect 352805 156454 353125 156486
rect 352805 156218 352847 156454
rect 353083 156218 353125 156454
rect 352805 156134 353125 156218
rect 352805 155898 352847 156134
rect 353083 155898 353125 156134
rect 352805 155866 353125 155898
rect 373874 156454 374194 156486
rect 373874 156218 373916 156454
rect 374152 156218 374194 156454
rect 373874 156134 374194 156218
rect 373874 155898 373916 156134
rect 374152 155898 374194 156134
rect 373874 155866 374194 155898
rect 379805 156454 380125 156486
rect 379805 156218 379847 156454
rect 380083 156218 380125 156454
rect 379805 156134 380125 156218
rect 379805 155898 379847 156134
rect 380083 155898 380125 156134
rect 379805 155866 380125 155898
rect 400874 156454 401194 156486
rect 400874 156218 400916 156454
rect 401152 156218 401194 156454
rect 400874 156134 401194 156218
rect 400874 155898 400916 156134
rect 401152 155898 401194 156134
rect 400874 155866 401194 155898
rect 406805 156454 407125 156486
rect 406805 156218 406847 156454
rect 407083 156218 407125 156454
rect 406805 156134 407125 156218
rect 406805 155898 406847 156134
rect 407083 155898 407125 156134
rect 406805 155866 407125 155898
rect 427874 156454 428194 156486
rect 427874 156218 427916 156454
rect 428152 156218 428194 156454
rect 427874 156134 428194 156218
rect 427874 155898 427916 156134
rect 428152 155898 428194 156134
rect 427874 155866 428194 155898
rect 433805 156454 434125 156486
rect 433805 156218 433847 156454
rect 434083 156218 434125 156454
rect 433805 156134 434125 156218
rect 433805 155898 433847 156134
rect 434083 155898 434125 156134
rect 433805 155866 434125 155898
rect 454874 156454 455194 156486
rect 454874 156218 454916 156454
rect 455152 156218 455194 156454
rect 454874 156134 455194 156218
rect 454874 155898 454916 156134
rect 455152 155898 455194 156134
rect 454874 155866 455194 155898
rect 460805 156454 461125 156486
rect 460805 156218 460847 156454
rect 461083 156218 461125 156454
rect 460805 156134 461125 156218
rect 460805 155898 460847 156134
rect 461083 155898 461125 156134
rect 460805 155866 461125 155898
rect 481874 156454 482194 156486
rect 481874 156218 481916 156454
rect 482152 156218 482194 156454
rect 481874 156134 482194 156218
rect 481874 155898 481916 156134
rect 482152 155898 482194 156134
rect 481874 155866 482194 155898
rect 487805 156454 488125 156486
rect 487805 156218 487847 156454
rect 488083 156218 488125 156454
rect 487805 156134 488125 156218
rect 487805 155898 487847 156134
rect 488083 155898 488125 156134
rect 487805 155866 488125 155898
rect 508874 156454 509194 156486
rect 508874 156218 508916 156454
rect 509152 156218 509194 156454
rect 508874 156134 509194 156218
rect 508874 155898 508916 156134
rect 509152 155898 509194 156134
rect 508874 155866 509194 155898
rect 514805 156454 515125 156486
rect 514805 156218 514847 156454
rect 515083 156218 515125 156454
rect 514805 156134 515125 156218
rect 514805 155898 514847 156134
rect 515083 155898 515125 156134
rect 514805 155866 515125 155898
rect 535874 156454 536194 156486
rect 535874 156218 535916 156454
rect 536152 156218 536194 156454
rect 535874 156134 536194 156218
rect 535874 155898 535916 156134
rect 536152 155898 536194 156134
rect 535874 155866 536194 155898
rect 541805 156454 542125 156486
rect 541805 156218 541847 156454
rect 542083 156218 542125 156454
rect 541805 156134 542125 156218
rect 541805 155898 541847 156134
rect 542083 155898 542125 156134
rect 541805 155866 542125 155898
rect 19794 147454 20414 149000
rect 19794 147218 19826 147454
rect 20062 147218 20146 147454
rect 20382 147218 20414 147454
rect 19794 147134 20414 147218
rect 19794 146898 19826 147134
rect 20062 146898 20146 147134
rect 20382 146898 20414 147134
rect 19794 146000 20414 146898
rect 28794 148394 29414 149000
rect 28794 148158 28826 148394
rect 29062 148158 29146 148394
rect 29382 148158 29414 148394
rect 28794 148074 29414 148158
rect 28794 147838 28826 148074
rect 29062 147838 29146 148074
rect 29382 147838 29414 148074
rect 28794 146000 29414 147838
rect 37794 147454 38414 149000
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 146000 38414 146898
rect 46794 148394 47414 149000
rect 46794 148158 46826 148394
rect 47062 148158 47146 148394
rect 47382 148158 47414 148394
rect 46794 148074 47414 148158
rect 46794 147838 46826 148074
rect 47062 147838 47146 148074
rect 47382 147838 47414 148074
rect 46794 146000 47414 147838
rect 55794 147454 56414 149000
rect 55794 147218 55826 147454
rect 56062 147218 56146 147454
rect 56382 147218 56414 147454
rect 55794 147134 56414 147218
rect 55794 146898 55826 147134
rect 56062 146898 56146 147134
rect 56382 146898 56414 147134
rect 55794 146000 56414 146898
rect 64794 148394 65414 149000
rect 64794 148158 64826 148394
rect 65062 148158 65146 148394
rect 65382 148158 65414 148394
rect 64794 148074 65414 148158
rect 64794 147838 64826 148074
rect 65062 147838 65146 148074
rect 65382 147838 65414 148074
rect 64794 146000 65414 147838
rect 73794 147454 74414 149000
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 146000 74414 146898
rect 82794 148394 83414 149000
rect 82794 148158 82826 148394
rect 83062 148158 83146 148394
rect 83382 148158 83414 148394
rect 82794 148074 83414 148158
rect 82794 147838 82826 148074
rect 83062 147838 83146 148074
rect 83382 147838 83414 148074
rect 82794 146000 83414 147838
rect 91794 147454 92414 149000
rect 91794 147218 91826 147454
rect 92062 147218 92146 147454
rect 92382 147218 92414 147454
rect 91794 147134 92414 147218
rect 91794 146898 91826 147134
rect 92062 146898 92146 147134
rect 92382 146898 92414 147134
rect 91794 146000 92414 146898
rect 100794 148394 101414 149000
rect 100794 148158 100826 148394
rect 101062 148158 101146 148394
rect 101382 148158 101414 148394
rect 100794 148074 101414 148158
rect 100794 147838 100826 148074
rect 101062 147838 101146 148074
rect 101382 147838 101414 148074
rect 100794 146000 101414 147838
rect 109794 147454 110414 149000
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 146000 110414 146898
rect 118794 148394 119414 149000
rect 118794 148158 118826 148394
rect 119062 148158 119146 148394
rect 119382 148158 119414 148394
rect 118794 148074 119414 148158
rect 118794 147838 118826 148074
rect 119062 147838 119146 148074
rect 119382 147838 119414 148074
rect 118794 146000 119414 147838
rect 127794 147454 128414 149000
rect 127794 147218 127826 147454
rect 128062 147218 128146 147454
rect 128382 147218 128414 147454
rect 127794 147134 128414 147218
rect 127794 146898 127826 147134
rect 128062 146898 128146 147134
rect 128382 146898 128414 147134
rect 127794 146000 128414 146898
rect 136794 148394 137414 149000
rect 136794 148158 136826 148394
rect 137062 148158 137146 148394
rect 137382 148158 137414 148394
rect 136794 148074 137414 148158
rect 136794 147838 136826 148074
rect 137062 147838 137146 148074
rect 137382 147838 137414 148074
rect 136794 146000 137414 147838
rect 145794 147454 146414 149000
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 146000 146414 146898
rect 154794 148394 155414 149000
rect 154794 148158 154826 148394
rect 155062 148158 155146 148394
rect 155382 148158 155414 148394
rect 154794 148074 155414 148158
rect 154794 147838 154826 148074
rect 155062 147838 155146 148074
rect 155382 147838 155414 148074
rect 154794 146000 155414 147838
rect 163794 147454 164414 149000
rect 163794 147218 163826 147454
rect 164062 147218 164146 147454
rect 164382 147218 164414 147454
rect 163794 147134 164414 147218
rect 163794 146898 163826 147134
rect 164062 146898 164146 147134
rect 164382 146898 164414 147134
rect 163794 146000 164414 146898
rect 172794 148394 173414 149000
rect 172794 148158 172826 148394
rect 173062 148158 173146 148394
rect 173382 148158 173414 148394
rect 172794 148074 173414 148158
rect 172794 147838 172826 148074
rect 173062 147838 173146 148074
rect 173382 147838 173414 148074
rect 172794 146000 173414 147838
rect 181794 147454 182414 149000
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 146000 182414 146898
rect 190794 148394 191414 149000
rect 190794 148158 190826 148394
rect 191062 148158 191146 148394
rect 191382 148158 191414 148394
rect 190794 148074 191414 148158
rect 190794 147838 190826 148074
rect 191062 147838 191146 148074
rect 191382 147838 191414 148074
rect 190794 146000 191414 147838
rect 199794 147454 200414 149000
rect 199794 147218 199826 147454
rect 200062 147218 200146 147454
rect 200382 147218 200414 147454
rect 199794 147134 200414 147218
rect 199794 146898 199826 147134
rect 200062 146898 200146 147134
rect 200382 146898 200414 147134
rect 199794 146000 200414 146898
rect 208794 148394 209414 149000
rect 208794 148158 208826 148394
rect 209062 148158 209146 148394
rect 209382 148158 209414 148394
rect 208794 148074 209414 148158
rect 208794 147838 208826 148074
rect 209062 147838 209146 148074
rect 209382 147838 209414 148074
rect 208794 146000 209414 147838
rect 217794 147454 218414 149000
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 146000 218414 146898
rect 226794 148394 227414 149000
rect 226794 148158 226826 148394
rect 227062 148158 227146 148394
rect 227382 148158 227414 148394
rect 226794 148074 227414 148158
rect 226794 147838 226826 148074
rect 227062 147838 227146 148074
rect 227382 147838 227414 148074
rect 226794 146000 227414 147838
rect 235794 147454 236414 149000
rect 235794 147218 235826 147454
rect 236062 147218 236146 147454
rect 236382 147218 236414 147454
rect 235794 147134 236414 147218
rect 235794 146898 235826 147134
rect 236062 146898 236146 147134
rect 236382 146898 236414 147134
rect 235794 146000 236414 146898
rect 244794 148394 245414 149000
rect 244794 148158 244826 148394
rect 245062 148158 245146 148394
rect 245382 148158 245414 148394
rect 244794 148074 245414 148158
rect 244794 147838 244826 148074
rect 245062 147838 245146 148074
rect 245382 147838 245414 148074
rect 244794 146000 245414 147838
rect 253794 147454 254414 149000
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 146000 254414 146898
rect 262794 148394 263414 149000
rect 262794 148158 262826 148394
rect 263062 148158 263146 148394
rect 263382 148158 263414 148394
rect 262794 148074 263414 148158
rect 262794 147838 262826 148074
rect 263062 147838 263146 148074
rect 263382 147838 263414 148074
rect 262794 146000 263414 147838
rect 271794 147454 272414 149000
rect 271794 147218 271826 147454
rect 272062 147218 272146 147454
rect 272382 147218 272414 147454
rect 271794 147134 272414 147218
rect 271794 146898 271826 147134
rect 272062 146898 272146 147134
rect 272382 146898 272414 147134
rect 271794 146000 272414 146898
rect 280794 148394 281414 149000
rect 280794 148158 280826 148394
rect 281062 148158 281146 148394
rect 281382 148158 281414 148394
rect 280794 148074 281414 148158
rect 280794 147838 280826 148074
rect 281062 147838 281146 148074
rect 281382 147838 281414 148074
rect 280794 146000 281414 147838
rect 289794 147454 290414 149000
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 146000 290414 146898
rect 298794 148394 299414 149000
rect 298794 148158 298826 148394
rect 299062 148158 299146 148394
rect 299382 148158 299414 148394
rect 298794 148074 299414 148158
rect 298794 147838 298826 148074
rect 299062 147838 299146 148074
rect 299382 147838 299414 148074
rect 298794 146000 299414 147838
rect 307794 147454 308414 149000
rect 307794 147218 307826 147454
rect 308062 147218 308146 147454
rect 308382 147218 308414 147454
rect 307794 147134 308414 147218
rect 307794 146898 307826 147134
rect 308062 146898 308146 147134
rect 308382 146898 308414 147134
rect 307794 146000 308414 146898
rect 316794 148394 317414 149000
rect 316794 148158 316826 148394
rect 317062 148158 317146 148394
rect 317382 148158 317414 148394
rect 316794 148074 317414 148158
rect 316794 147838 316826 148074
rect 317062 147838 317146 148074
rect 317382 147838 317414 148074
rect 316794 146000 317414 147838
rect 325794 147454 326414 149000
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 146000 326414 146898
rect 334794 148394 335414 149000
rect 334794 148158 334826 148394
rect 335062 148158 335146 148394
rect 335382 148158 335414 148394
rect 334794 148074 335414 148158
rect 334794 147838 334826 148074
rect 335062 147838 335146 148074
rect 335382 147838 335414 148074
rect 334794 146000 335414 147838
rect 343794 147454 344414 149000
rect 343794 147218 343826 147454
rect 344062 147218 344146 147454
rect 344382 147218 344414 147454
rect 343794 147134 344414 147218
rect 343794 146898 343826 147134
rect 344062 146898 344146 147134
rect 344382 146898 344414 147134
rect 343794 146000 344414 146898
rect 352794 148394 353414 149000
rect 352794 148158 352826 148394
rect 353062 148158 353146 148394
rect 353382 148158 353414 148394
rect 352794 148074 353414 148158
rect 352794 147838 352826 148074
rect 353062 147838 353146 148074
rect 353382 147838 353414 148074
rect 352794 146000 353414 147838
rect 361794 147454 362414 149000
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 146000 362414 146898
rect 370794 148394 371414 149000
rect 370794 148158 370826 148394
rect 371062 148158 371146 148394
rect 371382 148158 371414 148394
rect 370794 148074 371414 148158
rect 370794 147838 370826 148074
rect 371062 147838 371146 148074
rect 371382 147838 371414 148074
rect 370794 146000 371414 147838
rect 379794 147454 380414 149000
rect 379794 147218 379826 147454
rect 380062 147218 380146 147454
rect 380382 147218 380414 147454
rect 379794 147134 380414 147218
rect 379794 146898 379826 147134
rect 380062 146898 380146 147134
rect 380382 146898 380414 147134
rect 379794 146000 380414 146898
rect 388794 148394 389414 149000
rect 388794 148158 388826 148394
rect 389062 148158 389146 148394
rect 389382 148158 389414 148394
rect 388794 148074 389414 148158
rect 388794 147838 388826 148074
rect 389062 147838 389146 148074
rect 389382 147838 389414 148074
rect 388794 146000 389414 147838
rect 397794 147454 398414 149000
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 146000 398414 146898
rect 406794 148394 407414 149000
rect 406794 148158 406826 148394
rect 407062 148158 407146 148394
rect 407382 148158 407414 148394
rect 406794 148074 407414 148158
rect 406794 147838 406826 148074
rect 407062 147838 407146 148074
rect 407382 147838 407414 148074
rect 406794 146000 407414 147838
rect 415794 147454 416414 149000
rect 415794 147218 415826 147454
rect 416062 147218 416146 147454
rect 416382 147218 416414 147454
rect 415794 147134 416414 147218
rect 415794 146898 415826 147134
rect 416062 146898 416146 147134
rect 416382 146898 416414 147134
rect 415794 146000 416414 146898
rect 424794 148394 425414 149000
rect 424794 148158 424826 148394
rect 425062 148158 425146 148394
rect 425382 148158 425414 148394
rect 424794 148074 425414 148158
rect 424794 147838 424826 148074
rect 425062 147838 425146 148074
rect 425382 147838 425414 148074
rect 424794 146000 425414 147838
rect 433794 147454 434414 149000
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 146000 434414 146898
rect 442794 148394 443414 149000
rect 442794 148158 442826 148394
rect 443062 148158 443146 148394
rect 443382 148158 443414 148394
rect 442794 148074 443414 148158
rect 442794 147838 442826 148074
rect 443062 147838 443146 148074
rect 443382 147838 443414 148074
rect 442794 146000 443414 147838
rect 451794 147454 452414 149000
rect 451794 147218 451826 147454
rect 452062 147218 452146 147454
rect 452382 147218 452414 147454
rect 451794 147134 452414 147218
rect 451794 146898 451826 147134
rect 452062 146898 452146 147134
rect 452382 146898 452414 147134
rect 451794 146000 452414 146898
rect 460794 148394 461414 149000
rect 460794 148158 460826 148394
rect 461062 148158 461146 148394
rect 461382 148158 461414 148394
rect 460794 148074 461414 148158
rect 460794 147838 460826 148074
rect 461062 147838 461146 148074
rect 461382 147838 461414 148074
rect 460794 146000 461414 147838
rect 469794 147454 470414 149000
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 146000 470414 146898
rect 478794 148394 479414 149000
rect 478794 148158 478826 148394
rect 479062 148158 479146 148394
rect 479382 148158 479414 148394
rect 478794 148074 479414 148158
rect 478794 147838 478826 148074
rect 479062 147838 479146 148074
rect 479382 147838 479414 148074
rect 478794 146000 479414 147838
rect 487794 147454 488414 149000
rect 487794 147218 487826 147454
rect 488062 147218 488146 147454
rect 488382 147218 488414 147454
rect 487794 147134 488414 147218
rect 487794 146898 487826 147134
rect 488062 146898 488146 147134
rect 488382 146898 488414 147134
rect 487794 146000 488414 146898
rect 496794 148394 497414 149000
rect 496794 148158 496826 148394
rect 497062 148158 497146 148394
rect 497382 148158 497414 148394
rect 496794 148074 497414 148158
rect 496794 147838 496826 148074
rect 497062 147838 497146 148074
rect 497382 147838 497414 148074
rect 496794 146000 497414 147838
rect 505794 147454 506414 149000
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 146000 506414 146898
rect 514794 148394 515414 149000
rect 514794 148158 514826 148394
rect 515062 148158 515146 148394
rect 515382 148158 515414 148394
rect 514794 148074 515414 148158
rect 514794 147838 514826 148074
rect 515062 147838 515146 148074
rect 515382 147838 515414 148074
rect 514794 146000 515414 147838
rect 523794 147454 524414 149000
rect 523794 147218 523826 147454
rect 524062 147218 524146 147454
rect 524382 147218 524414 147454
rect 523794 147134 524414 147218
rect 523794 146898 523826 147134
rect 524062 146898 524146 147134
rect 524382 146898 524414 147134
rect 523794 146000 524414 146898
rect 532794 148394 533414 149000
rect 532794 148158 532826 148394
rect 533062 148158 533146 148394
rect 533382 148158 533414 148394
rect 532794 148074 533414 148158
rect 532794 147838 532826 148074
rect 533062 147838 533146 148074
rect 533382 147838 533414 148074
rect 532794 146000 533414 147838
rect 541794 147454 542414 149000
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 146000 542414 146898
rect 550794 148394 551414 149000
rect 550794 148158 550826 148394
rect 551062 148158 551146 148394
rect 551382 148158 551414 148394
rect 550794 148074 551414 148158
rect 550794 147838 550826 148074
rect 551062 147838 551146 148074
rect 551382 147838 551414 148074
rect 550794 146000 551414 147838
rect 559794 147454 560414 164898
rect 559794 147218 559826 147454
rect 560062 147218 560146 147454
rect 560382 147218 560414 147454
rect 559794 147134 560414 147218
rect 559794 146898 559826 147134
rect 560062 146898 560146 147134
rect 560382 146898 560414 147134
rect 10794 138218 10826 138454
rect 11062 138218 11146 138454
rect 11382 138218 11414 138454
rect 10794 138134 11414 138218
rect 10794 137898 10826 138134
rect 11062 137898 11146 138134
rect 11382 137898 11414 138134
rect 10794 120454 11414 137898
rect 22874 138454 23194 138486
rect 22874 138218 22916 138454
rect 23152 138218 23194 138454
rect 22874 138134 23194 138218
rect 22874 137898 22916 138134
rect 23152 137898 23194 138134
rect 22874 137866 23194 137898
rect 28805 138454 29125 138486
rect 28805 138218 28847 138454
rect 29083 138218 29125 138454
rect 28805 138134 29125 138218
rect 28805 137898 28847 138134
rect 29083 137898 29125 138134
rect 28805 137866 29125 137898
rect 49874 138454 50194 138486
rect 49874 138218 49916 138454
rect 50152 138218 50194 138454
rect 49874 138134 50194 138218
rect 49874 137898 49916 138134
rect 50152 137898 50194 138134
rect 49874 137866 50194 137898
rect 55805 138454 56125 138486
rect 55805 138218 55847 138454
rect 56083 138218 56125 138454
rect 55805 138134 56125 138218
rect 55805 137898 55847 138134
rect 56083 137898 56125 138134
rect 55805 137866 56125 137898
rect 76874 138454 77194 138486
rect 76874 138218 76916 138454
rect 77152 138218 77194 138454
rect 76874 138134 77194 138218
rect 76874 137898 76916 138134
rect 77152 137898 77194 138134
rect 76874 137866 77194 137898
rect 82805 138454 83125 138486
rect 82805 138218 82847 138454
rect 83083 138218 83125 138454
rect 82805 138134 83125 138218
rect 82805 137898 82847 138134
rect 83083 137898 83125 138134
rect 82805 137866 83125 137898
rect 103874 138454 104194 138486
rect 103874 138218 103916 138454
rect 104152 138218 104194 138454
rect 103874 138134 104194 138218
rect 103874 137898 103916 138134
rect 104152 137898 104194 138134
rect 103874 137866 104194 137898
rect 109805 138454 110125 138486
rect 109805 138218 109847 138454
rect 110083 138218 110125 138454
rect 109805 138134 110125 138218
rect 109805 137898 109847 138134
rect 110083 137898 110125 138134
rect 109805 137866 110125 137898
rect 130874 138454 131194 138486
rect 130874 138218 130916 138454
rect 131152 138218 131194 138454
rect 130874 138134 131194 138218
rect 130874 137898 130916 138134
rect 131152 137898 131194 138134
rect 130874 137866 131194 137898
rect 136805 138454 137125 138486
rect 136805 138218 136847 138454
rect 137083 138218 137125 138454
rect 136805 138134 137125 138218
rect 136805 137898 136847 138134
rect 137083 137898 137125 138134
rect 136805 137866 137125 137898
rect 157874 138454 158194 138486
rect 157874 138218 157916 138454
rect 158152 138218 158194 138454
rect 157874 138134 158194 138218
rect 157874 137898 157916 138134
rect 158152 137898 158194 138134
rect 157874 137866 158194 137898
rect 163805 138454 164125 138486
rect 163805 138218 163847 138454
rect 164083 138218 164125 138454
rect 163805 138134 164125 138218
rect 163805 137898 163847 138134
rect 164083 137898 164125 138134
rect 163805 137866 164125 137898
rect 184874 138454 185194 138486
rect 184874 138218 184916 138454
rect 185152 138218 185194 138454
rect 184874 138134 185194 138218
rect 184874 137898 184916 138134
rect 185152 137898 185194 138134
rect 184874 137866 185194 137898
rect 190805 138454 191125 138486
rect 190805 138218 190847 138454
rect 191083 138218 191125 138454
rect 190805 138134 191125 138218
rect 190805 137898 190847 138134
rect 191083 137898 191125 138134
rect 190805 137866 191125 137898
rect 211874 138454 212194 138486
rect 211874 138218 211916 138454
rect 212152 138218 212194 138454
rect 211874 138134 212194 138218
rect 211874 137898 211916 138134
rect 212152 137898 212194 138134
rect 211874 137866 212194 137898
rect 217805 138454 218125 138486
rect 217805 138218 217847 138454
rect 218083 138218 218125 138454
rect 217805 138134 218125 138218
rect 217805 137898 217847 138134
rect 218083 137898 218125 138134
rect 217805 137866 218125 137898
rect 238874 138454 239194 138486
rect 238874 138218 238916 138454
rect 239152 138218 239194 138454
rect 238874 138134 239194 138218
rect 238874 137898 238916 138134
rect 239152 137898 239194 138134
rect 238874 137866 239194 137898
rect 244805 138454 245125 138486
rect 244805 138218 244847 138454
rect 245083 138218 245125 138454
rect 244805 138134 245125 138218
rect 244805 137898 244847 138134
rect 245083 137898 245125 138134
rect 244805 137866 245125 137898
rect 265874 138454 266194 138486
rect 265874 138218 265916 138454
rect 266152 138218 266194 138454
rect 265874 138134 266194 138218
rect 265874 137898 265916 138134
rect 266152 137898 266194 138134
rect 265874 137866 266194 137898
rect 271805 138454 272125 138486
rect 271805 138218 271847 138454
rect 272083 138218 272125 138454
rect 271805 138134 272125 138218
rect 271805 137898 271847 138134
rect 272083 137898 272125 138134
rect 271805 137866 272125 137898
rect 292874 138454 293194 138486
rect 292874 138218 292916 138454
rect 293152 138218 293194 138454
rect 292874 138134 293194 138218
rect 292874 137898 292916 138134
rect 293152 137898 293194 138134
rect 292874 137866 293194 137898
rect 298805 138454 299125 138486
rect 298805 138218 298847 138454
rect 299083 138218 299125 138454
rect 298805 138134 299125 138218
rect 298805 137898 298847 138134
rect 299083 137898 299125 138134
rect 298805 137866 299125 137898
rect 319874 138454 320194 138486
rect 319874 138218 319916 138454
rect 320152 138218 320194 138454
rect 319874 138134 320194 138218
rect 319874 137898 319916 138134
rect 320152 137898 320194 138134
rect 319874 137866 320194 137898
rect 325805 138454 326125 138486
rect 325805 138218 325847 138454
rect 326083 138218 326125 138454
rect 325805 138134 326125 138218
rect 325805 137898 325847 138134
rect 326083 137898 326125 138134
rect 325805 137866 326125 137898
rect 346874 138454 347194 138486
rect 346874 138218 346916 138454
rect 347152 138218 347194 138454
rect 346874 138134 347194 138218
rect 346874 137898 346916 138134
rect 347152 137898 347194 138134
rect 346874 137866 347194 137898
rect 352805 138454 353125 138486
rect 352805 138218 352847 138454
rect 353083 138218 353125 138454
rect 352805 138134 353125 138218
rect 352805 137898 352847 138134
rect 353083 137898 353125 138134
rect 352805 137866 353125 137898
rect 373874 138454 374194 138486
rect 373874 138218 373916 138454
rect 374152 138218 374194 138454
rect 373874 138134 374194 138218
rect 373874 137898 373916 138134
rect 374152 137898 374194 138134
rect 373874 137866 374194 137898
rect 379805 138454 380125 138486
rect 379805 138218 379847 138454
rect 380083 138218 380125 138454
rect 379805 138134 380125 138218
rect 379805 137898 379847 138134
rect 380083 137898 380125 138134
rect 379805 137866 380125 137898
rect 400874 138454 401194 138486
rect 400874 138218 400916 138454
rect 401152 138218 401194 138454
rect 400874 138134 401194 138218
rect 400874 137898 400916 138134
rect 401152 137898 401194 138134
rect 400874 137866 401194 137898
rect 406805 138454 407125 138486
rect 406805 138218 406847 138454
rect 407083 138218 407125 138454
rect 406805 138134 407125 138218
rect 406805 137898 406847 138134
rect 407083 137898 407125 138134
rect 406805 137866 407125 137898
rect 427874 138454 428194 138486
rect 427874 138218 427916 138454
rect 428152 138218 428194 138454
rect 427874 138134 428194 138218
rect 427874 137898 427916 138134
rect 428152 137898 428194 138134
rect 427874 137866 428194 137898
rect 433805 138454 434125 138486
rect 433805 138218 433847 138454
rect 434083 138218 434125 138454
rect 433805 138134 434125 138218
rect 433805 137898 433847 138134
rect 434083 137898 434125 138134
rect 433805 137866 434125 137898
rect 454874 138454 455194 138486
rect 454874 138218 454916 138454
rect 455152 138218 455194 138454
rect 454874 138134 455194 138218
rect 454874 137898 454916 138134
rect 455152 137898 455194 138134
rect 454874 137866 455194 137898
rect 460805 138454 461125 138486
rect 460805 138218 460847 138454
rect 461083 138218 461125 138454
rect 460805 138134 461125 138218
rect 460805 137898 460847 138134
rect 461083 137898 461125 138134
rect 460805 137866 461125 137898
rect 481874 138454 482194 138486
rect 481874 138218 481916 138454
rect 482152 138218 482194 138454
rect 481874 138134 482194 138218
rect 481874 137898 481916 138134
rect 482152 137898 482194 138134
rect 481874 137866 482194 137898
rect 487805 138454 488125 138486
rect 487805 138218 487847 138454
rect 488083 138218 488125 138454
rect 487805 138134 488125 138218
rect 487805 137898 487847 138134
rect 488083 137898 488125 138134
rect 487805 137866 488125 137898
rect 508874 138454 509194 138486
rect 508874 138218 508916 138454
rect 509152 138218 509194 138454
rect 508874 138134 509194 138218
rect 508874 137898 508916 138134
rect 509152 137898 509194 138134
rect 508874 137866 509194 137898
rect 514805 138454 515125 138486
rect 514805 138218 514847 138454
rect 515083 138218 515125 138454
rect 514805 138134 515125 138218
rect 514805 137898 514847 138134
rect 515083 137898 515125 138134
rect 514805 137866 515125 137898
rect 535874 138454 536194 138486
rect 535874 138218 535916 138454
rect 536152 138218 536194 138454
rect 535874 138134 536194 138218
rect 535874 137898 535916 138134
rect 536152 137898 536194 138134
rect 535874 137866 536194 137898
rect 541805 138454 542125 138486
rect 541805 138218 541847 138454
rect 542083 138218 542125 138454
rect 541805 138134 542125 138218
rect 541805 137898 541847 138134
rect 542083 137898 542125 138134
rect 541805 137866 542125 137898
rect 19910 129454 20230 129486
rect 19910 129218 19952 129454
rect 20188 129218 20230 129454
rect 19910 129134 20230 129218
rect 19910 128898 19952 129134
rect 20188 128898 20230 129134
rect 19910 128866 20230 128898
rect 25840 129454 26160 129486
rect 25840 129218 25882 129454
rect 26118 129218 26160 129454
rect 25840 129134 26160 129218
rect 25840 128898 25882 129134
rect 26118 128898 26160 129134
rect 25840 128866 26160 128898
rect 31771 129454 32091 129486
rect 31771 129218 31813 129454
rect 32049 129218 32091 129454
rect 31771 129134 32091 129218
rect 31771 128898 31813 129134
rect 32049 128898 32091 129134
rect 31771 128866 32091 128898
rect 46910 129454 47230 129486
rect 46910 129218 46952 129454
rect 47188 129218 47230 129454
rect 46910 129134 47230 129218
rect 46910 128898 46952 129134
rect 47188 128898 47230 129134
rect 46910 128866 47230 128898
rect 52840 129454 53160 129486
rect 52840 129218 52882 129454
rect 53118 129218 53160 129454
rect 52840 129134 53160 129218
rect 52840 128898 52882 129134
rect 53118 128898 53160 129134
rect 52840 128866 53160 128898
rect 58771 129454 59091 129486
rect 58771 129218 58813 129454
rect 59049 129218 59091 129454
rect 58771 129134 59091 129218
rect 58771 128898 58813 129134
rect 59049 128898 59091 129134
rect 58771 128866 59091 128898
rect 73910 129454 74230 129486
rect 73910 129218 73952 129454
rect 74188 129218 74230 129454
rect 73910 129134 74230 129218
rect 73910 128898 73952 129134
rect 74188 128898 74230 129134
rect 73910 128866 74230 128898
rect 79840 129454 80160 129486
rect 79840 129218 79882 129454
rect 80118 129218 80160 129454
rect 79840 129134 80160 129218
rect 79840 128898 79882 129134
rect 80118 128898 80160 129134
rect 79840 128866 80160 128898
rect 85771 129454 86091 129486
rect 85771 129218 85813 129454
rect 86049 129218 86091 129454
rect 85771 129134 86091 129218
rect 85771 128898 85813 129134
rect 86049 128898 86091 129134
rect 85771 128866 86091 128898
rect 100910 129454 101230 129486
rect 100910 129218 100952 129454
rect 101188 129218 101230 129454
rect 100910 129134 101230 129218
rect 100910 128898 100952 129134
rect 101188 128898 101230 129134
rect 100910 128866 101230 128898
rect 106840 129454 107160 129486
rect 106840 129218 106882 129454
rect 107118 129218 107160 129454
rect 106840 129134 107160 129218
rect 106840 128898 106882 129134
rect 107118 128898 107160 129134
rect 106840 128866 107160 128898
rect 112771 129454 113091 129486
rect 112771 129218 112813 129454
rect 113049 129218 113091 129454
rect 112771 129134 113091 129218
rect 112771 128898 112813 129134
rect 113049 128898 113091 129134
rect 112771 128866 113091 128898
rect 127910 129454 128230 129486
rect 127910 129218 127952 129454
rect 128188 129218 128230 129454
rect 127910 129134 128230 129218
rect 127910 128898 127952 129134
rect 128188 128898 128230 129134
rect 127910 128866 128230 128898
rect 133840 129454 134160 129486
rect 133840 129218 133882 129454
rect 134118 129218 134160 129454
rect 133840 129134 134160 129218
rect 133840 128898 133882 129134
rect 134118 128898 134160 129134
rect 133840 128866 134160 128898
rect 139771 129454 140091 129486
rect 139771 129218 139813 129454
rect 140049 129218 140091 129454
rect 139771 129134 140091 129218
rect 139771 128898 139813 129134
rect 140049 128898 140091 129134
rect 139771 128866 140091 128898
rect 154910 129454 155230 129486
rect 154910 129218 154952 129454
rect 155188 129218 155230 129454
rect 154910 129134 155230 129218
rect 154910 128898 154952 129134
rect 155188 128898 155230 129134
rect 154910 128866 155230 128898
rect 160840 129454 161160 129486
rect 160840 129218 160882 129454
rect 161118 129218 161160 129454
rect 160840 129134 161160 129218
rect 160840 128898 160882 129134
rect 161118 128898 161160 129134
rect 160840 128866 161160 128898
rect 166771 129454 167091 129486
rect 166771 129218 166813 129454
rect 167049 129218 167091 129454
rect 166771 129134 167091 129218
rect 166771 128898 166813 129134
rect 167049 128898 167091 129134
rect 166771 128866 167091 128898
rect 181910 129454 182230 129486
rect 181910 129218 181952 129454
rect 182188 129218 182230 129454
rect 181910 129134 182230 129218
rect 181910 128898 181952 129134
rect 182188 128898 182230 129134
rect 181910 128866 182230 128898
rect 187840 129454 188160 129486
rect 187840 129218 187882 129454
rect 188118 129218 188160 129454
rect 187840 129134 188160 129218
rect 187840 128898 187882 129134
rect 188118 128898 188160 129134
rect 187840 128866 188160 128898
rect 193771 129454 194091 129486
rect 193771 129218 193813 129454
rect 194049 129218 194091 129454
rect 193771 129134 194091 129218
rect 193771 128898 193813 129134
rect 194049 128898 194091 129134
rect 193771 128866 194091 128898
rect 208910 129454 209230 129486
rect 208910 129218 208952 129454
rect 209188 129218 209230 129454
rect 208910 129134 209230 129218
rect 208910 128898 208952 129134
rect 209188 128898 209230 129134
rect 208910 128866 209230 128898
rect 214840 129454 215160 129486
rect 214840 129218 214882 129454
rect 215118 129218 215160 129454
rect 214840 129134 215160 129218
rect 214840 128898 214882 129134
rect 215118 128898 215160 129134
rect 214840 128866 215160 128898
rect 220771 129454 221091 129486
rect 220771 129218 220813 129454
rect 221049 129218 221091 129454
rect 220771 129134 221091 129218
rect 220771 128898 220813 129134
rect 221049 128898 221091 129134
rect 220771 128866 221091 128898
rect 235910 129454 236230 129486
rect 235910 129218 235952 129454
rect 236188 129218 236230 129454
rect 235910 129134 236230 129218
rect 235910 128898 235952 129134
rect 236188 128898 236230 129134
rect 235910 128866 236230 128898
rect 241840 129454 242160 129486
rect 241840 129218 241882 129454
rect 242118 129218 242160 129454
rect 241840 129134 242160 129218
rect 241840 128898 241882 129134
rect 242118 128898 242160 129134
rect 241840 128866 242160 128898
rect 247771 129454 248091 129486
rect 247771 129218 247813 129454
rect 248049 129218 248091 129454
rect 247771 129134 248091 129218
rect 247771 128898 247813 129134
rect 248049 128898 248091 129134
rect 247771 128866 248091 128898
rect 262910 129454 263230 129486
rect 262910 129218 262952 129454
rect 263188 129218 263230 129454
rect 262910 129134 263230 129218
rect 262910 128898 262952 129134
rect 263188 128898 263230 129134
rect 262910 128866 263230 128898
rect 268840 129454 269160 129486
rect 268840 129218 268882 129454
rect 269118 129218 269160 129454
rect 268840 129134 269160 129218
rect 268840 128898 268882 129134
rect 269118 128898 269160 129134
rect 268840 128866 269160 128898
rect 274771 129454 275091 129486
rect 274771 129218 274813 129454
rect 275049 129218 275091 129454
rect 274771 129134 275091 129218
rect 274771 128898 274813 129134
rect 275049 128898 275091 129134
rect 274771 128866 275091 128898
rect 289910 129454 290230 129486
rect 289910 129218 289952 129454
rect 290188 129218 290230 129454
rect 289910 129134 290230 129218
rect 289910 128898 289952 129134
rect 290188 128898 290230 129134
rect 289910 128866 290230 128898
rect 295840 129454 296160 129486
rect 295840 129218 295882 129454
rect 296118 129218 296160 129454
rect 295840 129134 296160 129218
rect 295840 128898 295882 129134
rect 296118 128898 296160 129134
rect 295840 128866 296160 128898
rect 301771 129454 302091 129486
rect 301771 129218 301813 129454
rect 302049 129218 302091 129454
rect 301771 129134 302091 129218
rect 301771 128898 301813 129134
rect 302049 128898 302091 129134
rect 301771 128866 302091 128898
rect 316910 129454 317230 129486
rect 316910 129218 316952 129454
rect 317188 129218 317230 129454
rect 316910 129134 317230 129218
rect 316910 128898 316952 129134
rect 317188 128898 317230 129134
rect 316910 128866 317230 128898
rect 322840 129454 323160 129486
rect 322840 129218 322882 129454
rect 323118 129218 323160 129454
rect 322840 129134 323160 129218
rect 322840 128898 322882 129134
rect 323118 128898 323160 129134
rect 322840 128866 323160 128898
rect 328771 129454 329091 129486
rect 328771 129218 328813 129454
rect 329049 129218 329091 129454
rect 328771 129134 329091 129218
rect 328771 128898 328813 129134
rect 329049 128898 329091 129134
rect 328771 128866 329091 128898
rect 343910 129454 344230 129486
rect 343910 129218 343952 129454
rect 344188 129218 344230 129454
rect 343910 129134 344230 129218
rect 343910 128898 343952 129134
rect 344188 128898 344230 129134
rect 343910 128866 344230 128898
rect 349840 129454 350160 129486
rect 349840 129218 349882 129454
rect 350118 129218 350160 129454
rect 349840 129134 350160 129218
rect 349840 128898 349882 129134
rect 350118 128898 350160 129134
rect 349840 128866 350160 128898
rect 355771 129454 356091 129486
rect 355771 129218 355813 129454
rect 356049 129218 356091 129454
rect 355771 129134 356091 129218
rect 355771 128898 355813 129134
rect 356049 128898 356091 129134
rect 355771 128866 356091 128898
rect 370910 129454 371230 129486
rect 370910 129218 370952 129454
rect 371188 129218 371230 129454
rect 370910 129134 371230 129218
rect 370910 128898 370952 129134
rect 371188 128898 371230 129134
rect 370910 128866 371230 128898
rect 376840 129454 377160 129486
rect 376840 129218 376882 129454
rect 377118 129218 377160 129454
rect 376840 129134 377160 129218
rect 376840 128898 376882 129134
rect 377118 128898 377160 129134
rect 376840 128866 377160 128898
rect 382771 129454 383091 129486
rect 382771 129218 382813 129454
rect 383049 129218 383091 129454
rect 382771 129134 383091 129218
rect 382771 128898 382813 129134
rect 383049 128898 383091 129134
rect 382771 128866 383091 128898
rect 397910 129454 398230 129486
rect 397910 129218 397952 129454
rect 398188 129218 398230 129454
rect 397910 129134 398230 129218
rect 397910 128898 397952 129134
rect 398188 128898 398230 129134
rect 397910 128866 398230 128898
rect 403840 129454 404160 129486
rect 403840 129218 403882 129454
rect 404118 129218 404160 129454
rect 403840 129134 404160 129218
rect 403840 128898 403882 129134
rect 404118 128898 404160 129134
rect 403840 128866 404160 128898
rect 409771 129454 410091 129486
rect 409771 129218 409813 129454
rect 410049 129218 410091 129454
rect 409771 129134 410091 129218
rect 409771 128898 409813 129134
rect 410049 128898 410091 129134
rect 409771 128866 410091 128898
rect 424910 129454 425230 129486
rect 424910 129218 424952 129454
rect 425188 129218 425230 129454
rect 424910 129134 425230 129218
rect 424910 128898 424952 129134
rect 425188 128898 425230 129134
rect 424910 128866 425230 128898
rect 430840 129454 431160 129486
rect 430840 129218 430882 129454
rect 431118 129218 431160 129454
rect 430840 129134 431160 129218
rect 430840 128898 430882 129134
rect 431118 128898 431160 129134
rect 430840 128866 431160 128898
rect 436771 129454 437091 129486
rect 436771 129218 436813 129454
rect 437049 129218 437091 129454
rect 436771 129134 437091 129218
rect 436771 128898 436813 129134
rect 437049 128898 437091 129134
rect 436771 128866 437091 128898
rect 451910 129454 452230 129486
rect 451910 129218 451952 129454
rect 452188 129218 452230 129454
rect 451910 129134 452230 129218
rect 451910 128898 451952 129134
rect 452188 128898 452230 129134
rect 451910 128866 452230 128898
rect 457840 129454 458160 129486
rect 457840 129218 457882 129454
rect 458118 129218 458160 129454
rect 457840 129134 458160 129218
rect 457840 128898 457882 129134
rect 458118 128898 458160 129134
rect 457840 128866 458160 128898
rect 463771 129454 464091 129486
rect 463771 129218 463813 129454
rect 464049 129218 464091 129454
rect 463771 129134 464091 129218
rect 463771 128898 463813 129134
rect 464049 128898 464091 129134
rect 463771 128866 464091 128898
rect 478910 129454 479230 129486
rect 478910 129218 478952 129454
rect 479188 129218 479230 129454
rect 478910 129134 479230 129218
rect 478910 128898 478952 129134
rect 479188 128898 479230 129134
rect 478910 128866 479230 128898
rect 484840 129454 485160 129486
rect 484840 129218 484882 129454
rect 485118 129218 485160 129454
rect 484840 129134 485160 129218
rect 484840 128898 484882 129134
rect 485118 128898 485160 129134
rect 484840 128866 485160 128898
rect 490771 129454 491091 129486
rect 490771 129218 490813 129454
rect 491049 129218 491091 129454
rect 490771 129134 491091 129218
rect 490771 128898 490813 129134
rect 491049 128898 491091 129134
rect 490771 128866 491091 128898
rect 505910 129454 506230 129486
rect 505910 129218 505952 129454
rect 506188 129218 506230 129454
rect 505910 129134 506230 129218
rect 505910 128898 505952 129134
rect 506188 128898 506230 129134
rect 505910 128866 506230 128898
rect 511840 129454 512160 129486
rect 511840 129218 511882 129454
rect 512118 129218 512160 129454
rect 511840 129134 512160 129218
rect 511840 128898 511882 129134
rect 512118 128898 512160 129134
rect 511840 128866 512160 128898
rect 517771 129454 518091 129486
rect 517771 129218 517813 129454
rect 518049 129218 518091 129454
rect 517771 129134 518091 129218
rect 517771 128898 517813 129134
rect 518049 128898 518091 129134
rect 517771 128866 518091 128898
rect 532910 129454 533230 129486
rect 532910 129218 532952 129454
rect 533188 129218 533230 129454
rect 532910 129134 533230 129218
rect 532910 128898 532952 129134
rect 533188 128898 533230 129134
rect 532910 128866 533230 128898
rect 538840 129454 539160 129486
rect 538840 129218 538882 129454
rect 539118 129218 539160 129454
rect 538840 129134 539160 129218
rect 538840 128898 538882 129134
rect 539118 128898 539160 129134
rect 538840 128866 539160 128898
rect 544771 129454 545091 129486
rect 544771 129218 544813 129454
rect 545049 129218 545091 129454
rect 544771 129134 545091 129218
rect 544771 128898 544813 129134
rect 545049 128898 545091 129134
rect 544771 128866 545091 128898
rect 559794 129454 560414 146898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 102454 11414 119898
rect 19794 121394 20414 122000
rect 19794 121158 19826 121394
rect 20062 121158 20146 121394
rect 20382 121158 20414 121394
rect 19794 121074 20414 121158
rect 19794 120838 19826 121074
rect 20062 120838 20146 121074
rect 20382 120838 20414 121074
rect 19794 119000 20414 120838
rect 28794 120454 29414 122000
rect 28794 120218 28826 120454
rect 29062 120218 29146 120454
rect 29382 120218 29414 120454
rect 28794 120134 29414 120218
rect 28794 119898 28826 120134
rect 29062 119898 29146 120134
rect 29382 119898 29414 120134
rect 28794 119000 29414 119898
rect 37794 121394 38414 122000
rect 37794 121158 37826 121394
rect 38062 121158 38146 121394
rect 38382 121158 38414 121394
rect 37794 121074 38414 121158
rect 37794 120838 37826 121074
rect 38062 120838 38146 121074
rect 38382 120838 38414 121074
rect 37794 119000 38414 120838
rect 46794 120454 47414 122000
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 119000 47414 119898
rect 55794 121394 56414 122000
rect 55794 121158 55826 121394
rect 56062 121158 56146 121394
rect 56382 121158 56414 121394
rect 55794 121074 56414 121158
rect 55794 120838 55826 121074
rect 56062 120838 56146 121074
rect 56382 120838 56414 121074
rect 55794 119000 56414 120838
rect 64794 120454 65414 122000
rect 64794 120218 64826 120454
rect 65062 120218 65146 120454
rect 65382 120218 65414 120454
rect 64794 120134 65414 120218
rect 64794 119898 64826 120134
rect 65062 119898 65146 120134
rect 65382 119898 65414 120134
rect 64794 119000 65414 119898
rect 73794 121394 74414 122000
rect 73794 121158 73826 121394
rect 74062 121158 74146 121394
rect 74382 121158 74414 121394
rect 73794 121074 74414 121158
rect 73794 120838 73826 121074
rect 74062 120838 74146 121074
rect 74382 120838 74414 121074
rect 73794 119000 74414 120838
rect 82794 120454 83414 122000
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 119000 83414 119898
rect 91794 121394 92414 122000
rect 91794 121158 91826 121394
rect 92062 121158 92146 121394
rect 92382 121158 92414 121394
rect 91794 121074 92414 121158
rect 91794 120838 91826 121074
rect 92062 120838 92146 121074
rect 92382 120838 92414 121074
rect 91794 119000 92414 120838
rect 100794 120454 101414 122000
rect 100794 120218 100826 120454
rect 101062 120218 101146 120454
rect 101382 120218 101414 120454
rect 100794 120134 101414 120218
rect 100794 119898 100826 120134
rect 101062 119898 101146 120134
rect 101382 119898 101414 120134
rect 100794 119000 101414 119898
rect 109794 121394 110414 122000
rect 109794 121158 109826 121394
rect 110062 121158 110146 121394
rect 110382 121158 110414 121394
rect 109794 121074 110414 121158
rect 109794 120838 109826 121074
rect 110062 120838 110146 121074
rect 110382 120838 110414 121074
rect 109794 119000 110414 120838
rect 118794 120454 119414 122000
rect 118794 120218 118826 120454
rect 119062 120218 119146 120454
rect 119382 120218 119414 120454
rect 118794 120134 119414 120218
rect 118794 119898 118826 120134
rect 119062 119898 119146 120134
rect 119382 119898 119414 120134
rect 118794 119000 119414 119898
rect 127794 121394 128414 122000
rect 127794 121158 127826 121394
rect 128062 121158 128146 121394
rect 128382 121158 128414 121394
rect 127794 121074 128414 121158
rect 127794 120838 127826 121074
rect 128062 120838 128146 121074
rect 128382 120838 128414 121074
rect 127794 119000 128414 120838
rect 136794 120454 137414 122000
rect 136794 120218 136826 120454
rect 137062 120218 137146 120454
rect 137382 120218 137414 120454
rect 136794 120134 137414 120218
rect 136794 119898 136826 120134
rect 137062 119898 137146 120134
rect 137382 119898 137414 120134
rect 136794 119000 137414 119898
rect 145794 121394 146414 122000
rect 145794 121158 145826 121394
rect 146062 121158 146146 121394
rect 146382 121158 146414 121394
rect 145794 121074 146414 121158
rect 145794 120838 145826 121074
rect 146062 120838 146146 121074
rect 146382 120838 146414 121074
rect 145794 119000 146414 120838
rect 154794 120454 155414 122000
rect 154794 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 155414 120454
rect 154794 120134 155414 120218
rect 154794 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 155414 120134
rect 154794 119000 155414 119898
rect 163794 121394 164414 122000
rect 163794 121158 163826 121394
rect 164062 121158 164146 121394
rect 164382 121158 164414 121394
rect 163794 121074 164414 121158
rect 163794 120838 163826 121074
rect 164062 120838 164146 121074
rect 164382 120838 164414 121074
rect 163794 119000 164414 120838
rect 172794 120454 173414 122000
rect 172794 120218 172826 120454
rect 173062 120218 173146 120454
rect 173382 120218 173414 120454
rect 172794 120134 173414 120218
rect 172794 119898 172826 120134
rect 173062 119898 173146 120134
rect 173382 119898 173414 120134
rect 172794 119000 173414 119898
rect 181794 121394 182414 122000
rect 181794 121158 181826 121394
rect 182062 121158 182146 121394
rect 182382 121158 182414 121394
rect 181794 121074 182414 121158
rect 181794 120838 181826 121074
rect 182062 120838 182146 121074
rect 182382 120838 182414 121074
rect 181794 119000 182414 120838
rect 190794 120454 191414 122000
rect 190794 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 191414 120454
rect 190794 120134 191414 120218
rect 190794 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 191414 120134
rect 190794 119000 191414 119898
rect 199794 121394 200414 122000
rect 199794 121158 199826 121394
rect 200062 121158 200146 121394
rect 200382 121158 200414 121394
rect 199794 121074 200414 121158
rect 199794 120838 199826 121074
rect 200062 120838 200146 121074
rect 200382 120838 200414 121074
rect 199794 119000 200414 120838
rect 208794 120454 209414 122000
rect 208794 120218 208826 120454
rect 209062 120218 209146 120454
rect 209382 120218 209414 120454
rect 208794 120134 209414 120218
rect 208794 119898 208826 120134
rect 209062 119898 209146 120134
rect 209382 119898 209414 120134
rect 208794 119000 209414 119898
rect 217794 121394 218414 122000
rect 217794 121158 217826 121394
rect 218062 121158 218146 121394
rect 218382 121158 218414 121394
rect 217794 121074 218414 121158
rect 217794 120838 217826 121074
rect 218062 120838 218146 121074
rect 218382 120838 218414 121074
rect 217794 119000 218414 120838
rect 226794 120454 227414 122000
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 119000 227414 119898
rect 235794 121394 236414 122000
rect 235794 121158 235826 121394
rect 236062 121158 236146 121394
rect 236382 121158 236414 121394
rect 235794 121074 236414 121158
rect 235794 120838 235826 121074
rect 236062 120838 236146 121074
rect 236382 120838 236414 121074
rect 235794 119000 236414 120838
rect 244794 120454 245414 122000
rect 244794 120218 244826 120454
rect 245062 120218 245146 120454
rect 245382 120218 245414 120454
rect 244794 120134 245414 120218
rect 244794 119898 244826 120134
rect 245062 119898 245146 120134
rect 245382 119898 245414 120134
rect 244794 119000 245414 119898
rect 253794 121394 254414 122000
rect 253794 121158 253826 121394
rect 254062 121158 254146 121394
rect 254382 121158 254414 121394
rect 253794 121074 254414 121158
rect 253794 120838 253826 121074
rect 254062 120838 254146 121074
rect 254382 120838 254414 121074
rect 253794 119000 254414 120838
rect 262794 120454 263414 122000
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 119000 263414 119898
rect 271794 121394 272414 122000
rect 271794 121158 271826 121394
rect 272062 121158 272146 121394
rect 272382 121158 272414 121394
rect 271794 121074 272414 121158
rect 271794 120838 271826 121074
rect 272062 120838 272146 121074
rect 272382 120838 272414 121074
rect 271794 119000 272414 120838
rect 280794 120454 281414 122000
rect 280794 120218 280826 120454
rect 281062 120218 281146 120454
rect 281382 120218 281414 120454
rect 280794 120134 281414 120218
rect 280794 119898 280826 120134
rect 281062 119898 281146 120134
rect 281382 119898 281414 120134
rect 280794 119000 281414 119898
rect 289794 121394 290414 122000
rect 289794 121158 289826 121394
rect 290062 121158 290146 121394
rect 290382 121158 290414 121394
rect 289794 121074 290414 121158
rect 289794 120838 289826 121074
rect 290062 120838 290146 121074
rect 290382 120838 290414 121074
rect 289794 119000 290414 120838
rect 298794 120454 299414 122000
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 119000 299414 119898
rect 307794 121394 308414 122000
rect 307794 121158 307826 121394
rect 308062 121158 308146 121394
rect 308382 121158 308414 121394
rect 307794 121074 308414 121158
rect 307794 120838 307826 121074
rect 308062 120838 308146 121074
rect 308382 120838 308414 121074
rect 307794 119000 308414 120838
rect 316794 120454 317414 122000
rect 316794 120218 316826 120454
rect 317062 120218 317146 120454
rect 317382 120218 317414 120454
rect 316794 120134 317414 120218
rect 316794 119898 316826 120134
rect 317062 119898 317146 120134
rect 317382 119898 317414 120134
rect 316794 119000 317414 119898
rect 325794 121394 326414 122000
rect 325794 121158 325826 121394
rect 326062 121158 326146 121394
rect 326382 121158 326414 121394
rect 325794 121074 326414 121158
rect 325794 120838 325826 121074
rect 326062 120838 326146 121074
rect 326382 120838 326414 121074
rect 325794 119000 326414 120838
rect 334794 120454 335414 122000
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 119000 335414 119898
rect 343794 121394 344414 122000
rect 343794 121158 343826 121394
rect 344062 121158 344146 121394
rect 344382 121158 344414 121394
rect 343794 121074 344414 121158
rect 343794 120838 343826 121074
rect 344062 120838 344146 121074
rect 344382 120838 344414 121074
rect 343794 119000 344414 120838
rect 352794 120454 353414 122000
rect 352794 120218 352826 120454
rect 353062 120218 353146 120454
rect 353382 120218 353414 120454
rect 352794 120134 353414 120218
rect 352794 119898 352826 120134
rect 353062 119898 353146 120134
rect 353382 119898 353414 120134
rect 352794 119000 353414 119898
rect 361794 121394 362414 122000
rect 361794 121158 361826 121394
rect 362062 121158 362146 121394
rect 362382 121158 362414 121394
rect 361794 121074 362414 121158
rect 361794 120838 361826 121074
rect 362062 120838 362146 121074
rect 362382 120838 362414 121074
rect 361794 119000 362414 120838
rect 370794 120454 371414 122000
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 119000 371414 119898
rect 379794 121394 380414 122000
rect 379794 121158 379826 121394
rect 380062 121158 380146 121394
rect 380382 121158 380414 121394
rect 379794 121074 380414 121158
rect 379794 120838 379826 121074
rect 380062 120838 380146 121074
rect 380382 120838 380414 121074
rect 379794 119000 380414 120838
rect 388794 120454 389414 122000
rect 388794 120218 388826 120454
rect 389062 120218 389146 120454
rect 389382 120218 389414 120454
rect 388794 120134 389414 120218
rect 388794 119898 388826 120134
rect 389062 119898 389146 120134
rect 389382 119898 389414 120134
rect 388794 119000 389414 119898
rect 397794 121394 398414 122000
rect 397794 121158 397826 121394
rect 398062 121158 398146 121394
rect 398382 121158 398414 121394
rect 397794 121074 398414 121158
rect 397794 120838 397826 121074
rect 398062 120838 398146 121074
rect 398382 120838 398414 121074
rect 397794 119000 398414 120838
rect 406794 120454 407414 122000
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 119000 407414 119898
rect 415794 121394 416414 122000
rect 415794 121158 415826 121394
rect 416062 121158 416146 121394
rect 416382 121158 416414 121394
rect 415794 121074 416414 121158
rect 415794 120838 415826 121074
rect 416062 120838 416146 121074
rect 416382 120838 416414 121074
rect 415794 119000 416414 120838
rect 424794 120454 425414 122000
rect 424794 120218 424826 120454
rect 425062 120218 425146 120454
rect 425382 120218 425414 120454
rect 424794 120134 425414 120218
rect 424794 119898 424826 120134
rect 425062 119898 425146 120134
rect 425382 119898 425414 120134
rect 424794 119000 425414 119898
rect 433794 121394 434414 122000
rect 433794 121158 433826 121394
rect 434062 121158 434146 121394
rect 434382 121158 434414 121394
rect 433794 121074 434414 121158
rect 433794 120838 433826 121074
rect 434062 120838 434146 121074
rect 434382 120838 434414 121074
rect 433794 119000 434414 120838
rect 442794 120454 443414 122000
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 119000 443414 119898
rect 451794 121394 452414 122000
rect 451794 121158 451826 121394
rect 452062 121158 452146 121394
rect 452382 121158 452414 121394
rect 451794 121074 452414 121158
rect 451794 120838 451826 121074
rect 452062 120838 452146 121074
rect 452382 120838 452414 121074
rect 451794 119000 452414 120838
rect 460794 120454 461414 122000
rect 460794 120218 460826 120454
rect 461062 120218 461146 120454
rect 461382 120218 461414 120454
rect 460794 120134 461414 120218
rect 460794 119898 460826 120134
rect 461062 119898 461146 120134
rect 461382 119898 461414 120134
rect 460794 119000 461414 119898
rect 469794 121394 470414 122000
rect 469794 121158 469826 121394
rect 470062 121158 470146 121394
rect 470382 121158 470414 121394
rect 469794 121074 470414 121158
rect 469794 120838 469826 121074
rect 470062 120838 470146 121074
rect 470382 120838 470414 121074
rect 469794 119000 470414 120838
rect 478794 120454 479414 122000
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 119000 479414 119898
rect 487794 121394 488414 122000
rect 487794 121158 487826 121394
rect 488062 121158 488146 121394
rect 488382 121158 488414 121394
rect 487794 121074 488414 121158
rect 487794 120838 487826 121074
rect 488062 120838 488146 121074
rect 488382 120838 488414 121074
rect 487794 119000 488414 120838
rect 496794 120454 497414 122000
rect 496794 120218 496826 120454
rect 497062 120218 497146 120454
rect 497382 120218 497414 120454
rect 496794 120134 497414 120218
rect 496794 119898 496826 120134
rect 497062 119898 497146 120134
rect 497382 119898 497414 120134
rect 496794 119000 497414 119898
rect 505794 121394 506414 122000
rect 505794 121158 505826 121394
rect 506062 121158 506146 121394
rect 506382 121158 506414 121394
rect 505794 121074 506414 121158
rect 505794 120838 505826 121074
rect 506062 120838 506146 121074
rect 506382 120838 506414 121074
rect 505794 119000 506414 120838
rect 514794 120454 515414 122000
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 119000 515414 119898
rect 523794 121394 524414 122000
rect 523794 121158 523826 121394
rect 524062 121158 524146 121394
rect 524382 121158 524414 121394
rect 523794 121074 524414 121158
rect 523794 120838 523826 121074
rect 524062 120838 524146 121074
rect 524382 120838 524414 121074
rect 523794 119000 524414 120838
rect 532794 120454 533414 122000
rect 532794 120218 532826 120454
rect 533062 120218 533146 120454
rect 533382 120218 533414 120454
rect 532794 120134 533414 120218
rect 532794 119898 532826 120134
rect 533062 119898 533146 120134
rect 533382 119898 533414 120134
rect 532794 119000 533414 119898
rect 541794 121394 542414 122000
rect 541794 121158 541826 121394
rect 542062 121158 542146 121394
rect 542382 121158 542414 121394
rect 541794 121074 542414 121158
rect 541794 120838 541826 121074
rect 542062 120838 542146 121074
rect 542382 120838 542414 121074
rect 541794 119000 542414 120838
rect 550794 120454 551414 122000
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 119000 551414 119898
rect 19910 111454 20230 111486
rect 19910 111218 19952 111454
rect 20188 111218 20230 111454
rect 19910 111134 20230 111218
rect 19910 110898 19952 111134
rect 20188 110898 20230 111134
rect 19910 110866 20230 110898
rect 25840 111454 26160 111486
rect 25840 111218 25882 111454
rect 26118 111218 26160 111454
rect 25840 111134 26160 111218
rect 25840 110898 25882 111134
rect 26118 110898 26160 111134
rect 25840 110866 26160 110898
rect 31771 111454 32091 111486
rect 31771 111218 31813 111454
rect 32049 111218 32091 111454
rect 31771 111134 32091 111218
rect 31771 110898 31813 111134
rect 32049 110898 32091 111134
rect 31771 110866 32091 110898
rect 46910 111454 47230 111486
rect 46910 111218 46952 111454
rect 47188 111218 47230 111454
rect 46910 111134 47230 111218
rect 46910 110898 46952 111134
rect 47188 110898 47230 111134
rect 46910 110866 47230 110898
rect 52840 111454 53160 111486
rect 52840 111218 52882 111454
rect 53118 111218 53160 111454
rect 52840 111134 53160 111218
rect 52840 110898 52882 111134
rect 53118 110898 53160 111134
rect 52840 110866 53160 110898
rect 58771 111454 59091 111486
rect 58771 111218 58813 111454
rect 59049 111218 59091 111454
rect 58771 111134 59091 111218
rect 58771 110898 58813 111134
rect 59049 110898 59091 111134
rect 58771 110866 59091 110898
rect 73910 111454 74230 111486
rect 73910 111218 73952 111454
rect 74188 111218 74230 111454
rect 73910 111134 74230 111218
rect 73910 110898 73952 111134
rect 74188 110898 74230 111134
rect 73910 110866 74230 110898
rect 79840 111454 80160 111486
rect 79840 111218 79882 111454
rect 80118 111218 80160 111454
rect 79840 111134 80160 111218
rect 79840 110898 79882 111134
rect 80118 110898 80160 111134
rect 79840 110866 80160 110898
rect 85771 111454 86091 111486
rect 85771 111218 85813 111454
rect 86049 111218 86091 111454
rect 85771 111134 86091 111218
rect 85771 110898 85813 111134
rect 86049 110898 86091 111134
rect 85771 110866 86091 110898
rect 100910 111454 101230 111486
rect 100910 111218 100952 111454
rect 101188 111218 101230 111454
rect 100910 111134 101230 111218
rect 100910 110898 100952 111134
rect 101188 110898 101230 111134
rect 100910 110866 101230 110898
rect 106840 111454 107160 111486
rect 106840 111218 106882 111454
rect 107118 111218 107160 111454
rect 106840 111134 107160 111218
rect 106840 110898 106882 111134
rect 107118 110898 107160 111134
rect 106840 110866 107160 110898
rect 112771 111454 113091 111486
rect 112771 111218 112813 111454
rect 113049 111218 113091 111454
rect 112771 111134 113091 111218
rect 112771 110898 112813 111134
rect 113049 110898 113091 111134
rect 112771 110866 113091 110898
rect 127910 111454 128230 111486
rect 127910 111218 127952 111454
rect 128188 111218 128230 111454
rect 127910 111134 128230 111218
rect 127910 110898 127952 111134
rect 128188 110898 128230 111134
rect 127910 110866 128230 110898
rect 133840 111454 134160 111486
rect 133840 111218 133882 111454
rect 134118 111218 134160 111454
rect 133840 111134 134160 111218
rect 133840 110898 133882 111134
rect 134118 110898 134160 111134
rect 133840 110866 134160 110898
rect 139771 111454 140091 111486
rect 139771 111218 139813 111454
rect 140049 111218 140091 111454
rect 139771 111134 140091 111218
rect 139771 110898 139813 111134
rect 140049 110898 140091 111134
rect 139771 110866 140091 110898
rect 154910 111454 155230 111486
rect 154910 111218 154952 111454
rect 155188 111218 155230 111454
rect 154910 111134 155230 111218
rect 154910 110898 154952 111134
rect 155188 110898 155230 111134
rect 154910 110866 155230 110898
rect 160840 111454 161160 111486
rect 160840 111218 160882 111454
rect 161118 111218 161160 111454
rect 160840 111134 161160 111218
rect 160840 110898 160882 111134
rect 161118 110898 161160 111134
rect 160840 110866 161160 110898
rect 166771 111454 167091 111486
rect 166771 111218 166813 111454
rect 167049 111218 167091 111454
rect 166771 111134 167091 111218
rect 166771 110898 166813 111134
rect 167049 110898 167091 111134
rect 166771 110866 167091 110898
rect 181910 111454 182230 111486
rect 181910 111218 181952 111454
rect 182188 111218 182230 111454
rect 181910 111134 182230 111218
rect 181910 110898 181952 111134
rect 182188 110898 182230 111134
rect 181910 110866 182230 110898
rect 187840 111454 188160 111486
rect 187840 111218 187882 111454
rect 188118 111218 188160 111454
rect 187840 111134 188160 111218
rect 187840 110898 187882 111134
rect 188118 110898 188160 111134
rect 187840 110866 188160 110898
rect 193771 111454 194091 111486
rect 193771 111218 193813 111454
rect 194049 111218 194091 111454
rect 193771 111134 194091 111218
rect 193771 110898 193813 111134
rect 194049 110898 194091 111134
rect 193771 110866 194091 110898
rect 208910 111454 209230 111486
rect 208910 111218 208952 111454
rect 209188 111218 209230 111454
rect 208910 111134 209230 111218
rect 208910 110898 208952 111134
rect 209188 110898 209230 111134
rect 208910 110866 209230 110898
rect 214840 111454 215160 111486
rect 214840 111218 214882 111454
rect 215118 111218 215160 111454
rect 214840 111134 215160 111218
rect 214840 110898 214882 111134
rect 215118 110898 215160 111134
rect 214840 110866 215160 110898
rect 220771 111454 221091 111486
rect 220771 111218 220813 111454
rect 221049 111218 221091 111454
rect 220771 111134 221091 111218
rect 220771 110898 220813 111134
rect 221049 110898 221091 111134
rect 220771 110866 221091 110898
rect 235910 111454 236230 111486
rect 235910 111218 235952 111454
rect 236188 111218 236230 111454
rect 235910 111134 236230 111218
rect 235910 110898 235952 111134
rect 236188 110898 236230 111134
rect 235910 110866 236230 110898
rect 241840 111454 242160 111486
rect 241840 111218 241882 111454
rect 242118 111218 242160 111454
rect 241840 111134 242160 111218
rect 241840 110898 241882 111134
rect 242118 110898 242160 111134
rect 241840 110866 242160 110898
rect 247771 111454 248091 111486
rect 247771 111218 247813 111454
rect 248049 111218 248091 111454
rect 247771 111134 248091 111218
rect 247771 110898 247813 111134
rect 248049 110898 248091 111134
rect 247771 110866 248091 110898
rect 262910 111454 263230 111486
rect 262910 111218 262952 111454
rect 263188 111218 263230 111454
rect 262910 111134 263230 111218
rect 262910 110898 262952 111134
rect 263188 110898 263230 111134
rect 262910 110866 263230 110898
rect 268840 111454 269160 111486
rect 268840 111218 268882 111454
rect 269118 111218 269160 111454
rect 268840 111134 269160 111218
rect 268840 110898 268882 111134
rect 269118 110898 269160 111134
rect 268840 110866 269160 110898
rect 274771 111454 275091 111486
rect 274771 111218 274813 111454
rect 275049 111218 275091 111454
rect 274771 111134 275091 111218
rect 274771 110898 274813 111134
rect 275049 110898 275091 111134
rect 274771 110866 275091 110898
rect 289910 111454 290230 111486
rect 289910 111218 289952 111454
rect 290188 111218 290230 111454
rect 289910 111134 290230 111218
rect 289910 110898 289952 111134
rect 290188 110898 290230 111134
rect 289910 110866 290230 110898
rect 295840 111454 296160 111486
rect 295840 111218 295882 111454
rect 296118 111218 296160 111454
rect 295840 111134 296160 111218
rect 295840 110898 295882 111134
rect 296118 110898 296160 111134
rect 295840 110866 296160 110898
rect 301771 111454 302091 111486
rect 301771 111218 301813 111454
rect 302049 111218 302091 111454
rect 301771 111134 302091 111218
rect 301771 110898 301813 111134
rect 302049 110898 302091 111134
rect 301771 110866 302091 110898
rect 316910 111454 317230 111486
rect 316910 111218 316952 111454
rect 317188 111218 317230 111454
rect 316910 111134 317230 111218
rect 316910 110898 316952 111134
rect 317188 110898 317230 111134
rect 316910 110866 317230 110898
rect 322840 111454 323160 111486
rect 322840 111218 322882 111454
rect 323118 111218 323160 111454
rect 322840 111134 323160 111218
rect 322840 110898 322882 111134
rect 323118 110898 323160 111134
rect 322840 110866 323160 110898
rect 328771 111454 329091 111486
rect 328771 111218 328813 111454
rect 329049 111218 329091 111454
rect 328771 111134 329091 111218
rect 328771 110898 328813 111134
rect 329049 110898 329091 111134
rect 328771 110866 329091 110898
rect 343910 111454 344230 111486
rect 343910 111218 343952 111454
rect 344188 111218 344230 111454
rect 343910 111134 344230 111218
rect 343910 110898 343952 111134
rect 344188 110898 344230 111134
rect 343910 110866 344230 110898
rect 349840 111454 350160 111486
rect 349840 111218 349882 111454
rect 350118 111218 350160 111454
rect 349840 111134 350160 111218
rect 349840 110898 349882 111134
rect 350118 110898 350160 111134
rect 349840 110866 350160 110898
rect 355771 111454 356091 111486
rect 355771 111218 355813 111454
rect 356049 111218 356091 111454
rect 355771 111134 356091 111218
rect 355771 110898 355813 111134
rect 356049 110898 356091 111134
rect 355771 110866 356091 110898
rect 370910 111454 371230 111486
rect 370910 111218 370952 111454
rect 371188 111218 371230 111454
rect 370910 111134 371230 111218
rect 370910 110898 370952 111134
rect 371188 110898 371230 111134
rect 370910 110866 371230 110898
rect 376840 111454 377160 111486
rect 376840 111218 376882 111454
rect 377118 111218 377160 111454
rect 376840 111134 377160 111218
rect 376840 110898 376882 111134
rect 377118 110898 377160 111134
rect 376840 110866 377160 110898
rect 382771 111454 383091 111486
rect 382771 111218 382813 111454
rect 383049 111218 383091 111454
rect 382771 111134 383091 111218
rect 382771 110898 382813 111134
rect 383049 110898 383091 111134
rect 382771 110866 383091 110898
rect 397910 111454 398230 111486
rect 397910 111218 397952 111454
rect 398188 111218 398230 111454
rect 397910 111134 398230 111218
rect 397910 110898 397952 111134
rect 398188 110898 398230 111134
rect 397910 110866 398230 110898
rect 403840 111454 404160 111486
rect 403840 111218 403882 111454
rect 404118 111218 404160 111454
rect 403840 111134 404160 111218
rect 403840 110898 403882 111134
rect 404118 110898 404160 111134
rect 403840 110866 404160 110898
rect 409771 111454 410091 111486
rect 409771 111218 409813 111454
rect 410049 111218 410091 111454
rect 409771 111134 410091 111218
rect 409771 110898 409813 111134
rect 410049 110898 410091 111134
rect 409771 110866 410091 110898
rect 424910 111454 425230 111486
rect 424910 111218 424952 111454
rect 425188 111218 425230 111454
rect 424910 111134 425230 111218
rect 424910 110898 424952 111134
rect 425188 110898 425230 111134
rect 424910 110866 425230 110898
rect 430840 111454 431160 111486
rect 430840 111218 430882 111454
rect 431118 111218 431160 111454
rect 430840 111134 431160 111218
rect 430840 110898 430882 111134
rect 431118 110898 431160 111134
rect 430840 110866 431160 110898
rect 436771 111454 437091 111486
rect 436771 111218 436813 111454
rect 437049 111218 437091 111454
rect 436771 111134 437091 111218
rect 436771 110898 436813 111134
rect 437049 110898 437091 111134
rect 436771 110866 437091 110898
rect 451910 111454 452230 111486
rect 451910 111218 451952 111454
rect 452188 111218 452230 111454
rect 451910 111134 452230 111218
rect 451910 110898 451952 111134
rect 452188 110898 452230 111134
rect 451910 110866 452230 110898
rect 457840 111454 458160 111486
rect 457840 111218 457882 111454
rect 458118 111218 458160 111454
rect 457840 111134 458160 111218
rect 457840 110898 457882 111134
rect 458118 110898 458160 111134
rect 457840 110866 458160 110898
rect 463771 111454 464091 111486
rect 463771 111218 463813 111454
rect 464049 111218 464091 111454
rect 463771 111134 464091 111218
rect 463771 110898 463813 111134
rect 464049 110898 464091 111134
rect 463771 110866 464091 110898
rect 478910 111454 479230 111486
rect 478910 111218 478952 111454
rect 479188 111218 479230 111454
rect 478910 111134 479230 111218
rect 478910 110898 478952 111134
rect 479188 110898 479230 111134
rect 478910 110866 479230 110898
rect 484840 111454 485160 111486
rect 484840 111218 484882 111454
rect 485118 111218 485160 111454
rect 484840 111134 485160 111218
rect 484840 110898 484882 111134
rect 485118 110898 485160 111134
rect 484840 110866 485160 110898
rect 490771 111454 491091 111486
rect 490771 111218 490813 111454
rect 491049 111218 491091 111454
rect 490771 111134 491091 111218
rect 490771 110898 490813 111134
rect 491049 110898 491091 111134
rect 490771 110866 491091 110898
rect 505910 111454 506230 111486
rect 505910 111218 505952 111454
rect 506188 111218 506230 111454
rect 505910 111134 506230 111218
rect 505910 110898 505952 111134
rect 506188 110898 506230 111134
rect 505910 110866 506230 110898
rect 511840 111454 512160 111486
rect 511840 111218 511882 111454
rect 512118 111218 512160 111454
rect 511840 111134 512160 111218
rect 511840 110898 511882 111134
rect 512118 110898 512160 111134
rect 511840 110866 512160 110898
rect 517771 111454 518091 111486
rect 517771 111218 517813 111454
rect 518049 111218 518091 111454
rect 517771 111134 518091 111218
rect 517771 110898 517813 111134
rect 518049 110898 518091 111134
rect 517771 110866 518091 110898
rect 532910 111454 533230 111486
rect 532910 111218 532952 111454
rect 533188 111218 533230 111454
rect 532910 111134 533230 111218
rect 532910 110898 532952 111134
rect 533188 110898 533230 111134
rect 532910 110866 533230 110898
rect 538840 111454 539160 111486
rect 538840 111218 538882 111454
rect 539118 111218 539160 111454
rect 538840 111134 539160 111218
rect 538840 110898 538882 111134
rect 539118 110898 539160 111134
rect 538840 110866 539160 110898
rect 544771 111454 545091 111486
rect 544771 111218 544813 111454
rect 545049 111218 545091 111454
rect 544771 111134 545091 111218
rect 544771 110898 544813 111134
rect 545049 110898 545091 111134
rect 544771 110866 545091 110898
rect 559794 111454 560414 128898
rect 559794 111218 559826 111454
rect 560062 111218 560146 111454
rect 560382 111218 560414 111454
rect 559794 111134 560414 111218
rect 559794 110898 559826 111134
rect 560062 110898 560146 111134
rect 560382 110898 560414 111134
rect 10794 102218 10826 102454
rect 11062 102218 11146 102454
rect 11382 102218 11414 102454
rect 10794 102134 11414 102218
rect 10794 101898 10826 102134
rect 11062 101898 11146 102134
rect 11382 101898 11414 102134
rect 10794 84454 11414 101898
rect 22874 102454 23194 102486
rect 22874 102218 22916 102454
rect 23152 102218 23194 102454
rect 22874 102134 23194 102218
rect 22874 101898 22916 102134
rect 23152 101898 23194 102134
rect 22874 101866 23194 101898
rect 28805 102454 29125 102486
rect 28805 102218 28847 102454
rect 29083 102218 29125 102454
rect 28805 102134 29125 102218
rect 28805 101898 28847 102134
rect 29083 101898 29125 102134
rect 28805 101866 29125 101898
rect 49874 102454 50194 102486
rect 49874 102218 49916 102454
rect 50152 102218 50194 102454
rect 49874 102134 50194 102218
rect 49874 101898 49916 102134
rect 50152 101898 50194 102134
rect 49874 101866 50194 101898
rect 55805 102454 56125 102486
rect 55805 102218 55847 102454
rect 56083 102218 56125 102454
rect 55805 102134 56125 102218
rect 55805 101898 55847 102134
rect 56083 101898 56125 102134
rect 55805 101866 56125 101898
rect 76874 102454 77194 102486
rect 76874 102218 76916 102454
rect 77152 102218 77194 102454
rect 76874 102134 77194 102218
rect 76874 101898 76916 102134
rect 77152 101898 77194 102134
rect 76874 101866 77194 101898
rect 82805 102454 83125 102486
rect 82805 102218 82847 102454
rect 83083 102218 83125 102454
rect 82805 102134 83125 102218
rect 82805 101898 82847 102134
rect 83083 101898 83125 102134
rect 82805 101866 83125 101898
rect 103874 102454 104194 102486
rect 103874 102218 103916 102454
rect 104152 102218 104194 102454
rect 103874 102134 104194 102218
rect 103874 101898 103916 102134
rect 104152 101898 104194 102134
rect 103874 101866 104194 101898
rect 109805 102454 110125 102486
rect 109805 102218 109847 102454
rect 110083 102218 110125 102454
rect 109805 102134 110125 102218
rect 109805 101898 109847 102134
rect 110083 101898 110125 102134
rect 109805 101866 110125 101898
rect 130874 102454 131194 102486
rect 130874 102218 130916 102454
rect 131152 102218 131194 102454
rect 130874 102134 131194 102218
rect 130874 101898 130916 102134
rect 131152 101898 131194 102134
rect 130874 101866 131194 101898
rect 136805 102454 137125 102486
rect 136805 102218 136847 102454
rect 137083 102218 137125 102454
rect 136805 102134 137125 102218
rect 136805 101898 136847 102134
rect 137083 101898 137125 102134
rect 136805 101866 137125 101898
rect 157874 102454 158194 102486
rect 157874 102218 157916 102454
rect 158152 102218 158194 102454
rect 157874 102134 158194 102218
rect 157874 101898 157916 102134
rect 158152 101898 158194 102134
rect 157874 101866 158194 101898
rect 163805 102454 164125 102486
rect 163805 102218 163847 102454
rect 164083 102218 164125 102454
rect 163805 102134 164125 102218
rect 163805 101898 163847 102134
rect 164083 101898 164125 102134
rect 163805 101866 164125 101898
rect 184874 102454 185194 102486
rect 184874 102218 184916 102454
rect 185152 102218 185194 102454
rect 184874 102134 185194 102218
rect 184874 101898 184916 102134
rect 185152 101898 185194 102134
rect 184874 101866 185194 101898
rect 190805 102454 191125 102486
rect 190805 102218 190847 102454
rect 191083 102218 191125 102454
rect 190805 102134 191125 102218
rect 190805 101898 190847 102134
rect 191083 101898 191125 102134
rect 190805 101866 191125 101898
rect 211874 102454 212194 102486
rect 211874 102218 211916 102454
rect 212152 102218 212194 102454
rect 211874 102134 212194 102218
rect 211874 101898 211916 102134
rect 212152 101898 212194 102134
rect 211874 101866 212194 101898
rect 217805 102454 218125 102486
rect 217805 102218 217847 102454
rect 218083 102218 218125 102454
rect 217805 102134 218125 102218
rect 217805 101898 217847 102134
rect 218083 101898 218125 102134
rect 217805 101866 218125 101898
rect 238874 102454 239194 102486
rect 238874 102218 238916 102454
rect 239152 102218 239194 102454
rect 238874 102134 239194 102218
rect 238874 101898 238916 102134
rect 239152 101898 239194 102134
rect 238874 101866 239194 101898
rect 244805 102454 245125 102486
rect 244805 102218 244847 102454
rect 245083 102218 245125 102454
rect 244805 102134 245125 102218
rect 244805 101898 244847 102134
rect 245083 101898 245125 102134
rect 244805 101866 245125 101898
rect 265874 102454 266194 102486
rect 265874 102218 265916 102454
rect 266152 102218 266194 102454
rect 265874 102134 266194 102218
rect 265874 101898 265916 102134
rect 266152 101898 266194 102134
rect 265874 101866 266194 101898
rect 271805 102454 272125 102486
rect 271805 102218 271847 102454
rect 272083 102218 272125 102454
rect 271805 102134 272125 102218
rect 271805 101898 271847 102134
rect 272083 101898 272125 102134
rect 271805 101866 272125 101898
rect 292874 102454 293194 102486
rect 292874 102218 292916 102454
rect 293152 102218 293194 102454
rect 292874 102134 293194 102218
rect 292874 101898 292916 102134
rect 293152 101898 293194 102134
rect 292874 101866 293194 101898
rect 298805 102454 299125 102486
rect 298805 102218 298847 102454
rect 299083 102218 299125 102454
rect 298805 102134 299125 102218
rect 298805 101898 298847 102134
rect 299083 101898 299125 102134
rect 298805 101866 299125 101898
rect 319874 102454 320194 102486
rect 319874 102218 319916 102454
rect 320152 102218 320194 102454
rect 319874 102134 320194 102218
rect 319874 101898 319916 102134
rect 320152 101898 320194 102134
rect 319874 101866 320194 101898
rect 325805 102454 326125 102486
rect 325805 102218 325847 102454
rect 326083 102218 326125 102454
rect 325805 102134 326125 102218
rect 325805 101898 325847 102134
rect 326083 101898 326125 102134
rect 325805 101866 326125 101898
rect 346874 102454 347194 102486
rect 346874 102218 346916 102454
rect 347152 102218 347194 102454
rect 346874 102134 347194 102218
rect 346874 101898 346916 102134
rect 347152 101898 347194 102134
rect 346874 101866 347194 101898
rect 352805 102454 353125 102486
rect 352805 102218 352847 102454
rect 353083 102218 353125 102454
rect 352805 102134 353125 102218
rect 352805 101898 352847 102134
rect 353083 101898 353125 102134
rect 352805 101866 353125 101898
rect 373874 102454 374194 102486
rect 373874 102218 373916 102454
rect 374152 102218 374194 102454
rect 373874 102134 374194 102218
rect 373874 101898 373916 102134
rect 374152 101898 374194 102134
rect 373874 101866 374194 101898
rect 379805 102454 380125 102486
rect 379805 102218 379847 102454
rect 380083 102218 380125 102454
rect 379805 102134 380125 102218
rect 379805 101898 379847 102134
rect 380083 101898 380125 102134
rect 379805 101866 380125 101898
rect 400874 102454 401194 102486
rect 400874 102218 400916 102454
rect 401152 102218 401194 102454
rect 400874 102134 401194 102218
rect 400874 101898 400916 102134
rect 401152 101898 401194 102134
rect 400874 101866 401194 101898
rect 406805 102454 407125 102486
rect 406805 102218 406847 102454
rect 407083 102218 407125 102454
rect 406805 102134 407125 102218
rect 406805 101898 406847 102134
rect 407083 101898 407125 102134
rect 406805 101866 407125 101898
rect 427874 102454 428194 102486
rect 427874 102218 427916 102454
rect 428152 102218 428194 102454
rect 427874 102134 428194 102218
rect 427874 101898 427916 102134
rect 428152 101898 428194 102134
rect 427874 101866 428194 101898
rect 433805 102454 434125 102486
rect 433805 102218 433847 102454
rect 434083 102218 434125 102454
rect 433805 102134 434125 102218
rect 433805 101898 433847 102134
rect 434083 101898 434125 102134
rect 433805 101866 434125 101898
rect 454874 102454 455194 102486
rect 454874 102218 454916 102454
rect 455152 102218 455194 102454
rect 454874 102134 455194 102218
rect 454874 101898 454916 102134
rect 455152 101898 455194 102134
rect 454874 101866 455194 101898
rect 460805 102454 461125 102486
rect 460805 102218 460847 102454
rect 461083 102218 461125 102454
rect 460805 102134 461125 102218
rect 460805 101898 460847 102134
rect 461083 101898 461125 102134
rect 460805 101866 461125 101898
rect 481874 102454 482194 102486
rect 481874 102218 481916 102454
rect 482152 102218 482194 102454
rect 481874 102134 482194 102218
rect 481874 101898 481916 102134
rect 482152 101898 482194 102134
rect 481874 101866 482194 101898
rect 487805 102454 488125 102486
rect 487805 102218 487847 102454
rect 488083 102218 488125 102454
rect 487805 102134 488125 102218
rect 487805 101898 487847 102134
rect 488083 101898 488125 102134
rect 487805 101866 488125 101898
rect 508874 102454 509194 102486
rect 508874 102218 508916 102454
rect 509152 102218 509194 102454
rect 508874 102134 509194 102218
rect 508874 101898 508916 102134
rect 509152 101898 509194 102134
rect 508874 101866 509194 101898
rect 514805 102454 515125 102486
rect 514805 102218 514847 102454
rect 515083 102218 515125 102454
rect 514805 102134 515125 102218
rect 514805 101898 514847 102134
rect 515083 101898 515125 102134
rect 514805 101866 515125 101898
rect 535874 102454 536194 102486
rect 535874 102218 535916 102454
rect 536152 102218 536194 102454
rect 535874 102134 536194 102218
rect 535874 101898 535916 102134
rect 536152 101898 536194 102134
rect 535874 101866 536194 101898
rect 541805 102454 542125 102486
rect 541805 102218 541847 102454
rect 542083 102218 542125 102454
rect 541805 102134 542125 102218
rect 541805 101898 541847 102134
rect 542083 101898 542125 102134
rect 541805 101866 542125 101898
rect 19794 93454 20414 95000
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 92000 20414 92898
rect 28794 94394 29414 95000
rect 28794 94158 28826 94394
rect 29062 94158 29146 94394
rect 29382 94158 29414 94394
rect 28794 94074 29414 94158
rect 28794 93838 28826 94074
rect 29062 93838 29146 94074
rect 29382 93838 29414 94074
rect 28794 92000 29414 93838
rect 37794 93454 38414 95000
rect 37794 93218 37826 93454
rect 38062 93218 38146 93454
rect 38382 93218 38414 93454
rect 37794 93134 38414 93218
rect 37794 92898 37826 93134
rect 38062 92898 38146 93134
rect 38382 92898 38414 93134
rect 37794 92000 38414 92898
rect 46794 94394 47414 95000
rect 46794 94158 46826 94394
rect 47062 94158 47146 94394
rect 47382 94158 47414 94394
rect 46794 94074 47414 94158
rect 46794 93838 46826 94074
rect 47062 93838 47146 94074
rect 47382 93838 47414 94074
rect 46794 92000 47414 93838
rect 55794 93454 56414 95000
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 92000 56414 92898
rect 64794 94394 65414 95000
rect 64794 94158 64826 94394
rect 65062 94158 65146 94394
rect 65382 94158 65414 94394
rect 64794 94074 65414 94158
rect 64794 93838 64826 94074
rect 65062 93838 65146 94074
rect 65382 93838 65414 94074
rect 64794 92000 65414 93838
rect 73794 93454 74414 95000
rect 73794 93218 73826 93454
rect 74062 93218 74146 93454
rect 74382 93218 74414 93454
rect 73794 93134 74414 93218
rect 73794 92898 73826 93134
rect 74062 92898 74146 93134
rect 74382 92898 74414 93134
rect 73794 92000 74414 92898
rect 82794 94394 83414 95000
rect 82794 94158 82826 94394
rect 83062 94158 83146 94394
rect 83382 94158 83414 94394
rect 82794 94074 83414 94158
rect 82794 93838 82826 94074
rect 83062 93838 83146 94074
rect 83382 93838 83414 94074
rect 82794 92000 83414 93838
rect 91794 93454 92414 95000
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 92000 92414 92898
rect 100794 94394 101414 95000
rect 100794 94158 100826 94394
rect 101062 94158 101146 94394
rect 101382 94158 101414 94394
rect 100794 94074 101414 94158
rect 100794 93838 100826 94074
rect 101062 93838 101146 94074
rect 101382 93838 101414 94074
rect 100794 92000 101414 93838
rect 109794 93454 110414 95000
rect 109794 93218 109826 93454
rect 110062 93218 110146 93454
rect 110382 93218 110414 93454
rect 109794 93134 110414 93218
rect 109794 92898 109826 93134
rect 110062 92898 110146 93134
rect 110382 92898 110414 93134
rect 109794 92000 110414 92898
rect 118794 94394 119414 95000
rect 118794 94158 118826 94394
rect 119062 94158 119146 94394
rect 119382 94158 119414 94394
rect 118794 94074 119414 94158
rect 118794 93838 118826 94074
rect 119062 93838 119146 94074
rect 119382 93838 119414 94074
rect 118794 92000 119414 93838
rect 127794 93454 128414 95000
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 92000 128414 92898
rect 136794 94394 137414 95000
rect 136794 94158 136826 94394
rect 137062 94158 137146 94394
rect 137382 94158 137414 94394
rect 136794 94074 137414 94158
rect 136794 93838 136826 94074
rect 137062 93838 137146 94074
rect 137382 93838 137414 94074
rect 136794 92000 137414 93838
rect 145794 93454 146414 95000
rect 145794 93218 145826 93454
rect 146062 93218 146146 93454
rect 146382 93218 146414 93454
rect 145794 93134 146414 93218
rect 145794 92898 145826 93134
rect 146062 92898 146146 93134
rect 146382 92898 146414 93134
rect 145794 92000 146414 92898
rect 154794 94394 155414 95000
rect 154794 94158 154826 94394
rect 155062 94158 155146 94394
rect 155382 94158 155414 94394
rect 154794 94074 155414 94158
rect 154794 93838 154826 94074
rect 155062 93838 155146 94074
rect 155382 93838 155414 94074
rect 154794 92000 155414 93838
rect 163794 93454 164414 95000
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 92000 164414 92898
rect 172794 94394 173414 95000
rect 172794 94158 172826 94394
rect 173062 94158 173146 94394
rect 173382 94158 173414 94394
rect 172794 94074 173414 94158
rect 172794 93838 172826 94074
rect 173062 93838 173146 94074
rect 173382 93838 173414 94074
rect 172794 92000 173414 93838
rect 181794 93454 182414 95000
rect 181794 93218 181826 93454
rect 182062 93218 182146 93454
rect 182382 93218 182414 93454
rect 181794 93134 182414 93218
rect 181794 92898 181826 93134
rect 182062 92898 182146 93134
rect 182382 92898 182414 93134
rect 181794 92000 182414 92898
rect 190794 94394 191414 95000
rect 190794 94158 190826 94394
rect 191062 94158 191146 94394
rect 191382 94158 191414 94394
rect 190794 94074 191414 94158
rect 190794 93838 190826 94074
rect 191062 93838 191146 94074
rect 191382 93838 191414 94074
rect 190794 92000 191414 93838
rect 199794 93454 200414 95000
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 92000 200414 92898
rect 208794 94394 209414 95000
rect 208794 94158 208826 94394
rect 209062 94158 209146 94394
rect 209382 94158 209414 94394
rect 208794 94074 209414 94158
rect 208794 93838 208826 94074
rect 209062 93838 209146 94074
rect 209382 93838 209414 94074
rect 208794 92000 209414 93838
rect 217794 93454 218414 95000
rect 217794 93218 217826 93454
rect 218062 93218 218146 93454
rect 218382 93218 218414 93454
rect 217794 93134 218414 93218
rect 217794 92898 217826 93134
rect 218062 92898 218146 93134
rect 218382 92898 218414 93134
rect 217794 92000 218414 92898
rect 226794 94394 227414 95000
rect 226794 94158 226826 94394
rect 227062 94158 227146 94394
rect 227382 94158 227414 94394
rect 226794 94074 227414 94158
rect 226794 93838 226826 94074
rect 227062 93838 227146 94074
rect 227382 93838 227414 94074
rect 226794 92000 227414 93838
rect 235794 93454 236414 95000
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 92000 236414 92898
rect 244794 94394 245414 95000
rect 244794 94158 244826 94394
rect 245062 94158 245146 94394
rect 245382 94158 245414 94394
rect 244794 94074 245414 94158
rect 244794 93838 244826 94074
rect 245062 93838 245146 94074
rect 245382 93838 245414 94074
rect 244794 92000 245414 93838
rect 253794 93454 254414 95000
rect 253794 93218 253826 93454
rect 254062 93218 254146 93454
rect 254382 93218 254414 93454
rect 253794 93134 254414 93218
rect 253794 92898 253826 93134
rect 254062 92898 254146 93134
rect 254382 92898 254414 93134
rect 253794 92000 254414 92898
rect 262794 94394 263414 95000
rect 262794 94158 262826 94394
rect 263062 94158 263146 94394
rect 263382 94158 263414 94394
rect 262794 94074 263414 94158
rect 262794 93838 262826 94074
rect 263062 93838 263146 94074
rect 263382 93838 263414 94074
rect 262794 92000 263414 93838
rect 271794 93454 272414 95000
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 92000 272414 92898
rect 280794 94394 281414 95000
rect 280794 94158 280826 94394
rect 281062 94158 281146 94394
rect 281382 94158 281414 94394
rect 280794 94074 281414 94158
rect 280794 93838 280826 94074
rect 281062 93838 281146 94074
rect 281382 93838 281414 94074
rect 280794 92000 281414 93838
rect 289794 93454 290414 95000
rect 289794 93218 289826 93454
rect 290062 93218 290146 93454
rect 290382 93218 290414 93454
rect 289794 93134 290414 93218
rect 289794 92898 289826 93134
rect 290062 92898 290146 93134
rect 290382 92898 290414 93134
rect 289794 92000 290414 92898
rect 298794 94394 299414 95000
rect 298794 94158 298826 94394
rect 299062 94158 299146 94394
rect 299382 94158 299414 94394
rect 298794 94074 299414 94158
rect 298794 93838 298826 94074
rect 299062 93838 299146 94074
rect 299382 93838 299414 94074
rect 298794 92000 299414 93838
rect 307794 93454 308414 95000
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 92000 308414 92898
rect 316794 94394 317414 95000
rect 316794 94158 316826 94394
rect 317062 94158 317146 94394
rect 317382 94158 317414 94394
rect 316794 94074 317414 94158
rect 316794 93838 316826 94074
rect 317062 93838 317146 94074
rect 317382 93838 317414 94074
rect 316794 92000 317414 93838
rect 325794 93454 326414 95000
rect 325794 93218 325826 93454
rect 326062 93218 326146 93454
rect 326382 93218 326414 93454
rect 325794 93134 326414 93218
rect 325794 92898 325826 93134
rect 326062 92898 326146 93134
rect 326382 92898 326414 93134
rect 325794 92000 326414 92898
rect 334794 94394 335414 95000
rect 334794 94158 334826 94394
rect 335062 94158 335146 94394
rect 335382 94158 335414 94394
rect 334794 94074 335414 94158
rect 334794 93838 334826 94074
rect 335062 93838 335146 94074
rect 335382 93838 335414 94074
rect 334794 92000 335414 93838
rect 343794 93454 344414 95000
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 92000 344414 92898
rect 352794 94394 353414 95000
rect 352794 94158 352826 94394
rect 353062 94158 353146 94394
rect 353382 94158 353414 94394
rect 352794 94074 353414 94158
rect 352794 93838 352826 94074
rect 353062 93838 353146 94074
rect 353382 93838 353414 94074
rect 352794 92000 353414 93838
rect 361794 93454 362414 95000
rect 361794 93218 361826 93454
rect 362062 93218 362146 93454
rect 362382 93218 362414 93454
rect 361794 93134 362414 93218
rect 361794 92898 361826 93134
rect 362062 92898 362146 93134
rect 362382 92898 362414 93134
rect 361794 92000 362414 92898
rect 370794 94394 371414 95000
rect 370794 94158 370826 94394
rect 371062 94158 371146 94394
rect 371382 94158 371414 94394
rect 370794 94074 371414 94158
rect 370794 93838 370826 94074
rect 371062 93838 371146 94074
rect 371382 93838 371414 94074
rect 370794 92000 371414 93838
rect 379794 93454 380414 95000
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 92000 380414 92898
rect 388794 94394 389414 95000
rect 388794 94158 388826 94394
rect 389062 94158 389146 94394
rect 389382 94158 389414 94394
rect 388794 94074 389414 94158
rect 388794 93838 388826 94074
rect 389062 93838 389146 94074
rect 389382 93838 389414 94074
rect 388794 92000 389414 93838
rect 397794 93454 398414 95000
rect 397794 93218 397826 93454
rect 398062 93218 398146 93454
rect 398382 93218 398414 93454
rect 397794 93134 398414 93218
rect 397794 92898 397826 93134
rect 398062 92898 398146 93134
rect 398382 92898 398414 93134
rect 397794 92000 398414 92898
rect 406794 94394 407414 95000
rect 406794 94158 406826 94394
rect 407062 94158 407146 94394
rect 407382 94158 407414 94394
rect 406794 94074 407414 94158
rect 406794 93838 406826 94074
rect 407062 93838 407146 94074
rect 407382 93838 407414 94074
rect 406794 92000 407414 93838
rect 415794 93454 416414 95000
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 92000 416414 92898
rect 424794 94394 425414 95000
rect 424794 94158 424826 94394
rect 425062 94158 425146 94394
rect 425382 94158 425414 94394
rect 424794 94074 425414 94158
rect 424794 93838 424826 94074
rect 425062 93838 425146 94074
rect 425382 93838 425414 94074
rect 424794 92000 425414 93838
rect 433794 93454 434414 95000
rect 433794 93218 433826 93454
rect 434062 93218 434146 93454
rect 434382 93218 434414 93454
rect 433794 93134 434414 93218
rect 433794 92898 433826 93134
rect 434062 92898 434146 93134
rect 434382 92898 434414 93134
rect 433794 92000 434414 92898
rect 442794 94394 443414 95000
rect 442794 94158 442826 94394
rect 443062 94158 443146 94394
rect 443382 94158 443414 94394
rect 442794 94074 443414 94158
rect 442794 93838 442826 94074
rect 443062 93838 443146 94074
rect 443382 93838 443414 94074
rect 442794 92000 443414 93838
rect 451794 93454 452414 95000
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 92000 452414 92898
rect 460794 94394 461414 95000
rect 460794 94158 460826 94394
rect 461062 94158 461146 94394
rect 461382 94158 461414 94394
rect 460794 94074 461414 94158
rect 460794 93838 460826 94074
rect 461062 93838 461146 94074
rect 461382 93838 461414 94074
rect 460794 92000 461414 93838
rect 469794 93454 470414 95000
rect 469794 93218 469826 93454
rect 470062 93218 470146 93454
rect 470382 93218 470414 93454
rect 469794 93134 470414 93218
rect 469794 92898 469826 93134
rect 470062 92898 470146 93134
rect 470382 92898 470414 93134
rect 469794 92000 470414 92898
rect 478794 94394 479414 95000
rect 478794 94158 478826 94394
rect 479062 94158 479146 94394
rect 479382 94158 479414 94394
rect 478794 94074 479414 94158
rect 478794 93838 478826 94074
rect 479062 93838 479146 94074
rect 479382 93838 479414 94074
rect 478794 92000 479414 93838
rect 487794 93454 488414 95000
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 92000 488414 92898
rect 496794 94394 497414 95000
rect 496794 94158 496826 94394
rect 497062 94158 497146 94394
rect 497382 94158 497414 94394
rect 496794 94074 497414 94158
rect 496794 93838 496826 94074
rect 497062 93838 497146 94074
rect 497382 93838 497414 94074
rect 496794 92000 497414 93838
rect 505794 93454 506414 95000
rect 505794 93218 505826 93454
rect 506062 93218 506146 93454
rect 506382 93218 506414 93454
rect 505794 93134 506414 93218
rect 505794 92898 505826 93134
rect 506062 92898 506146 93134
rect 506382 92898 506414 93134
rect 505794 92000 506414 92898
rect 514794 94394 515414 95000
rect 514794 94158 514826 94394
rect 515062 94158 515146 94394
rect 515382 94158 515414 94394
rect 514794 94074 515414 94158
rect 514794 93838 514826 94074
rect 515062 93838 515146 94074
rect 515382 93838 515414 94074
rect 514794 92000 515414 93838
rect 523794 93454 524414 95000
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 92000 524414 92898
rect 532794 94394 533414 95000
rect 532794 94158 532826 94394
rect 533062 94158 533146 94394
rect 533382 94158 533414 94394
rect 532794 94074 533414 94158
rect 532794 93838 532826 94074
rect 533062 93838 533146 94074
rect 533382 93838 533414 94074
rect 532794 92000 533414 93838
rect 541794 93454 542414 95000
rect 541794 93218 541826 93454
rect 542062 93218 542146 93454
rect 542382 93218 542414 93454
rect 541794 93134 542414 93218
rect 541794 92898 541826 93134
rect 542062 92898 542146 93134
rect 542382 92898 542414 93134
rect 541794 92000 542414 92898
rect 550794 94394 551414 95000
rect 550794 94158 550826 94394
rect 551062 94158 551146 94394
rect 551382 94158 551414 94394
rect 550794 94074 551414 94158
rect 550794 93838 550826 94074
rect 551062 93838 551146 94074
rect 551382 93838 551414 94074
rect 550794 92000 551414 93838
rect 559794 93454 560414 110898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 66454 11414 83898
rect 22874 84454 23194 84486
rect 22874 84218 22916 84454
rect 23152 84218 23194 84454
rect 22874 84134 23194 84218
rect 22874 83898 22916 84134
rect 23152 83898 23194 84134
rect 22874 83866 23194 83898
rect 28805 84454 29125 84486
rect 28805 84218 28847 84454
rect 29083 84218 29125 84454
rect 28805 84134 29125 84218
rect 28805 83898 28847 84134
rect 29083 83898 29125 84134
rect 28805 83866 29125 83898
rect 49874 84454 50194 84486
rect 49874 84218 49916 84454
rect 50152 84218 50194 84454
rect 49874 84134 50194 84218
rect 49874 83898 49916 84134
rect 50152 83898 50194 84134
rect 49874 83866 50194 83898
rect 55805 84454 56125 84486
rect 55805 84218 55847 84454
rect 56083 84218 56125 84454
rect 55805 84134 56125 84218
rect 55805 83898 55847 84134
rect 56083 83898 56125 84134
rect 55805 83866 56125 83898
rect 76874 84454 77194 84486
rect 76874 84218 76916 84454
rect 77152 84218 77194 84454
rect 76874 84134 77194 84218
rect 76874 83898 76916 84134
rect 77152 83898 77194 84134
rect 76874 83866 77194 83898
rect 82805 84454 83125 84486
rect 82805 84218 82847 84454
rect 83083 84218 83125 84454
rect 82805 84134 83125 84218
rect 82805 83898 82847 84134
rect 83083 83898 83125 84134
rect 82805 83866 83125 83898
rect 103874 84454 104194 84486
rect 103874 84218 103916 84454
rect 104152 84218 104194 84454
rect 103874 84134 104194 84218
rect 103874 83898 103916 84134
rect 104152 83898 104194 84134
rect 103874 83866 104194 83898
rect 109805 84454 110125 84486
rect 109805 84218 109847 84454
rect 110083 84218 110125 84454
rect 109805 84134 110125 84218
rect 109805 83898 109847 84134
rect 110083 83898 110125 84134
rect 109805 83866 110125 83898
rect 130874 84454 131194 84486
rect 130874 84218 130916 84454
rect 131152 84218 131194 84454
rect 130874 84134 131194 84218
rect 130874 83898 130916 84134
rect 131152 83898 131194 84134
rect 130874 83866 131194 83898
rect 136805 84454 137125 84486
rect 136805 84218 136847 84454
rect 137083 84218 137125 84454
rect 136805 84134 137125 84218
rect 136805 83898 136847 84134
rect 137083 83898 137125 84134
rect 136805 83866 137125 83898
rect 157874 84454 158194 84486
rect 157874 84218 157916 84454
rect 158152 84218 158194 84454
rect 157874 84134 158194 84218
rect 157874 83898 157916 84134
rect 158152 83898 158194 84134
rect 157874 83866 158194 83898
rect 163805 84454 164125 84486
rect 163805 84218 163847 84454
rect 164083 84218 164125 84454
rect 163805 84134 164125 84218
rect 163805 83898 163847 84134
rect 164083 83898 164125 84134
rect 163805 83866 164125 83898
rect 184874 84454 185194 84486
rect 184874 84218 184916 84454
rect 185152 84218 185194 84454
rect 184874 84134 185194 84218
rect 184874 83898 184916 84134
rect 185152 83898 185194 84134
rect 184874 83866 185194 83898
rect 190805 84454 191125 84486
rect 190805 84218 190847 84454
rect 191083 84218 191125 84454
rect 190805 84134 191125 84218
rect 190805 83898 190847 84134
rect 191083 83898 191125 84134
rect 190805 83866 191125 83898
rect 211874 84454 212194 84486
rect 211874 84218 211916 84454
rect 212152 84218 212194 84454
rect 211874 84134 212194 84218
rect 211874 83898 211916 84134
rect 212152 83898 212194 84134
rect 211874 83866 212194 83898
rect 217805 84454 218125 84486
rect 217805 84218 217847 84454
rect 218083 84218 218125 84454
rect 217805 84134 218125 84218
rect 217805 83898 217847 84134
rect 218083 83898 218125 84134
rect 217805 83866 218125 83898
rect 238874 84454 239194 84486
rect 238874 84218 238916 84454
rect 239152 84218 239194 84454
rect 238874 84134 239194 84218
rect 238874 83898 238916 84134
rect 239152 83898 239194 84134
rect 238874 83866 239194 83898
rect 244805 84454 245125 84486
rect 244805 84218 244847 84454
rect 245083 84218 245125 84454
rect 244805 84134 245125 84218
rect 244805 83898 244847 84134
rect 245083 83898 245125 84134
rect 244805 83866 245125 83898
rect 265874 84454 266194 84486
rect 265874 84218 265916 84454
rect 266152 84218 266194 84454
rect 265874 84134 266194 84218
rect 265874 83898 265916 84134
rect 266152 83898 266194 84134
rect 265874 83866 266194 83898
rect 271805 84454 272125 84486
rect 271805 84218 271847 84454
rect 272083 84218 272125 84454
rect 271805 84134 272125 84218
rect 271805 83898 271847 84134
rect 272083 83898 272125 84134
rect 271805 83866 272125 83898
rect 292874 84454 293194 84486
rect 292874 84218 292916 84454
rect 293152 84218 293194 84454
rect 292874 84134 293194 84218
rect 292874 83898 292916 84134
rect 293152 83898 293194 84134
rect 292874 83866 293194 83898
rect 298805 84454 299125 84486
rect 298805 84218 298847 84454
rect 299083 84218 299125 84454
rect 298805 84134 299125 84218
rect 298805 83898 298847 84134
rect 299083 83898 299125 84134
rect 298805 83866 299125 83898
rect 319874 84454 320194 84486
rect 319874 84218 319916 84454
rect 320152 84218 320194 84454
rect 319874 84134 320194 84218
rect 319874 83898 319916 84134
rect 320152 83898 320194 84134
rect 319874 83866 320194 83898
rect 325805 84454 326125 84486
rect 325805 84218 325847 84454
rect 326083 84218 326125 84454
rect 325805 84134 326125 84218
rect 325805 83898 325847 84134
rect 326083 83898 326125 84134
rect 325805 83866 326125 83898
rect 346874 84454 347194 84486
rect 346874 84218 346916 84454
rect 347152 84218 347194 84454
rect 346874 84134 347194 84218
rect 346874 83898 346916 84134
rect 347152 83898 347194 84134
rect 346874 83866 347194 83898
rect 352805 84454 353125 84486
rect 352805 84218 352847 84454
rect 353083 84218 353125 84454
rect 352805 84134 353125 84218
rect 352805 83898 352847 84134
rect 353083 83898 353125 84134
rect 352805 83866 353125 83898
rect 373874 84454 374194 84486
rect 373874 84218 373916 84454
rect 374152 84218 374194 84454
rect 373874 84134 374194 84218
rect 373874 83898 373916 84134
rect 374152 83898 374194 84134
rect 373874 83866 374194 83898
rect 379805 84454 380125 84486
rect 379805 84218 379847 84454
rect 380083 84218 380125 84454
rect 379805 84134 380125 84218
rect 379805 83898 379847 84134
rect 380083 83898 380125 84134
rect 379805 83866 380125 83898
rect 400874 84454 401194 84486
rect 400874 84218 400916 84454
rect 401152 84218 401194 84454
rect 400874 84134 401194 84218
rect 400874 83898 400916 84134
rect 401152 83898 401194 84134
rect 400874 83866 401194 83898
rect 406805 84454 407125 84486
rect 406805 84218 406847 84454
rect 407083 84218 407125 84454
rect 406805 84134 407125 84218
rect 406805 83898 406847 84134
rect 407083 83898 407125 84134
rect 406805 83866 407125 83898
rect 427874 84454 428194 84486
rect 427874 84218 427916 84454
rect 428152 84218 428194 84454
rect 427874 84134 428194 84218
rect 427874 83898 427916 84134
rect 428152 83898 428194 84134
rect 427874 83866 428194 83898
rect 433805 84454 434125 84486
rect 433805 84218 433847 84454
rect 434083 84218 434125 84454
rect 433805 84134 434125 84218
rect 433805 83898 433847 84134
rect 434083 83898 434125 84134
rect 433805 83866 434125 83898
rect 454874 84454 455194 84486
rect 454874 84218 454916 84454
rect 455152 84218 455194 84454
rect 454874 84134 455194 84218
rect 454874 83898 454916 84134
rect 455152 83898 455194 84134
rect 454874 83866 455194 83898
rect 460805 84454 461125 84486
rect 460805 84218 460847 84454
rect 461083 84218 461125 84454
rect 460805 84134 461125 84218
rect 460805 83898 460847 84134
rect 461083 83898 461125 84134
rect 460805 83866 461125 83898
rect 481874 84454 482194 84486
rect 481874 84218 481916 84454
rect 482152 84218 482194 84454
rect 481874 84134 482194 84218
rect 481874 83898 481916 84134
rect 482152 83898 482194 84134
rect 481874 83866 482194 83898
rect 487805 84454 488125 84486
rect 487805 84218 487847 84454
rect 488083 84218 488125 84454
rect 487805 84134 488125 84218
rect 487805 83898 487847 84134
rect 488083 83898 488125 84134
rect 487805 83866 488125 83898
rect 508874 84454 509194 84486
rect 508874 84218 508916 84454
rect 509152 84218 509194 84454
rect 508874 84134 509194 84218
rect 508874 83898 508916 84134
rect 509152 83898 509194 84134
rect 508874 83866 509194 83898
rect 514805 84454 515125 84486
rect 514805 84218 514847 84454
rect 515083 84218 515125 84454
rect 514805 84134 515125 84218
rect 514805 83898 514847 84134
rect 515083 83898 515125 84134
rect 514805 83866 515125 83898
rect 535874 84454 536194 84486
rect 535874 84218 535916 84454
rect 536152 84218 536194 84454
rect 535874 84134 536194 84218
rect 535874 83898 535916 84134
rect 536152 83898 536194 84134
rect 535874 83866 536194 83898
rect 541805 84454 542125 84486
rect 541805 84218 541847 84454
rect 542083 84218 542125 84454
rect 541805 84134 542125 84218
rect 541805 83898 541847 84134
rect 542083 83898 542125 84134
rect 541805 83866 542125 83898
rect 19910 75454 20230 75486
rect 19910 75218 19952 75454
rect 20188 75218 20230 75454
rect 19910 75134 20230 75218
rect 19910 74898 19952 75134
rect 20188 74898 20230 75134
rect 19910 74866 20230 74898
rect 25840 75454 26160 75486
rect 25840 75218 25882 75454
rect 26118 75218 26160 75454
rect 25840 75134 26160 75218
rect 25840 74898 25882 75134
rect 26118 74898 26160 75134
rect 25840 74866 26160 74898
rect 31771 75454 32091 75486
rect 31771 75218 31813 75454
rect 32049 75218 32091 75454
rect 31771 75134 32091 75218
rect 31771 74898 31813 75134
rect 32049 74898 32091 75134
rect 31771 74866 32091 74898
rect 46910 75454 47230 75486
rect 46910 75218 46952 75454
rect 47188 75218 47230 75454
rect 46910 75134 47230 75218
rect 46910 74898 46952 75134
rect 47188 74898 47230 75134
rect 46910 74866 47230 74898
rect 52840 75454 53160 75486
rect 52840 75218 52882 75454
rect 53118 75218 53160 75454
rect 52840 75134 53160 75218
rect 52840 74898 52882 75134
rect 53118 74898 53160 75134
rect 52840 74866 53160 74898
rect 58771 75454 59091 75486
rect 58771 75218 58813 75454
rect 59049 75218 59091 75454
rect 58771 75134 59091 75218
rect 58771 74898 58813 75134
rect 59049 74898 59091 75134
rect 58771 74866 59091 74898
rect 73910 75454 74230 75486
rect 73910 75218 73952 75454
rect 74188 75218 74230 75454
rect 73910 75134 74230 75218
rect 73910 74898 73952 75134
rect 74188 74898 74230 75134
rect 73910 74866 74230 74898
rect 79840 75454 80160 75486
rect 79840 75218 79882 75454
rect 80118 75218 80160 75454
rect 79840 75134 80160 75218
rect 79840 74898 79882 75134
rect 80118 74898 80160 75134
rect 79840 74866 80160 74898
rect 85771 75454 86091 75486
rect 85771 75218 85813 75454
rect 86049 75218 86091 75454
rect 85771 75134 86091 75218
rect 85771 74898 85813 75134
rect 86049 74898 86091 75134
rect 85771 74866 86091 74898
rect 100910 75454 101230 75486
rect 100910 75218 100952 75454
rect 101188 75218 101230 75454
rect 100910 75134 101230 75218
rect 100910 74898 100952 75134
rect 101188 74898 101230 75134
rect 100910 74866 101230 74898
rect 106840 75454 107160 75486
rect 106840 75218 106882 75454
rect 107118 75218 107160 75454
rect 106840 75134 107160 75218
rect 106840 74898 106882 75134
rect 107118 74898 107160 75134
rect 106840 74866 107160 74898
rect 112771 75454 113091 75486
rect 112771 75218 112813 75454
rect 113049 75218 113091 75454
rect 112771 75134 113091 75218
rect 112771 74898 112813 75134
rect 113049 74898 113091 75134
rect 112771 74866 113091 74898
rect 127910 75454 128230 75486
rect 127910 75218 127952 75454
rect 128188 75218 128230 75454
rect 127910 75134 128230 75218
rect 127910 74898 127952 75134
rect 128188 74898 128230 75134
rect 127910 74866 128230 74898
rect 133840 75454 134160 75486
rect 133840 75218 133882 75454
rect 134118 75218 134160 75454
rect 133840 75134 134160 75218
rect 133840 74898 133882 75134
rect 134118 74898 134160 75134
rect 133840 74866 134160 74898
rect 139771 75454 140091 75486
rect 139771 75218 139813 75454
rect 140049 75218 140091 75454
rect 139771 75134 140091 75218
rect 139771 74898 139813 75134
rect 140049 74898 140091 75134
rect 139771 74866 140091 74898
rect 154910 75454 155230 75486
rect 154910 75218 154952 75454
rect 155188 75218 155230 75454
rect 154910 75134 155230 75218
rect 154910 74898 154952 75134
rect 155188 74898 155230 75134
rect 154910 74866 155230 74898
rect 160840 75454 161160 75486
rect 160840 75218 160882 75454
rect 161118 75218 161160 75454
rect 160840 75134 161160 75218
rect 160840 74898 160882 75134
rect 161118 74898 161160 75134
rect 160840 74866 161160 74898
rect 166771 75454 167091 75486
rect 166771 75218 166813 75454
rect 167049 75218 167091 75454
rect 166771 75134 167091 75218
rect 166771 74898 166813 75134
rect 167049 74898 167091 75134
rect 166771 74866 167091 74898
rect 181910 75454 182230 75486
rect 181910 75218 181952 75454
rect 182188 75218 182230 75454
rect 181910 75134 182230 75218
rect 181910 74898 181952 75134
rect 182188 74898 182230 75134
rect 181910 74866 182230 74898
rect 187840 75454 188160 75486
rect 187840 75218 187882 75454
rect 188118 75218 188160 75454
rect 187840 75134 188160 75218
rect 187840 74898 187882 75134
rect 188118 74898 188160 75134
rect 187840 74866 188160 74898
rect 193771 75454 194091 75486
rect 193771 75218 193813 75454
rect 194049 75218 194091 75454
rect 193771 75134 194091 75218
rect 193771 74898 193813 75134
rect 194049 74898 194091 75134
rect 193771 74866 194091 74898
rect 208910 75454 209230 75486
rect 208910 75218 208952 75454
rect 209188 75218 209230 75454
rect 208910 75134 209230 75218
rect 208910 74898 208952 75134
rect 209188 74898 209230 75134
rect 208910 74866 209230 74898
rect 214840 75454 215160 75486
rect 214840 75218 214882 75454
rect 215118 75218 215160 75454
rect 214840 75134 215160 75218
rect 214840 74898 214882 75134
rect 215118 74898 215160 75134
rect 214840 74866 215160 74898
rect 220771 75454 221091 75486
rect 220771 75218 220813 75454
rect 221049 75218 221091 75454
rect 220771 75134 221091 75218
rect 220771 74898 220813 75134
rect 221049 74898 221091 75134
rect 220771 74866 221091 74898
rect 235910 75454 236230 75486
rect 235910 75218 235952 75454
rect 236188 75218 236230 75454
rect 235910 75134 236230 75218
rect 235910 74898 235952 75134
rect 236188 74898 236230 75134
rect 235910 74866 236230 74898
rect 241840 75454 242160 75486
rect 241840 75218 241882 75454
rect 242118 75218 242160 75454
rect 241840 75134 242160 75218
rect 241840 74898 241882 75134
rect 242118 74898 242160 75134
rect 241840 74866 242160 74898
rect 247771 75454 248091 75486
rect 247771 75218 247813 75454
rect 248049 75218 248091 75454
rect 247771 75134 248091 75218
rect 247771 74898 247813 75134
rect 248049 74898 248091 75134
rect 247771 74866 248091 74898
rect 262910 75454 263230 75486
rect 262910 75218 262952 75454
rect 263188 75218 263230 75454
rect 262910 75134 263230 75218
rect 262910 74898 262952 75134
rect 263188 74898 263230 75134
rect 262910 74866 263230 74898
rect 268840 75454 269160 75486
rect 268840 75218 268882 75454
rect 269118 75218 269160 75454
rect 268840 75134 269160 75218
rect 268840 74898 268882 75134
rect 269118 74898 269160 75134
rect 268840 74866 269160 74898
rect 274771 75454 275091 75486
rect 274771 75218 274813 75454
rect 275049 75218 275091 75454
rect 274771 75134 275091 75218
rect 274771 74898 274813 75134
rect 275049 74898 275091 75134
rect 274771 74866 275091 74898
rect 289910 75454 290230 75486
rect 289910 75218 289952 75454
rect 290188 75218 290230 75454
rect 289910 75134 290230 75218
rect 289910 74898 289952 75134
rect 290188 74898 290230 75134
rect 289910 74866 290230 74898
rect 295840 75454 296160 75486
rect 295840 75218 295882 75454
rect 296118 75218 296160 75454
rect 295840 75134 296160 75218
rect 295840 74898 295882 75134
rect 296118 74898 296160 75134
rect 295840 74866 296160 74898
rect 301771 75454 302091 75486
rect 301771 75218 301813 75454
rect 302049 75218 302091 75454
rect 301771 75134 302091 75218
rect 301771 74898 301813 75134
rect 302049 74898 302091 75134
rect 301771 74866 302091 74898
rect 316910 75454 317230 75486
rect 316910 75218 316952 75454
rect 317188 75218 317230 75454
rect 316910 75134 317230 75218
rect 316910 74898 316952 75134
rect 317188 74898 317230 75134
rect 316910 74866 317230 74898
rect 322840 75454 323160 75486
rect 322840 75218 322882 75454
rect 323118 75218 323160 75454
rect 322840 75134 323160 75218
rect 322840 74898 322882 75134
rect 323118 74898 323160 75134
rect 322840 74866 323160 74898
rect 328771 75454 329091 75486
rect 328771 75218 328813 75454
rect 329049 75218 329091 75454
rect 328771 75134 329091 75218
rect 328771 74898 328813 75134
rect 329049 74898 329091 75134
rect 328771 74866 329091 74898
rect 343910 75454 344230 75486
rect 343910 75218 343952 75454
rect 344188 75218 344230 75454
rect 343910 75134 344230 75218
rect 343910 74898 343952 75134
rect 344188 74898 344230 75134
rect 343910 74866 344230 74898
rect 349840 75454 350160 75486
rect 349840 75218 349882 75454
rect 350118 75218 350160 75454
rect 349840 75134 350160 75218
rect 349840 74898 349882 75134
rect 350118 74898 350160 75134
rect 349840 74866 350160 74898
rect 355771 75454 356091 75486
rect 355771 75218 355813 75454
rect 356049 75218 356091 75454
rect 355771 75134 356091 75218
rect 355771 74898 355813 75134
rect 356049 74898 356091 75134
rect 355771 74866 356091 74898
rect 370910 75454 371230 75486
rect 370910 75218 370952 75454
rect 371188 75218 371230 75454
rect 370910 75134 371230 75218
rect 370910 74898 370952 75134
rect 371188 74898 371230 75134
rect 370910 74866 371230 74898
rect 376840 75454 377160 75486
rect 376840 75218 376882 75454
rect 377118 75218 377160 75454
rect 376840 75134 377160 75218
rect 376840 74898 376882 75134
rect 377118 74898 377160 75134
rect 376840 74866 377160 74898
rect 382771 75454 383091 75486
rect 382771 75218 382813 75454
rect 383049 75218 383091 75454
rect 382771 75134 383091 75218
rect 382771 74898 382813 75134
rect 383049 74898 383091 75134
rect 382771 74866 383091 74898
rect 397910 75454 398230 75486
rect 397910 75218 397952 75454
rect 398188 75218 398230 75454
rect 397910 75134 398230 75218
rect 397910 74898 397952 75134
rect 398188 74898 398230 75134
rect 397910 74866 398230 74898
rect 403840 75454 404160 75486
rect 403840 75218 403882 75454
rect 404118 75218 404160 75454
rect 403840 75134 404160 75218
rect 403840 74898 403882 75134
rect 404118 74898 404160 75134
rect 403840 74866 404160 74898
rect 409771 75454 410091 75486
rect 409771 75218 409813 75454
rect 410049 75218 410091 75454
rect 409771 75134 410091 75218
rect 409771 74898 409813 75134
rect 410049 74898 410091 75134
rect 409771 74866 410091 74898
rect 424910 75454 425230 75486
rect 424910 75218 424952 75454
rect 425188 75218 425230 75454
rect 424910 75134 425230 75218
rect 424910 74898 424952 75134
rect 425188 74898 425230 75134
rect 424910 74866 425230 74898
rect 430840 75454 431160 75486
rect 430840 75218 430882 75454
rect 431118 75218 431160 75454
rect 430840 75134 431160 75218
rect 430840 74898 430882 75134
rect 431118 74898 431160 75134
rect 430840 74866 431160 74898
rect 436771 75454 437091 75486
rect 436771 75218 436813 75454
rect 437049 75218 437091 75454
rect 436771 75134 437091 75218
rect 436771 74898 436813 75134
rect 437049 74898 437091 75134
rect 436771 74866 437091 74898
rect 451910 75454 452230 75486
rect 451910 75218 451952 75454
rect 452188 75218 452230 75454
rect 451910 75134 452230 75218
rect 451910 74898 451952 75134
rect 452188 74898 452230 75134
rect 451910 74866 452230 74898
rect 457840 75454 458160 75486
rect 457840 75218 457882 75454
rect 458118 75218 458160 75454
rect 457840 75134 458160 75218
rect 457840 74898 457882 75134
rect 458118 74898 458160 75134
rect 457840 74866 458160 74898
rect 463771 75454 464091 75486
rect 463771 75218 463813 75454
rect 464049 75218 464091 75454
rect 463771 75134 464091 75218
rect 463771 74898 463813 75134
rect 464049 74898 464091 75134
rect 463771 74866 464091 74898
rect 478910 75454 479230 75486
rect 478910 75218 478952 75454
rect 479188 75218 479230 75454
rect 478910 75134 479230 75218
rect 478910 74898 478952 75134
rect 479188 74898 479230 75134
rect 478910 74866 479230 74898
rect 484840 75454 485160 75486
rect 484840 75218 484882 75454
rect 485118 75218 485160 75454
rect 484840 75134 485160 75218
rect 484840 74898 484882 75134
rect 485118 74898 485160 75134
rect 484840 74866 485160 74898
rect 490771 75454 491091 75486
rect 490771 75218 490813 75454
rect 491049 75218 491091 75454
rect 490771 75134 491091 75218
rect 490771 74898 490813 75134
rect 491049 74898 491091 75134
rect 490771 74866 491091 74898
rect 505910 75454 506230 75486
rect 505910 75218 505952 75454
rect 506188 75218 506230 75454
rect 505910 75134 506230 75218
rect 505910 74898 505952 75134
rect 506188 74898 506230 75134
rect 505910 74866 506230 74898
rect 511840 75454 512160 75486
rect 511840 75218 511882 75454
rect 512118 75218 512160 75454
rect 511840 75134 512160 75218
rect 511840 74898 511882 75134
rect 512118 74898 512160 75134
rect 511840 74866 512160 74898
rect 517771 75454 518091 75486
rect 517771 75218 517813 75454
rect 518049 75218 518091 75454
rect 517771 75134 518091 75218
rect 517771 74898 517813 75134
rect 518049 74898 518091 75134
rect 517771 74866 518091 74898
rect 532910 75454 533230 75486
rect 532910 75218 532952 75454
rect 533188 75218 533230 75454
rect 532910 75134 533230 75218
rect 532910 74898 532952 75134
rect 533188 74898 533230 75134
rect 532910 74866 533230 74898
rect 538840 75454 539160 75486
rect 538840 75218 538882 75454
rect 539118 75218 539160 75454
rect 538840 75134 539160 75218
rect 538840 74898 538882 75134
rect 539118 74898 539160 75134
rect 538840 74866 539160 74898
rect 544771 75454 545091 75486
rect 544771 75218 544813 75454
rect 545049 75218 545091 75454
rect 544771 75134 545091 75218
rect 544771 74898 544813 75134
rect 545049 74898 545091 75134
rect 544771 74866 545091 74898
rect 559794 75454 560414 92898
rect 559794 75218 559826 75454
rect 560062 75218 560146 75454
rect 560382 75218 560414 75454
rect 559794 75134 560414 75218
rect 559794 74898 559826 75134
rect 560062 74898 560146 75134
rect 560382 74898 560414 75134
rect 10794 66218 10826 66454
rect 11062 66218 11146 66454
rect 11382 66218 11414 66454
rect 10794 66134 11414 66218
rect 10794 65898 10826 66134
rect 11062 65898 11146 66134
rect 11382 65898 11414 66134
rect 10794 48454 11414 65898
rect 19794 67394 20414 68000
rect 19794 67158 19826 67394
rect 20062 67158 20146 67394
rect 20382 67158 20414 67394
rect 19794 67074 20414 67158
rect 19794 66838 19826 67074
rect 20062 66838 20146 67074
rect 20382 66838 20414 67074
rect 19794 65000 20414 66838
rect 28794 66454 29414 68000
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 65000 29414 65898
rect 37794 67394 38414 68000
rect 37794 67158 37826 67394
rect 38062 67158 38146 67394
rect 38382 67158 38414 67394
rect 37794 67074 38414 67158
rect 37794 66838 37826 67074
rect 38062 66838 38146 67074
rect 38382 66838 38414 67074
rect 37794 65000 38414 66838
rect 46794 66454 47414 68000
rect 46794 66218 46826 66454
rect 47062 66218 47146 66454
rect 47382 66218 47414 66454
rect 46794 66134 47414 66218
rect 46794 65898 46826 66134
rect 47062 65898 47146 66134
rect 47382 65898 47414 66134
rect 46794 65000 47414 65898
rect 55794 67394 56414 68000
rect 55794 67158 55826 67394
rect 56062 67158 56146 67394
rect 56382 67158 56414 67394
rect 55794 67074 56414 67158
rect 55794 66838 55826 67074
rect 56062 66838 56146 67074
rect 56382 66838 56414 67074
rect 55794 65000 56414 66838
rect 64794 66454 65414 68000
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 65000 65414 65898
rect 73794 67394 74414 68000
rect 73794 67158 73826 67394
rect 74062 67158 74146 67394
rect 74382 67158 74414 67394
rect 73794 67074 74414 67158
rect 73794 66838 73826 67074
rect 74062 66838 74146 67074
rect 74382 66838 74414 67074
rect 73794 65000 74414 66838
rect 82794 66454 83414 68000
rect 82794 66218 82826 66454
rect 83062 66218 83146 66454
rect 83382 66218 83414 66454
rect 82794 66134 83414 66218
rect 82794 65898 82826 66134
rect 83062 65898 83146 66134
rect 83382 65898 83414 66134
rect 82794 65000 83414 65898
rect 91794 67394 92414 68000
rect 91794 67158 91826 67394
rect 92062 67158 92146 67394
rect 92382 67158 92414 67394
rect 91794 67074 92414 67158
rect 91794 66838 91826 67074
rect 92062 66838 92146 67074
rect 92382 66838 92414 67074
rect 91794 65000 92414 66838
rect 100794 66454 101414 68000
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 65000 101414 65898
rect 109794 67394 110414 68000
rect 109794 67158 109826 67394
rect 110062 67158 110146 67394
rect 110382 67158 110414 67394
rect 109794 67074 110414 67158
rect 109794 66838 109826 67074
rect 110062 66838 110146 67074
rect 110382 66838 110414 67074
rect 109794 65000 110414 66838
rect 118794 66454 119414 68000
rect 118794 66218 118826 66454
rect 119062 66218 119146 66454
rect 119382 66218 119414 66454
rect 118794 66134 119414 66218
rect 118794 65898 118826 66134
rect 119062 65898 119146 66134
rect 119382 65898 119414 66134
rect 118794 65000 119414 65898
rect 127794 67394 128414 68000
rect 127794 67158 127826 67394
rect 128062 67158 128146 67394
rect 128382 67158 128414 67394
rect 127794 67074 128414 67158
rect 127794 66838 127826 67074
rect 128062 66838 128146 67074
rect 128382 66838 128414 67074
rect 127794 65000 128414 66838
rect 136794 66454 137414 68000
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 65000 137414 65898
rect 145794 67394 146414 68000
rect 145794 67158 145826 67394
rect 146062 67158 146146 67394
rect 146382 67158 146414 67394
rect 145794 67074 146414 67158
rect 145794 66838 145826 67074
rect 146062 66838 146146 67074
rect 146382 66838 146414 67074
rect 145794 65000 146414 66838
rect 154794 66454 155414 68000
rect 154794 66218 154826 66454
rect 155062 66218 155146 66454
rect 155382 66218 155414 66454
rect 154794 66134 155414 66218
rect 154794 65898 154826 66134
rect 155062 65898 155146 66134
rect 155382 65898 155414 66134
rect 154794 65000 155414 65898
rect 163794 67394 164414 68000
rect 163794 67158 163826 67394
rect 164062 67158 164146 67394
rect 164382 67158 164414 67394
rect 163794 67074 164414 67158
rect 163794 66838 163826 67074
rect 164062 66838 164146 67074
rect 164382 66838 164414 67074
rect 163794 65000 164414 66838
rect 172794 66454 173414 68000
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172794 65000 173414 65898
rect 181794 67394 182414 68000
rect 181794 67158 181826 67394
rect 182062 67158 182146 67394
rect 182382 67158 182414 67394
rect 181794 67074 182414 67158
rect 181794 66838 181826 67074
rect 182062 66838 182146 67074
rect 182382 66838 182414 67074
rect 181794 65000 182414 66838
rect 190794 66454 191414 68000
rect 190794 66218 190826 66454
rect 191062 66218 191146 66454
rect 191382 66218 191414 66454
rect 190794 66134 191414 66218
rect 190794 65898 190826 66134
rect 191062 65898 191146 66134
rect 191382 65898 191414 66134
rect 190794 65000 191414 65898
rect 199794 67394 200414 68000
rect 199794 67158 199826 67394
rect 200062 67158 200146 67394
rect 200382 67158 200414 67394
rect 199794 67074 200414 67158
rect 199794 66838 199826 67074
rect 200062 66838 200146 67074
rect 200382 66838 200414 67074
rect 199794 65000 200414 66838
rect 208794 66454 209414 68000
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 65000 209414 65898
rect 217794 67394 218414 68000
rect 217794 67158 217826 67394
rect 218062 67158 218146 67394
rect 218382 67158 218414 67394
rect 217794 67074 218414 67158
rect 217794 66838 217826 67074
rect 218062 66838 218146 67074
rect 218382 66838 218414 67074
rect 217794 65000 218414 66838
rect 226794 66454 227414 68000
rect 226794 66218 226826 66454
rect 227062 66218 227146 66454
rect 227382 66218 227414 66454
rect 226794 66134 227414 66218
rect 226794 65898 226826 66134
rect 227062 65898 227146 66134
rect 227382 65898 227414 66134
rect 226794 65000 227414 65898
rect 235794 67394 236414 68000
rect 235794 67158 235826 67394
rect 236062 67158 236146 67394
rect 236382 67158 236414 67394
rect 235794 67074 236414 67158
rect 235794 66838 235826 67074
rect 236062 66838 236146 67074
rect 236382 66838 236414 67074
rect 235794 65000 236414 66838
rect 244794 66454 245414 68000
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 65000 245414 65898
rect 253794 67394 254414 68000
rect 253794 67158 253826 67394
rect 254062 67158 254146 67394
rect 254382 67158 254414 67394
rect 253794 67074 254414 67158
rect 253794 66838 253826 67074
rect 254062 66838 254146 67074
rect 254382 66838 254414 67074
rect 253794 65000 254414 66838
rect 262794 66454 263414 68000
rect 262794 66218 262826 66454
rect 263062 66218 263146 66454
rect 263382 66218 263414 66454
rect 262794 66134 263414 66218
rect 262794 65898 262826 66134
rect 263062 65898 263146 66134
rect 263382 65898 263414 66134
rect 262794 65000 263414 65898
rect 271794 67394 272414 68000
rect 271794 67158 271826 67394
rect 272062 67158 272146 67394
rect 272382 67158 272414 67394
rect 271794 67074 272414 67158
rect 271794 66838 271826 67074
rect 272062 66838 272146 67074
rect 272382 66838 272414 67074
rect 271794 65000 272414 66838
rect 280794 66454 281414 68000
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 65000 281414 65898
rect 289794 67394 290414 68000
rect 289794 67158 289826 67394
rect 290062 67158 290146 67394
rect 290382 67158 290414 67394
rect 289794 67074 290414 67158
rect 289794 66838 289826 67074
rect 290062 66838 290146 67074
rect 290382 66838 290414 67074
rect 289794 65000 290414 66838
rect 298794 66454 299414 68000
rect 298794 66218 298826 66454
rect 299062 66218 299146 66454
rect 299382 66218 299414 66454
rect 298794 66134 299414 66218
rect 298794 65898 298826 66134
rect 299062 65898 299146 66134
rect 299382 65898 299414 66134
rect 298794 65000 299414 65898
rect 307794 67394 308414 68000
rect 307794 67158 307826 67394
rect 308062 67158 308146 67394
rect 308382 67158 308414 67394
rect 307794 67074 308414 67158
rect 307794 66838 307826 67074
rect 308062 66838 308146 67074
rect 308382 66838 308414 67074
rect 307794 65000 308414 66838
rect 316794 66454 317414 68000
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 65000 317414 65898
rect 325794 67394 326414 68000
rect 325794 67158 325826 67394
rect 326062 67158 326146 67394
rect 326382 67158 326414 67394
rect 325794 67074 326414 67158
rect 325794 66838 325826 67074
rect 326062 66838 326146 67074
rect 326382 66838 326414 67074
rect 325794 65000 326414 66838
rect 334794 66454 335414 68000
rect 334794 66218 334826 66454
rect 335062 66218 335146 66454
rect 335382 66218 335414 66454
rect 334794 66134 335414 66218
rect 334794 65898 334826 66134
rect 335062 65898 335146 66134
rect 335382 65898 335414 66134
rect 334794 65000 335414 65898
rect 343794 67394 344414 68000
rect 343794 67158 343826 67394
rect 344062 67158 344146 67394
rect 344382 67158 344414 67394
rect 343794 67074 344414 67158
rect 343794 66838 343826 67074
rect 344062 66838 344146 67074
rect 344382 66838 344414 67074
rect 343794 65000 344414 66838
rect 352794 66454 353414 68000
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 65000 353414 65898
rect 361794 67394 362414 68000
rect 361794 67158 361826 67394
rect 362062 67158 362146 67394
rect 362382 67158 362414 67394
rect 361794 67074 362414 67158
rect 361794 66838 361826 67074
rect 362062 66838 362146 67074
rect 362382 66838 362414 67074
rect 361794 65000 362414 66838
rect 370794 66454 371414 68000
rect 370794 66218 370826 66454
rect 371062 66218 371146 66454
rect 371382 66218 371414 66454
rect 370794 66134 371414 66218
rect 370794 65898 370826 66134
rect 371062 65898 371146 66134
rect 371382 65898 371414 66134
rect 370794 65000 371414 65898
rect 379794 67394 380414 68000
rect 379794 67158 379826 67394
rect 380062 67158 380146 67394
rect 380382 67158 380414 67394
rect 379794 67074 380414 67158
rect 379794 66838 379826 67074
rect 380062 66838 380146 67074
rect 380382 66838 380414 67074
rect 379794 65000 380414 66838
rect 388794 66454 389414 68000
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 65000 389414 65898
rect 397794 67394 398414 68000
rect 397794 67158 397826 67394
rect 398062 67158 398146 67394
rect 398382 67158 398414 67394
rect 397794 67074 398414 67158
rect 397794 66838 397826 67074
rect 398062 66838 398146 67074
rect 398382 66838 398414 67074
rect 397794 65000 398414 66838
rect 406794 66454 407414 68000
rect 406794 66218 406826 66454
rect 407062 66218 407146 66454
rect 407382 66218 407414 66454
rect 406794 66134 407414 66218
rect 406794 65898 406826 66134
rect 407062 65898 407146 66134
rect 407382 65898 407414 66134
rect 406794 65000 407414 65898
rect 415794 67394 416414 68000
rect 415794 67158 415826 67394
rect 416062 67158 416146 67394
rect 416382 67158 416414 67394
rect 415794 67074 416414 67158
rect 415794 66838 415826 67074
rect 416062 66838 416146 67074
rect 416382 66838 416414 67074
rect 415794 65000 416414 66838
rect 424794 66454 425414 68000
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 65000 425414 65898
rect 433794 67394 434414 68000
rect 433794 67158 433826 67394
rect 434062 67158 434146 67394
rect 434382 67158 434414 67394
rect 433794 67074 434414 67158
rect 433794 66838 433826 67074
rect 434062 66838 434146 67074
rect 434382 66838 434414 67074
rect 433794 65000 434414 66838
rect 442794 66454 443414 68000
rect 442794 66218 442826 66454
rect 443062 66218 443146 66454
rect 443382 66218 443414 66454
rect 442794 66134 443414 66218
rect 442794 65898 442826 66134
rect 443062 65898 443146 66134
rect 443382 65898 443414 66134
rect 442794 65000 443414 65898
rect 451794 67394 452414 68000
rect 451794 67158 451826 67394
rect 452062 67158 452146 67394
rect 452382 67158 452414 67394
rect 451794 67074 452414 67158
rect 451794 66838 451826 67074
rect 452062 66838 452146 67074
rect 452382 66838 452414 67074
rect 451794 65000 452414 66838
rect 460794 66454 461414 68000
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 65000 461414 65898
rect 469794 67394 470414 68000
rect 469794 67158 469826 67394
rect 470062 67158 470146 67394
rect 470382 67158 470414 67394
rect 469794 67074 470414 67158
rect 469794 66838 469826 67074
rect 470062 66838 470146 67074
rect 470382 66838 470414 67074
rect 469794 65000 470414 66838
rect 478794 66454 479414 68000
rect 478794 66218 478826 66454
rect 479062 66218 479146 66454
rect 479382 66218 479414 66454
rect 478794 66134 479414 66218
rect 478794 65898 478826 66134
rect 479062 65898 479146 66134
rect 479382 65898 479414 66134
rect 478794 65000 479414 65898
rect 487794 67394 488414 68000
rect 487794 67158 487826 67394
rect 488062 67158 488146 67394
rect 488382 67158 488414 67394
rect 487794 67074 488414 67158
rect 487794 66838 487826 67074
rect 488062 66838 488146 67074
rect 488382 66838 488414 67074
rect 487794 65000 488414 66838
rect 496794 66454 497414 68000
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 65000 497414 65898
rect 505794 67394 506414 68000
rect 505794 67158 505826 67394
rect 506062 67158 506146 67394
rect 506382 67158 506414 67394
rect 505794 67074 506414 67158
rect 505794 66838 505826 67074
rect 506062 66838 506146 67074
rect 506382 66838 506414 67074
rect 505794 65000 506414 66838
rect 514794 66454 515414 68000
rect 514794 66218 514826 66454
rect 515062 66218 515146 66454
rect 515382 66218 515414 66454
rect 514794 66134 515414 66218
rect 514794 65898 514826 66134
rect 515062 65898 515146 66134
rect 515382 65898 515414 66134
rect 514794 65000 515414 65898
rect 523794 67394 524414 68000
rect 523794 67158 523826 67394
rect 524062 67158 524146 67394
rect 524382 67158 524414 67394
rect 523794 67074 524414 67158
rect 523794 66838 523826 67074
rect 524062 66838 524146 67074
rect 524382 66838 524414 67074
rect 523794 65000 524414 66838
rect 532794 66454 533414 68000
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 65000 533414 65898
rect 541794 67394 542414 68000
rect 541794 67158 541826 67394
rect 542062 67158 542146 67394
rect 542382 67158 542414 67394
rect 541794 67074 542414 67158
rect 541794 66838 541826 67074
rect 542062 66838 542146 67074
rect 542382 66838 542414 67074
rect 541794 65000 542414 66838
rect 550794 66454 551414 68000
rect 550794 66218 550826 66454
rect 551062 66218 551146 66454
rect 551382 66218 551414 66454
rect 550794 66134 551414 66218
rect 550794 65898 550826 66134
rect 551062 65898 551146 66134
rect 551382 65898 551414 66134
rect 550794 65000 551414 65898
rect 19910 57454 20230 57486
rect 19910 57218 19952 57454
rect 20188 57218 20230 57454
rect 19910 57134 20230 57218
rect 19910 56898 19952 57134
rect 20188 56898 20230 57134
rect 19910 56866 20230 56898
rect 25840 57454 26160 57486
rect 25840 57218 25882 57454
rect 26118 57218 26160 57454
rect 25840 57134 26160 57218
rect 25840 56898 25882 57134
rect 26118 56898 26160 57134
rect 25840 56866 26160 56898
rect 31771 57454 32091 57486
rect 31771 57218 31813 57454
rect 32049 57218 32091 57454
rect 31771 57134 32091 57218
rect 31771 56898 31813 57134
rect 32049 56898 32091 57134
rect 31771 56866 32091 56898
rect 46910 57454 47230 57486
rect 46910 57218 46952 57454
rect 47188 57218 47230 57454
rect 46910 57134 47230 57218
rect 46910 56898 46952 57134
rect 47188 56898 47230 57134
rect 46910 56866 47230 56898
rect 52840 57454 53160 57486
rect 52840 57218 52882 57454
rect 53118 57218 53160 57454
rect 52840 57134 53160 57218
rect 52840 56898 52882 57134
rect 53118 56898 53160 57134
rect 52840 56866 53160 56898
rect 58771 57454 59091 57486
rect 58771 57218 58813 57454
rect 59049 57218 59091 57454
rect 58771 57134 59091 57218
rect 58771 56898 58813 57134
rect 59049 56898 59091 57134
rect 58771 56866 59091 56898
rect 73910 57454 74230 57486
rect 73910 57218 73952 57454
rect 74188 57218 74230 57454
rect 73910 57134 74230 57218
rect 73910 56898 73952 57134
rect 74188 56898 74230 57134
rect 73910 56866 74230 56898
rect 79840 57454 80160 57486
rect 79840 57218 79882 57454
rect 80118 57218 80160 57454
rect 79840 57134 80160 57218
rect 79840 56898 79882 57134
rect 80118 56898 80160 57134
rect 79840 56866 80160 56898
rect 85771 57454 86091 57486
rect 85771 57218 85813 57454
rect 86049 57218 86091 57454
rect 85771 57134 86091 57218
rect 85771 56898 85813 57134
rect 86049 56898 86091 57134
rect 85771 56866 86091 56898
rect 100910 57454 101230 57486
rect 100910 57218 100952 57454
rect 101188 57218 101230 57454
rect 100910 57134 101230 57218
rect 100910 56898 100952 57134
rect 101188 56898 101230 57134
rect 100910 56866 101230 56898
rect 106840 57454 107160 57486
rect 106840 57218 106882 57454
rect 107118 57218 107160 57454
rect 106840 57134 107160 57218
rect 106840 56898 106882 57134
rect 107118 56898 107160 57134
rect 106840 56866 107160 56898
rect 112771 57454 113091 57486
rect 112771 57218 112813 57454
rect 113049 57218 113091 57454
rect 112771 57134 113091 57218
rect 112771 56898 112813 57134
rect 113049 56898 113091 57134
rect 112771 56866 113091 56898
rect 127910 57454 128230 57486
rect 127910 57218 127952 57454
rect 128188 57218 128230 57454
rect 127910 57134 128230 57218
rect 127910 56898 127952 57134
rect 128188 56898 128230 57134
rect 127910 56866 128230 56898
rect 133840 57454 134160 57486
rect 133840 57218 133882 57454
rect 134118 57218 134160 57454
rect 133840 57134 134160 57218
rect 133840 56898 133882 57134
rect 134118 56898 134160 57134
rect 133840 56866 134160 56898
rect 139771 57454 140091 57486
rect 139771 57218 139813 57454
rect 140049 57218 140091 57454
rect 139771 57134 140091 57218
rect 139771 56898 139813 57134
rect 140049 56898 140091 57134
rect 139771 56866 140091 56898
rect 154910 57454 155230 57486
rect 154910 57218 154952 57454
rect 155188 57218 155230 57454
rect 154910 57134 155230 57218
rect 154910 56898 154952 57134
rect 155188 56898 155230 57134
rect 154910 56866 155230 56898
rect 160840 57454 161160 57486
rect 160840 57218 160882 57454
rect 161118 57218 161160 57454
rect 160840 57134 161160 57218
rect 160840 56898 160882 57134
rect 161118 56898 161160 57134
rect 160840 56866 161160 56898
rect 166771 57454 167091 57486
rect 166771 57218 166813 57454
rect 167049 57218 167091 57454
rect 166771 57134 167091 57218
rect 166771 56898 166813 57134
rect 167049 56898 167091 57134
rect 166771 56866 167091 56898
rect 181910 57454 182230 57486
rect 181910 57218 181952 57454
rect 182188 57218 182230 57454
rect 181910 57134 182230 57218
rect 181910 56898 181952 57134
rect 182188 56898 182230 57134
rect 181910 56866 182230 56898
rect 187840 57454 188160 57486
rect 187840 57218 187882 57454
rect 188118 57218 188160 57454
rect 187840 57134 188160 57218
rect 187840 56898 187882 57134
rect 188118 56898 188160 57134
rect 187840 56866 188160 56898
rect 193771 57454 194091 57486
rect 193771 57218 193813 57454
rect 194049 57218 194091 57454
rect 193771 57134 194091 57218
rect 193771 56898 193813 57134
rect 194049 56898 194091 57134
rect 193771 56866 194091 56898
rect 208910 57454 209230 57486
rect 208910 57218 208952 57454
rect 209188 57218 209230 57454
rect 208910 57134 209230 57218
rect 208910 56898 208952 57134
rect 209188 56898 209230 57134
rect 208910 56866 209230 56898
rect 214840 57454 215160 57486
rect 214840 57218 214882 57454
rect 215118 57218 215160 57454
rect 214840 57134 215160 57218
rect 214840 56898 214882 57134
rect 215118 56898 215160 57134
rect 214840 56866 215160 56898
rect 220771 57454 221091 57486
rect 220771 57218 220813 57454
rect 221049 57218 221091 57454
rect 220771 57134 221091 57218
rect 220771 56898 220813 57134
rect 221049 56898 221091 57134
rect 220771 56866 221091 56898
rect 235910 57454 236230 57486
rect 235910 57218 235952 57454
rect 236188 57218 236230 57454
rect 235910 57134 236230 57218
rect 235910 56898 235952 57134
rect 236188 56898 236230 57134
rect 235910 56866 236230 56898
rect 241840 57454 242160 57486
rect 241840 57218 241882 57454
rect 242118 57218 242160 57454
rect 241840 57134 242160 57218
rect 241840 56898 241882 57134
rect 242118 56898 242160 57134
rect 241840 56866 242160 56898
rect 247771 57454 248091 57486
rect 247771 57218 247813 57454
rect 248049 57218 248091 57454
rect 247771 57134 248091 57218
rect 247771 56898 247813 57134
rect 248049 56898 248091 57134
rect 247771 56866 248091 56898
rect 262910 57454 263230 57486
rect 262910 57218 262952 57454
rect 263188 57218 263230 57454
rect 262910 57134 263230 57218
rect 262910 56898 262952 57134
rect 263188 56898 263230 57134
rect 262910 56866 263230 56898
rect 268840 57454 269160 57486
rect 268840 57218 268882 57454
rect 269118 57218 269160 57454
rect 268840 57134 269160 57218
rect 268840 56898 268882 57134
rect 269118 56898 269160 57134
rect 268840 56866 269160 56898
rect 274771 57454 275091 57486
rect 274771 57218 274813 57454
rect 275049 57218 275091 57454
rect 274771 57134 275091 57218
rect 274771 56898 274813 57134
rect 275049 56898 275091 57134
rect 274771 56866 275091 56898
rect 289910 57454 290230 57486
rect 289910 57218 289952 57454
rect 290188 57218 290230 57454
rect 289910 57134 290230 57218
rect 289910 56898 289952 57134
rect 290188 56898 290230 57134
rect 289910 56866 290230 56898
rect 295840 57454 296160 57486
rect 295840 57218 295882 57454
rect 296118 57218 296160 57454
rect 295840 57134 296160 57218
rect 295840 56898 295882 57134
rect 296118 56898 296160 57134
rect 295840 56866 296160 56898
rect 301771 57454 302091 57486
rect 301771 57218 301813 57454
rect 302049 57218 302091 57454
rect 301771 57134 302091 57218
rect 301771 56898 301813 57134
rect 302049 56898 302091 57134
rect 301771 56866 302091 56898
rect 316910 57454 317230 57486
rect 316910 57218 316952 57454
rect 317188 57218 317230 57454
rect 316910 57134 317230 57218
rect 316910 56898 316952 57134
rect 317188 56898 317230 57134
rect 316910 56866 317230 56898
rect 322840 57454 323160 57486
rect 322840 57218 322882 57454
rect 323118 57218 323160 57454
rect 322840 57134 323160 57218
rect 322840 56898 322882 57134
rect 323118 56898 323160 57134
rect 322840 56866 323160 56898
rect 328771 57454 329091 57486
rect 328771 57218 328813 57454
rect 329049 57218 329091 57454
rect 328771 57134 329091 57218
rect 328771 56898 328813 57134
rect 329049 56898 329091 57134
rect 328771 56866 329091 56898
rect 343910 57454 344230 57486
rect 343910 57218 343952 57454
rect 344188 57218 344230 57454
rect 343910 57134 344230 57218
rect 343910 56898 343952 57134
rect 344188 56898 344230 57134
rect 343910 56866 344230 56898
rect 349840 57454 350160 57486
rect 349840 57218 349882 57454
rect 350118 57218 350160 57454
rect 349840 57134 350160 57218
rect 349840 56898 349882 57134
rect 350118 56898 350160 57134
rect 349840 56866 350160 56898
rect 355771 57454 356091 57486
rect 355771 57218 355813 57454
rect 356049 57218 356091 57454
rect 355771 57134 356091 57218
rect 355771 56898 355813 57134
rect 356049 56898 356091 57134
rect 355771 56866 356091 56898
rect 370910 57454 371230 57486
rect 370910 57218 370952 57454
rect 371188 57218 371230 57454
rect 370910 57134 371230 57218
rect 370910 56898 370952 57134
rect 371188 56898 371230 57134
rect 370910 56866 371230 56898
rect 376840 57454 377160 57486
rect 376840 57218 376882 57454
rect 377118 57218 377160 57454
rect 376840 57134 377160 57218
rect 376840 56898 376882 57134
rect 377118 56898 377160 57134
rect 376840 56866 377160 56898
rect 382771 57454 383091 57486
rect 382771 57218 382813 57454
rect 383049 57218 383091 57454
rect 382771 57134 383091 57218
rect 382771 56898 382813 57134
rect 383049 56898 383091 57134
rect 382771 56866 383091 56898
rect 397910 57454 398230 57486
rect 397910 57218 397952 57454
rect 398188 57218 398230 57454
rect 397910 57134 398230 57218
rect 397910 56898 397952 57134
rect 398188 56898 398230 57134
rect 397910 56866 398230 56898
rect 403840 57454 404160 57486
rect 403840 57218 403882 57454
rect 404118 57218 404160 57454
rect 403840 57134 404160 57218
rect 403840 56898 403882 57134
rect 404118 56898 404160 57134
rect 403840 56866 404160 56898
rect 409771 57454 410091 57486
rect 409771 57218 409813 57454
rect 410049 57218 410091 57454
rect 409771 57134 410091 57218
rect 409771 56898 409813 57134
rect 410049 56898 410091 57134
rect 409771 56866 410091 56898
rect 424910 57454 425230 57486
rect 424910 57218 424952 57454
rect 425188 57218 425230 57454
rect 424910 57134 425230 57218
rect 424910 56898 424952 57134
rect 425188 56898 425230 57134
rect 424910 56866 425230 56898
rect 430840 57454 431160 57486
rect 430840 57218 430882 57454
rect 431118 57218 431160 57454
rect 430840 57134 431160 57218
rect 430840 56898 430882 57134
rect 431118 56898 431160 57134
rect 430840 56866 431160 56898
rect 436771 57454 437091 57486
rect 436771 57218 436813 57454
rect 437049 57218 437091 57454
rect 436771 57134 437091 57218
rect 436771 56898 436813 57134
rect 437049 56898 437091 57134
rect 436771 56866 437091 56898
rect 451910 57454 452230 57486
rect 451910 57218 451952 57454
rect 452188 57218 452230 57454
rect 451910 57134 452230 57218
rect 451910 56898 451952 57134
rect 452188 56898 452230 57134
rect 451910 56866 452230 56898
rect 457840 57454 458160 57486
rect 457840 57218 457882 57454
rect 458118 57218 458160 57454
rect 457840 57134 458160 57218
rect 457840 56898 457882 57134
rect 458118 56898 458160 57134
rect 457840 56866 458160 56898
rect 463771 57454 464091 57486
rect 463771 57218 463813 57454
rect 464049 57218 464091 57454
rect 463771 57134 464091 57218
rect 463771 56898 463813 57134
rect 464049 56898 464091 57134
rect 463771 56866 464091 56898
rect 478910 57454 479230 57486
rect 478910 57218 478952 57454
rect 479188 57218 479230 57454
rect 478910 57134 479230 57218
rect 478910 56898 478952 57134
rect 479188 56898 479230 57134
rect 478910 56866 479230 56898
rect 484840 57454 485160 57486
rect 484840 57218 484882 57454
rect 485118 57218 485160 57454
rect 484840 57134 485160 57218
rect 484840 56898 484882 57134
rect 485118 56898 485160 57134
rect 484840 56866 485160 56898
rect 490771 57454 491091 57486
rect 490771 57218 490813 57454
rect 491049 57218 491091 57454
rect 490771 57134 491091 57218
rect 490771 56898 490813 57134
rect 491049 56898 491091 57134
rect 490771 56866 491091 56898
rect 505910 57454 506230 57486
rect 505910 57218 505952 57454
rect 506188 57218 506230 57454
rect 505910 57134 506230 57218
rect 505910 56898 505952 57134
rect 506188 56898 506230 57134
rect 505910 56866 506230 56898
rect 511840 57454 512160 57486
rect 511840 57218 511882 57454
rect 512118 57218 512160 57454
rect 511840 57134 512160 57218
rect 511840 56898 511882 57134
rect 512118 56898 512160 57134
rect 511840 56866 512160 56898
rect 517771 57454 518091 57486
rect 517771 57218 517813 57454
rect 518049 57218 518091 57454
rect 517771 57134 518091 57218
rect 517771 56898 517813 57134
rect 518049 56898 518091 57134
rect 517771 56866 518091 56898
rect 532910 57454 533230 57486
rect 532910 57218 532952 57454
rect 533188 57218 533230 57454
rect 532910 57134 533230 57218
rect 532910 56898 532952 57134
rect 533188 56898 533230 57134
rect 532910 56866 533230 56898
rect 538840 57454 539160 57486
rect 538840 57218 538882 57454
rect 539118 57218 539160 57454
rect 538840 57134 539160 57218
rect 538840 56898 538882 57134
rect 539118 56898 539160 57134
rect 538840 56866 539160 56898
rect 544771 57454 545091 57486
rect 544771 57218 544813 57454
rect 545049 57218 545091 57454
rect 544771 57134 545091 57218
rect 544771 56898 544813 57134
rect 545049 56898 545091 57134
rect 544771 56866 545091 56898
rect 559794 57454 560414 74898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 30454 11414 47898
rect 22874 48454 23194 48486
rect 22874 48218 22916 48454
rect 23152 48218 23194 48454
rect 22874 48134 23194 48218
rect 22874 47898 22916 48134
rect 23152 47898 23194 48134
rect 22874 47866 23194 47898
rect 28805 48454 29125 48486
rect 28805 48218 28847 48454
rect 29083 48218 29125 48454
rect 28805 48134 29125 48218
rect 28805 47898 28847 48134
rect 29083 47898 29125 48134
rect 28805 47866 29125 47898
rect 49874 48454 50194 48486
rect 49874 48218 49916 48454
rect 50152 48218 50194 48454
rect 49874 48134 50194 48218
rect 49874 47898 49916 48134
rect 50152 47898 50194 48134
rect 49874 47866 50194 47898
rect 55805 48454 56125 48486
rect 55805 48218 55847 48454
rect 56083 48218 56125 48454
rect 55805 48134 56125 48218
rect 55805 47898 55847 48134
rect 56083 47898 56125 48134
rect 55805 47866 56125 47898
rect 76874 48454 77194 48486
rect 76874 48218 76916 48454
rect 77152 48218 77194 48454
rect 76874 48134 77194 48218
rect 76874 47898 76916 48134
rect 77152 47898 77194 48134
rect 76874 47866 77194 47898
rect 82805 48454 83125 48486
rect 82805 48218 82847 48454
rect 83083 48218 83125 48454
rect 82805 48134 83125 48218
rect 82805 47898 82847 48134
rect 83083 47898 83125 48134
rect 82805 47866 83125 47898
rect 103874 48454 104194 48486
rect 103874 48218 103916 48454
rect 104152 48218 104194 48454
rect 103874 48134 104194 48218
rect 103874 47898 103916 48134
rect 104152 47898 104194 48134
rect 103874 47866 104194 47898
rect 109805 48454 110125 48486
rect 109805 48218 109847 48454
rect 110083 48218 110125 48454
rect 109805 48134 110125 48218
rect 109805 47898 109847 48134
rect 110083 47898 110125 48134
rect 109805 47866 110125 47898
rect 130874 48454 131194 48486
rect 130874 48218 130916 48454
rect 131152 48218 131194 48454
rect 130874 48134 131194 48218
rect 130874 47898 130916 48134
rect 131152 47898 131194 48134
rect 130874 47866 131194 47898
rect 136805 48454 137125 48486
rect 136805 48218 136847 48454
rect 137083 48218 137125 48454
rect 136805 48134 137125 48218
rect 136805 47898 136847 48134
rect 137083 47898 137125 48134
rect 136805 47866 137125 47898
rect 157874 48454 158194 48486
rect 157874 48218 157916 48454
rect 158152 48218 158194 48454
rect 157874 48134 158194 48218
rect 157874 47898 157916 48134
rect 158152 47898 158194 48134
rect 157874 47866 158194 47898
rect 163805 48454 164125 48486
rect 163805 48218 163847 48454
rect 164083 48218 164125 48454
rect 163805 48134 164125 48218
rect 163805 47898 163847 48134
rect 164083 47898 164125 48134
rect 163805 47866 164125 47898
rect 184874 48454 185194 48486
rect 184874 48218 184916 48454
rect 185152 48218 185194 48454
rect 184874 48134 185194 48218
rect 184874 47898 184916 48134
rect 185152 47898 185194 48134
rect 184874 47866 185194 47898
rect 190805 48454 191125 48486
rect 190805 48218 190847 48454
rect 191083 48218 191125 48454
rect 190805 48134 191125 48218
rect 190805 47898 190847 48134
rect 191083 47898 191125 48134
rect 190805 47866 191125 47898
rect 211874 48454 212194 48486
rect 211874 48218 211916 48454
rect 212152 48218 212194 48454
rect 211874 48134 212194 48218
rect 211874 47898 211916 48134
rect 212152 47898 212194 48134
rect 211874 47866 212194 47898
rect 217805 48454 218125 48486
rect 217805 48218 217847 48454
rect 218083 48218 218125 48454
rect 217805 48134 218125 48218
rect 217805 47898 217847 48134
rect 218083 47898 218125 48134
rect 217805 47866 218125 47898
rect 238874 48454 239194 48486
rect 238874 48218 238916 48454
rect 239152 48218 239194 48454
rect 238874 48134 239194 48218
rect 238874 47898 238916 48134
rect 239152 47898 239194 48134
rect 238874 47866 239194 47898
rect 244805 48454 245125 48486
rect 244805 48218 244847 48454
rect 245083 48218 245125 48454
rect 244805 48134 245125 48218
rect 244805 47898 244847 48134
rect 245083 47898 245125 48134
rect 244805 47866 245125 47898
rect 265874 48454 266194 48486
rect 265874 48218 265916 48454
rect 266152 48218 266194 48454
rect 265874 48134 266194 48218
rect 265874 47898 265916 48134
rect 266152 47898 266194 48134
rect 265874 47866 266194 47898
rect 271805 48454 272125 48486
rect 271805 48218 271847 48454
rect 272083 48218 272125 48454
rect 271805 48134 272125 48218
rect 271805 47898 271847 48134
rect 272083 47898 272125 48134
rect 271805 47866 272125 47898
rect 292874 48454 293194 48486
rect 292874 48218 292916 48454
rect 293152 48218 293194 48454
rect 292874 48134 293194 48218
rect 292874 47898 292916 48134
rect 293152 47898 293194 48134
rect 292874 47866 293194 47898
rect 298805 48454 299125 48486
rect 298805 48218 298847 48454
rect 299083 48218 299125 48454
rect 298805 48134 299125 48218
rect 298805 47898 298847 48134
rect 299083 47898 299125 48134
rect 298805 47866 299125 47898
rect 319874 48454 320194 48486
rect 319874 48218 319916 48454
rect 320152 48218 320194 48454
rect 319874 48134 320194 48218
rect 319874 47898 319916 48134
rect 320152 47898 320194 48134
rect 319874 47866 320194 47898
rect 325805 48454 326125 48486
rect 325805 48218 325847 48454
rect 326083 48218 326125 48454
rect 325805 48134 326125 48218
rect 325805 47898 325847 48134
rect 326083 47898 326125 48134
rect 325805 47866 326125 47898
rect 346874 48454 347194 48486
rect 346874 48218 346916 48454
rect 347152 48218 347194 48454
rect 346874 48134 347194 48218
rect 346874 47898 346916 48134
rect 347152 47898 347194 48134
rect 346874 47866 347194 47898
rect 352805 48454 353125 48486
rect 352805 48218 352847 48454
rect 353083 48218 353125 48454
rect 352805 48134 353125 48218
rect 352805 47898 352847 48134
rect 353083 47898 353125 48134
rect 352805 47866 353125 47898
rect 373874 48454 374194 48486
rect 373874 48218 373916 48454
rect 374152 48218 374194 48454
rect 373874 48134 374194 48218
rect 373874 47898 373916 48134
rect 374152 47898 374194 48134
rect 373874 47866 374194 47898
rect 379805 48454 380125 48486
rect 379805 48218 379847 48454
rect 380083 48218 380125 48454
rect 379805 48134 380125 48218
rect 379805 47898 379847 48134
rect 380083 47898 380125 48134
rect 379805 47866 380125 47898
rect 400874 48454 401194 48486
rect 400874 48218 400916 48454
rect 401152 48218 401194 48454
rect 400874 48134 401194 48218
rect 400874 47898 400916 48134
rect 401152 47898 401194 48134
rect 400874 47866 401194 47898
rect 406805 48454 407125 48486
rect 406805 48218 406847 48454
rect 407083 48218 407125 48454
rect 406805 48134 407125 48218
rect 406805 47898 406847 48134
rect 407083 47898 407125 48134
rect 406805 47866 407125 47898
rect 427874 48454 428194 48486
rect 427874 48218 427916 48454
rect 428152 48218 428194 48454
rect 427874 48134 428194 48218
rect 427874 47898 427916 48134
rect 428152 47898 428194 48134
rect 427874 47866 428194 47898
rect 433805 48454 434125 48486
rect 433805 48218 433847 48454
rect 434083 48218 434125 48454
rect 433805 48134 434125 48218
rect 433805 47898 433847 48134
rect 434083 47898 434125 48134
rect 433805 47866 434125 47898
rect 454874 48454 455194 48486
rect 454874 48218 454916 48454
rect 455152 48218 455194 48454
rect 454874 48134 455194 48218
rect 454874 47898 454916 48134
rect 455152 47898 455194 48134
rect 454874 47866 455194 47898
rect 460805 48454 461125 48486
rect 460805 48218 460847 48454
rect 461083 48218 461125 48454
rect 460805 48134 461125 48218
rect 460805 47898 460847 48134
rect 461083 47898 461125 48134
rect 460805 47866 461125 47898
rect 481874 48454 482194 48486
rect 481874 48218 481916 48454
rect 482152 48218 482194 48454
rect 481874 48134 482194 48218
rect 481874 47898 481916 48134
rect 482152 47898 482194 48134
rect 481874 47866 482194 47898
rect 487805 48454 488125 48486
rect 487805 48218 487847 48454
rect 488083 48218 488125 48454
rect 487805 48134 488125 48218
rect 487805 47898 487847 48134
rect 488083 47898 488125 48134
rect 487805 47866 488125 47898
rect 508874 48454 509194 48486
rect 508874 48218 508916 48454
rect 509152 48218 509194 48454
rect 508874 48134 509194 48218
rect 508874 47898 508916 48134
rect 509152 47898 509194 48134
rect 508874 47866 509194 47898
rect 514805 48454 515125 48486
rect 514805 48218 514847 48454
rect 515083 48218 515125 48454
rect 514805 48134 515125 48218
rect 514805 47898 514847 48134
rect 515083 47898 515125 48134
rect 514805 47866 515125 47898
rect 535874 48454 536194 48486
rect 535874 48218 535916 48454
rect 536152 48218 536194 48454
rect 535874 48134 536194 48218
rect 535874 47898 535916 48134
rect 536152 47898 536194 48134
rect 535874 47866 536194 47898
rect 541805 48454 542125 48486
rect 541805 48218 541847 48454
rect 542083 48218 542125 48454
rect 541805 48134 542125 48218
rect 541805 47898 541847 48134
rect 542083 47898 542125 48134
rect 541805 47866 542125 47898
rect 19794 39454 20414 41000
rect 19794 39218 19826 39454
rect 20062 39218 20146 39454
rect 20382 39218 20414 39454
rect 19794 39134 20414 39218
rect 19794 38898 19826 39134
rect 20062 38898 20146 39134
rect 20382 38898 20414 39134
rect 19794 38000 20414 38898
rect 28794 40394 29414 41000
rect 28794 40158 28826 40394
rect 29062 40158 29146 40394
rect 29382 40158 29414 40394
rect 28794 40074 29414 40158
rect 28794 39838 28826 40074
rect 29062 39838 29146 40074
rect 29382 39838 29414 40074
rect 28794 38000 29414 39838
rect 37794 39454 38414 41000
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 38000 38414 38898
rect 46794 40394 47414 41000
rect 46794 40158 46826 40394
rect 47062 40158 47146 40394
rect 47382 40158 47414 40394
rect 46794 40074 47414 40158
rect 46794 39838 46826 40074
rect 47062 39838 47146 40074
rect 47382 39838 47414 40074
rect 46794 38000 47414 39838
rect 55794 39454 56414 41000
rect 55794 39218 55826 39454
rect 56062 39218 56146 39454
rect 56382 39218 56414 39454
rect 55794 39134 56414 39218
rect 55794 38898 55826 39134
rect 56062 38898 56146 39134
rect 56382 38898 56414 39134
rect 55794 38000 56414 38898
rect 64794 40394 65414 41000
rect 64794 40158 64826 40394
rect 65062 40158 65146 40394
rect 65382 40158 65414 40394
rect 64794 40074 65414 40158
rect 64794 39838 64826 40074
rect 65062 39838 65146 40074
rect 65382 39838 65414 40074
rect 64794 38000 65414 39838
rect 73794 39454 74414 41000
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 38000 74414 38898
rect 82794 40394 83414 41000
rect 82794 40158 82826 40394
rect 83062 40158 83146 40394
rect 83382 40158 83414 40394
rect 82794 40074 83414 40158
rect 82794 39838 82826 40074
rect 83062 39838 83146 40074
rect 83382 39838 83414 40074
rect 82794 38000 83414 39838
rect 91794 39454 92414 41000
rect 91794 39218 91826 39454
rect 92062 39218 92146 39454
rect 92382 39218 92414 39454
rect 91794 39134 92414 39218
rect 91794 38898 91826 39134
rect 92062 38898 92146 39134
rect 92382 38898 92414 39134
rect 91794 38000 92414 38898
rect 100794 40394 101414 41000
rect 100794 40158 100826 40394
rect 101062 40158 101146 40394
rect 101382 40158 101414 40394
rect 100794 40074 101414 40158
rect 100794 39838 100826 40074
rect 101062 39838 101146 40074
rect 101382 39838 101414 40074
rect 100794 38000 101414 39838
rect 109794 39454 110414 41000
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 38000 110414 38898
rect 118794 40394 119414 41000
rect 118794 40158 118826 40394
rect 119062 40158 119146 40394
rect 119382 40158 119414 40394
rect 118794 40074 119414 40158
rect 118794 39838 118826 40074
rect 119062 39838 119146 40074
rect 119382 39838 119414 40074
rect 118794 38000 119414 39838
rect 127794 39454 128414 41000
rect 127794 39218 127826 39454
rect 128062 39218 128146 39454
rect 128382 39218 128414 39454
rect 127794 39134 128414 39218
rect 127794 38898 127826 39134
rect 128062 38898 128146 39134
rect 128382 38898 128414 39134
rect 127794 38000 128414 38898
rect 136794 40394 137414 41000
rect 136794 40158 136826 40394
rect 137062 40158 137146 40394
rect 137382 40158 137414 40394
rect 136794 40074 137414 40158
rect 136794 39838 136826 40074
rect 137062 39838 137146 40074
rect 137382 39838 137414 40074
rect 136794 38000 137414 39838
rect 145794 39454 146414 41000
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 38000 146414 38898
rect 154794 40394 155414 41000
rect 154794 40158 154826 40394
rect 155062 40158 155146 40394
rect 155382 40158 155414 40394
rect 154794 40074 155414 40158
rect 154794 39838 154826 40074
rect 155062 39838 155146 40074
rect 155382 39838 155414 40074
rect 154794 38000 155414 39838
rect 163794 39454 164414 41000
rect 163794 39218 163826 39454
rect 164062 39218 164146 39454
rect 164382 39218 164414 39454
rect 163794 39134 164414 39218
rect 163794 38898 163826 39134
rect 164062 38898 164146 39134
rect 164382 38898 164414 39134
rect 163794 38000 164414 38898
rect 172794 40394 173414 41000
rect 172794 40158 172826 40394
rect 173062 40158 173146 40394
rect 173382 40158 173414 40394
rect 172794 40074 173414 40158
rect 172794 39838 172826 40074
rect 173062 39838 173146 40074
rect 173382 39838 173414 40074
rect 172794 38000 173414 39838
rect 181794 39454 182414 41000
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 38000 182414 38898
rect 190794 40394 191414 41000
rect 190794 40158 190826 40394
rect 191062 40158 191146 40394
rect 191382 40158 191414 40394
rect 190794 40074 191414 40158
rect 190794 39838 190826 40074
rect 191062 39838 191146 40074
rect 191382 39838 191414 40074
rect 190794 38000 191414 39838
rect 199794 39454 200414 41000
rect 199794 39218 199826 39454
rect 200062 39218 200146 39454
rect 200382 39218 200414 39454
rect 199794 39134 200414 39218
rect 199794 38898 199826 39134
rect 200062 38898 200146 39134
rect 200382 38898 200414 39134
rect 199794 38000 200414 38898
rect 208794 40394 209414 41000
rect 208794 40158 208826 40394
rect 209062 40158 209146 40394
rect 209382 40158 209414 40394
rect 208794 40074 209414 40158
rect 208794 39838 208826 40074
rect 209062 39838 209146 40074
rect 209382 39838 209414 40074
rect 208794 38000 209414 39838
rect 217794 39454 218414 41000
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 38000 218414 38898
rect 226794 40394 227414 41000
rect 226794 40158 226826 40394
rect 227062 40158 227146 40394
rect 227382 40158 227414 40394
rect 226794 40074 227414 40158
rect 226794 39838 226826 40074
rect 227062 39838 227146 40074
rect 227382 39838 227414 40074
rect 226794 38000 227414 39838
rect 235794 39454 236414 41000
rect 235794 39218 235826 39454
rect 236062 39218 236146 39454
rect 236382 39218 236414 39454
rect 235794 39134 236414 39218
rect 235794 38898 235826 39134
rect 236062 38898 236146 39134
rect 236382 38898 236414 39134
rect 235794 38000 236414 38898
rect 244794 40394 245414 41000
rect 244794 40158 244826 40394
rect 245062 40158 245146 40394
rect 245382 40158 245414 40394
rect 244794 40074 245414 40158
rect 244794 39838 244826 40074
rect 245062 39838 245146 40074
rect 245382 39838 245414 40074
rect 244794 38000 245414 39838
rect 253794 39454 254414 41000
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 38000 254414 38898
rect 262794 40394 263414 41000
rect 262794 40158 262826 40394
rect 263062 40158 263146 40394
rect 263382 40158 263414 40394
rect 262794 40074 263414 40158
rect 262794 39838 262826 40074
rect 263062 39838 263146 40074
rect 263382 39838 263414 40074
rect 262794 38000 263414 39838
rect 271794 39454 272414 41000
rect 271794 39218 271826 39454
rect 272062 39218 272146 39454
rect 272382 39218 272414 39454
rect 271794 39134 272414 39218
rect 271794 38898 271826 39134
rect 272062 38898 272146 39134
rect 272382 38898 272414 39134
rect 271794 38000 272414 38898
rect 280794 40394 281414 41000
rect 280794 40158 280826 40394
rect 281062 40158 281146 40394
rect 281382 40158 281414 40394
rect 280794 40074 281414 40158
rect 280794 39838 280826 40074
rect 281062 39838 281146 40074
rect 281382 39838 281414 40074
rect 280794 38000 281414 39838
rect 289794 39454 290414 41000
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 38000 290414 38898
rect 298794 40394 299414 41000
rect 298794 40158 298826 40394
rect 299062 40158 299146 40394
rect 299382 40158 299414 40394
rect 298794 40074 299414 40158
rect 298794 39838 298826 40074
rect 299062 39838 299146 40074
rect 299382 39838 299414 40074
rect 298794 38000 299414 39838
rect 307794 39454 308414 41000
rect 307794 39218 307826 39454
rect 308062 39218 308146 39454
rect 308382 39218 308414 39454
rect 307794 39134 308414 39218
rect 307794 38898 307826 39134
rect 308062 38898 308146 39134
rect 308382 38898 308414 39134
rect 307794 38000 308414 38898
rect 316794 40394 317414 41000
rect 316794 40158 316826 40394
rect 317062 40158 317146 40394
rect 317382 40158 317414 40394
rect 316794 40074 317414 40158
rect 316794 39838 316826 40074
rect 317062 39838 317146 40074
rect 317382 39838 317414 40074
rect 316794 38000 317414 39838
rect 325794 39454 326414 41000
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 38000 326414 38898
rect 334794 40394 335414 41000
rect 334794 40158 334826 40394
rect 335062 40158 335146 40394
rect 335382 40158 335414 40394
rect 334794 40074 335414 40158
rect 334794 39838 334826 40074
rect 335062 39838 335146 40074
rect 335382 39838 335414 40074
rect 334794 38000 335414 39838
rect 343794 39454 344414 41000
rect 343794 39218 343826 39454
rect 344062 39218 344146 39454
rect 344382 39218 344414 39454
rect 343794 39134 344414 39218
rect 343794 38898 343826 39134
rect 344062 38898 344146 39134
rect 344382 38898 344414 39134
rect 343794 38000 344414 38898
rect 352794 40394 353414 41000
rect 352794 40158 352826 40394
rect 353062 40158 353146 40394
rect 353382 40158 353414 40394
rect 352794 40074 353414 40158
rect 352794 39838 352826 40074
rect 353062 39838 353146 40074
rect 353382 39838 353414 40074
rect 352794 38000 353414 39838
rect 361794 39454 362414 41000
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 38000 362414 38898
rect 370794 40394 371414 41000
rect 370794 40158 370826 40394
rect 371062 40158 371146 40394
rect 371382 40158 371414 40394
rect 370794 40074 371414 40158
rect 370794 39838 370826 40074
rect 371062 39838 371146 40074
rect 371382 39838 371414 40074
rect 370794 38000 371414 39838
rect 379794 39454 380414 41000
rect 379794 39218 379826 39454
rect 380062 39218 380146 39454
rect 380382 39218 380414 39454
rect 379794 39134 380414 39218
rect 379794 38898 379826 39134
rect 380062 38898 380146 39134
rect 380382 38898 380414 39134
rect 379794 38000 380414 38898
rect 388794 40394 389414 41000
rect 388794 40158 388826 40394
rect 389062 40158 389146 40394
rect 389382 40158 389414 40394
rect 388794 40074 389414 40158
rect 388794 39838 388826 40074
rect 389062 39838 389146 40074
rect 389382 39838 389414 40074
rect 388794 38000 389414 39838
rect 397794 39454 398414 41000
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 38000 398414 38898
rect 406794 40394 407414 41000
rect 406794 40158 406826 40394
rect 407062 40158 407146 40394
rect 407382 40158 407414 40394
rect 406794 40074 407414 40158
rect 406794 39838 406826 40074
rect 407062 39838 407146 40074
rect 407382 39838 407414 40074
rect 406794 38000 407414 39838
rect 415794 39454 416414 41000
rect 415794 39218 415826 39454
rect 416062 39218 416146 39454
rect 416382 39218 416414 39454
rect 415794 39134 416414 39218
rect 415794 38898 415826 39134
rect 416062 38898 416146 39134
rect 416382 38898 416414 39134
rect 415794 38000 416414 38898
rect 424794 40394 425414 41000
rect 424794 40158 424826 40394
rect 425062 40158 425146 40394
rect 425382 40158 425414 40394
rect 424794 40074 425414 40158
rect 424794 39838 424826 40074
rect 425062 39838 425146 40074
rect 425382 39838 425414 40074
rect 424794 38000 425414 39838
rect 433794 39454 434414 41000
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 38000 434414 38898
rect 442794 40394 443414 41000
rect 442794 40158 442826 40394
rect 443062 40158 443146 40394
rect 443382 40158 443414 40394
rect 442794 40074 443414 40158
rect 442794 39838 442826 40074
rect 443062 39838 443146 40074
rect 443382 39838 443414 40074
rect 442794 38000 443414 39838
rect 451794 39454 452414 41000
rect 451794 39218 451826 39454
rect 452062 39218 452146 39454
rect 452382 39218 452414 39454
rect 451794 39134 452414 39218
rect 451794 38898 451826 39134
rect 452062 38898 452146 39134
rect 452382 38898 452414 39134
rect 451794 38000 452414 38898
rect 460794 40394 461414 41000
rect 460794 40158 460826 40394
rect 461062 40158 461146 40394
rect 461382 40158 461414 40394
rect 460794 40074 461414 40158
rect 460794 39838 460826 40074
rect 461062 39838 461146 40074
rect 461382 39838 461414 40074
rect 460794 38000 461414 39838
rect 469794 39454 470414 41000
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 38000 470414 38898
rect 478794 40394 479414 41000
rect 478794 40158 478826 40394
rect 479062 40158 479146 40394
rect 479382 40158 479414 40394
rect 478794 40074 479414 40158
rect 478794 39838 478826 40074
rect 479062 39838 479146 40074
rect 479382 39838 479414 40074
rect 478794 38000 479414 39838
rect 487794 39454 488414 41000
rect 487794 39218 487826 39454
rect 488062 39218 488146 39454
rect 488382 39218 488414 39454
rect 487794 39134 488414 39218
rect 487794 38898 487826 39134
rect 488062 38898 488146 39134
rect 488382 38898 488414 39134
rect 487794 38000 488414 38898
rect 496794 40394 497414 41000
rect 496794 40158 496826 40394
rect 497062 40158 497146 40394
rect 497382 40158 497414 40394
rect 496794 40074 497414 40158
rect 496794 39838 496826 40074
rect 497062 39838 497146 40074
rect 497382 39838 497414 40074
rect 496794 38000 497414 39838
rect 505794 39454 506414 41000
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 38000 506414 38898
rect 514794 40394 515414 41000
rect 514794 40158 514826 40394
rect 515062 40158 515146 40394
rect 515382 40158 515414 40394
rect 514794 40074 515414 40158
rect 514794 39838 514826 40074
rect 515062 39838 515146 40074
rect 515382 39838 515414 40074
rect 514794 38000 515414 39838
rect 523794 39454 524414 41000
rect 523794 39218 523826 39454
rect 524062 39218 524146 39454
rect 524382 39218 524414 39454
rect 523794 39134 524414 39218
rect 523794 38898 523826 39134
rect 524062 38898 524146 39134
rect 524382 38898 524414 39134
rect 523794 38000 524414 38898
rect 532794 40394 533414 41000
rect 532794 40158 532826 40394
rect 533062 40158 533146 40394
rect 533382 40158 533414 40394
rect 532794 40074 533414 40158
rect 532794 39838 532826 40074
rect 533062 39838 533146 40074
rect 533382 39838 533414 40074
rect 532794 38000 533414 39838
rect 541794 39454 542414 41000
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 38000 542414 38898
rect 550794 40394 551414 41000
rect 550794 40158 550826 40394
rect 551062 40158 551146 40394
rect 551382 40158 551414 40394
rect 550794 40074 551414 40158
rect 550794 39838 550826 40074
rect 551062 39838 551146 40074
rect 551382 39838 551414 40074
rect 550794 38000 551414 39838
rect 559794 39454 560414 56898
rect 559794 39218 559826 39454
rect 560062 39218 560146 39454
rect 560382 39218 560414 39454
rect 559794 39134 560414 39218
rect 559794 38898 559826 39134
rect 560062 38898 560146 39134
rect 560382 38898 560414 39134
rect 10794 30218 10826 30454
rect 11062 30218 11146 30454
rect 11382 30218 11414 30454
rect 10794 30134 11414 30218
rect 10794 29898 10826 30134
rect 11062 29898 11146 30134
rect 11382 29898 11414 30134
rect 10794 12454 11414 29898
rect 22874 30454 23194 30486
rect 22874 30218 22916 30454
rect 23152 30218 23194 30454
rect 22874 30134 23194 30218
rect 22874 29898 22916 30134
rect 23152 29898 23194 30134
rect 22874 29866 23194 29898
rect 28805 30454 29125 30486
rect 28805 30218 28847 30454
rect 29083 30218 29125 30454
rect 28805 30134 29125 30218
rect 28805 29898 28847 30134
rect 29083 29898 29125 30134
rect 28805 29866 29125 29898
rect 49874 30454 50194 30486
rect 49874 30218 49916 30454
rect 50152 30218 50194 30454
rect 49874 30134 50194 30218
rect 49874 29898 49916 30134
rect 50152 29898 50194 30134
rect 49874 29866 50194 29898
rect 55805 30454 56125 30486
rect 55805 30218 55847 30454
rect 56083 30218 56125 30454
rect 55805 30134 56125 30218
rect 55805 29898 55847 30134
rect 56083 29898 56125 30134
rect 55805 29866 56125 29898
rect 76874 30454 77194 30486
rect 76874 30218 76916 30454
rect 77152 30218 77194 30454
rect 76874 30134 77194 30218
rect 76874 29898 76916 30134
rect 77152 29898 77194 30134
rect 76874 29866 77194 29898
rect 82805 30454 83125 30486
rect 82805 30218 82847 30454
rect 83083 30218 83125 30454
rect 82805 30134 83125 30218
rect 82805 29898 82847 30134
rect 83083 29898 83125 30134
rect 82805 29866 83125 29898
rect 103874 30454 104194 30486
rect 103874 30218 103916 30454
rect 104152 30218 104194 30454
rect 103874 30134 104194 30218
rect 103874 29898 103916 30134
rect 104152 29898 104194 30134
rect 103874 29866 104194 29898
rect 109805 30454 110125 30486
rect 109805 30218 109847 30454
rect 110083 30218 110125 30454
rect 109805 30134 110125 30218
rect 109805 29898 109847 30134
rect 110083 29898 110125 30134
rect 109805 29866 110125 29898
rect 130874 30454 131194 30486
rect 130874 30218 130916 30454
rect 131152 30218 131194 30454
rect 130874 30134 131194 30218
rect 130874 29898 130916 30134
rect 131152 29898 131194 30134
rect 130874 29866 131194 29898
rect 136805 30454 137125 30486
rect 136805 30218 136847 30454
rect 137083 30218 137125 30454
rect 136805 30134 137125 30218
rect 136805 29898 136847 30134
rect 137083 29898 137125 30134
rect 136805 29866 137125 29898
rect 157874 30454 158194 30486
rect 157874 30218 157916 30454
rect 158152 30218 158194 30454
rect 157874 30134 158194 30218
rect 157874 29898 157916 30134
rect 158152 29898 158194 30134
rect 157874 29866 158194 29898
rect 163805 30454 164125 30486
rect 163805 30218 163847 30454
rect 164083 30218 164125 30454
rect 163805 30134 164125 30218
rect 163805 29898 163847 30134
rect 164083 29898 164125 30134
rect 163805 29866 164125 29898
rect 184874 30454 185194 30486
rect 184874 30218 184916 30454
rect 185152 30218 185194 30454
rect 184874 30134 185194 30218
rect 184874 29898 184916 30134
rect 185152 29898 185194 30134
rect 184874 29866 185194 29898
rect 190805 30454 191125 30486
rect 190805 30218 190847 30454
rect 191083 30218 191125 30454
rect 190805 30134 191125 30218
rect 190805 29898 190847 30134
rect 191083 29898 191125 30134
rect 190805 29866 191125 29898
rect 211874 30454 212194 30486
rect 211874 30218 211916 30454
rect 212152 30218 212194 30454
rect 211874 30134 212194 30218
rect 211874 29898 211916 30134
rect 212152 29898 212194 30134
rect 211874 29866 212194 29898
rect 217805 30454 218125 30486
rect 217805 30218 217847 30454
rect 218083 30218 218125 30454
rect 217805 30134 218125 30218
rect 217805 29898 217847 30134
rect 218083 29898 218125 30134
rect 217805 29866 218125 29898
rect 238874 30454 239194 30486
rect 238874 30218 238916 30454
rect 239152 30218 239194 30454
rect 238874 30134 239194 30218
rect 238874 29898 238916 30134
rect 239152 29898 239194 30134
rect 238874 29866 239194 29898
rect 244805 30454 245125 30486
rect 244805 30218 244847 30454
rect 245083 30218 245125 30454
rect 244805 30134 245125 30218
rect 244805 29898 244847 30134
rect 245083 29898 245125 30134
rect 244805 29866 245125 29898
rect 265874 30454 266194 30486
rect 265874 30218 265916 30454
rect 266152 30218 266194 30454
rect 265874 30134 266194 30218
rect 265874 29898 265916 30134
rect 266152 29898 266194 30134
rect 265874 29866 266194 29898
rect 271805 30454 272125 30486
rect 271805 30218 271847 30454
rect 272083 30218 272125 30454
rect 271805 30134 272125 30218
rect 271805 29898 271847 30134
rect 272083 29898 272125 30134
rect 271805 29866 272125 29898
rect 292874 30454 293194 30486
rect 292874 30218 292916 30454
rect 293152 30218 293194 30454
rect 292874 30134 293194 30218
rect 292874 29898 292916 30134
rect 293152 29898 293194 30134
rect 292874 29866 293194 29898
rect 298805 30454 299125 30486
rect 298805 30218 298847 30454
rect 299083 30218 299125 30454
rect 298805 30134 299125 30218
rect 298805 29898 298847 30134
rect 299083 29898 299125 30134
rect 298805 29866 299125 29898
rect 319874 30454 320194 30486
rect 319874 30218 319916 30454
rect 320152 30218 320194 30454
rect 319874 30134 320194 30218
rect 319874 29898 319916 30134
rect 320152 29898 320194 30134
rect 319874 29866 320194 29898
rect 325805 30454 326125 30486
rect 325805 30218 325847 30454
rect 326083 30218 326125 30454
rect 325805 30134 326125 30218
rect 325805 29898 325847 30134
rect 326083 29898 326125 30134
rect 325805 29866 326125 29898
rect 346874 30454 347194 30486
rect 346874 30218 346916 30454
rect 347152 30218 347194 30454
rect 346874 30134 347194 30218
rect 346874 29898 346916 30134
rect 347152 29898 347194 30134
rect 346874 29866 347194 29898
rect 352805 30454 353125 30486
rect 352805 30218 352847 30454
rect 353083 30218 353125 30454
rect 352805 30134 353125 30218
rect 352805 29898 352847 30134
rect 353083 29898 353125 30134
rect 352805 29866 353125 29898
rect 373874 30454 374194 30486
rect 373874 30218 373916 30454
rect 374152 30218 374194 30454
rect 373874 30134 374194 30218
rect 373874 29898 373916 30134
rect 374152 29898 374194 30134
rect 373874 29866 374194 29898
rect 379805 30454 380125 30486
rect 379805 30218 379847 30454
rect 380083 30218 380125 30454
rect 379805 30134 380125 30218
rect 379805 29898 379847 30134
rect 380083 29898 380125 30134
rect 379805 29866 380125 29898
rect 400874 30454 401194 30486
rect 400874 30218 400916 30454
rect 401152 30218 401194 30454
rect 400874 30134 401194 30218
rect 400874 29898 400916 30134
rect 401152 29898 401194 30134
rect 400874 29866 401194 29898
rect 406805 30454 407125 30486
rect 406805 30218 406847 30454
rect 407083 30218 407125 30454
rect 406805 30134 407125 30218
rect 406805 29898 406847 30134
rect 407083 29898 407125 30134
rect 406805 29866 407125 29898
rect 427874 30454 428194 30486
rect 427874 30218 427916 30454
rect 428152 30218 428194 30454
rect 427874 30134 428194 30218
rect 427874 29898 427916 30134
rect 428152 29898 428194 30134
rect 427874 29866 428194 29898
rect 433805 30454 434125 30486
rect 433805 30218 433847 30454
rect 434083 30218 434125 30454
rect 433805 30134 434125 30218
rect 433805 29898 433847 30134
rect 434083 29898 434125 30134
rect 433805 29866 434125 29898
rect 454874 30454 455194 30486
rect 454874 30218 454916 30454
rect 455152 30218 455194 30454
rect 454874 30134 455194 30218
rect 454874 29898 454916 30134
rect 455152 29898 455194 30134
rect 454874 29866 455194 29898
rect 460805 30454 461125 30486
rect 460805 30218 460847 30454
rect 461083 30218 461125 30454
rect 460805 30134 461125 30218
rect 460805 29898 460847 30134
rect 461083 29898 461125 30134
rect 460805 29866 461125 29898
rect 481874 30454 482194 30486
rect 481874 30218 481916 30454
rect 482152 30218 482194 30454
rect 481874 30134 482194 30218
rect 481874 29898 481916 30134
rect 482152 29898 482194 30134
rect 481874 29866 482194 29898
rect 487805 30454 488125 30486
rect 487805 30218 487847 30454
rect 488083 30218 488125 30454
rect 487805 30134 488125 30218
rect 487805 29898 487847 30134
rect 488083 29898 488125 30134
rect 487805 29866 488125 29898
rect 508874 30454 509194 30486
rect 508874 30218 508916 30454
rect 509152 30218 509194 30454
rect 508874 30134 509194 30218
rect 508874 29898 508916 30134
rect 509152 29898 509194 30134
rect 508874 29866 509194 29898
rect 514805 30454 515125 30486
rect 514805 30218 514847 30454
rect 515083 30218 515125 30454
rect 514805 30134 515125 30218
rect 514805 29898 514847 30134
rect 515083 29898 515125 30134
rect 514805 29866 515125 29898
rect 535874 30454 536194 30486
rect 535874 30218 535916 30454
rect 536152 30218 536194 30454
rect 535874 30134 536194 30218
rect 535874 29898 535916 30134
rect 536152 29898 536194 30134
rect 535874 29866 536194 29898
rect 541805 30454 542125 30486
rect 541805 30218 541847 30454
rect 542083 30218 542125 30454
rect 541805 30134 542125 30218
rect 541805 29898 541847 30134
rect 542083 29898 542125 30134
rect 541805 29866 542125 29898
rect 19910 21454 20230 21486
rect 19910 21218 19952 21454
rect 20188 21218 20230 21454
rect 19910 21134 20230 21218
rect 19910 20898 19952 21134
rect 20188 20898 20230 21134
rect 19910 20866 20230 20898
rect 25840 21454 26160 21486
rect 25840 21218 25882 21454
rect 26118 21218 26160 21454
rect 25840 21134 26160 21218
rect 25840 20898 25882 21134
rect 26118 20898 26160 21134
rect 25840 20866 26160 20898
rect 31771 21454 32091 21486
rect 31771 21218 31813 21454
rect 32049 21218 32091 21454
rect 31771 21134 32091 21218
rect 31771 20898 31813 21134
rect 32049 20898 32091 21134
rect 31771 20866 32091 20898
rect 46910 21454 47230 21486
rect 46910 21218 46952 21454
rect 47188 21218 47230 21454
rect 46910 21134 47230 21218
rect 46910 20898 46952 21134
rect 47188 20898 47230 21134
rect 46910 20866 47230 20898
rect 52840 21454 53160 21486
rect 52840 21218 52882 21454
rect 53118 21218 53160 21454
rect 52840 21134 53160 21218
rect 52840 20898 52882 21134
rect 53118 20898 53160 21134
rect 52840 20866 53160 20898
rect 58771 21454 59091 21486
rect 58771 21218 58813 21454
rect 59049 21218 59091 21454
rect 58771 21134 59091 21218
rect 58771 20898 58813 21134
rect 59049 20898 59091 21134
rect 58771 20866 59091 20898
rect 73910 21454 74230 21486
rect 73910 21218 73952 21454
rect 74188 21218 74230 21454
rect 73910 21134 74230 21218
rect 73910 20898 73952 21134
rect 74188 20898 74230 21134
rect 73910 20866 74230 20898
rect 79840 21454 80160 21486
rect 79840 21218 79882 21454
rect 80118 21218 80160 21454
rect 79840 21134 80160 21218
rect 79840 20898 79882 21134
rect 80118 20898 80160 21134
rect 79840 20866 80160 20898
rect 85771 21454 86091 21486
rect 85771 21218 85813 21454
rect 86049 21218 86091 21454
rect 85771 21134 86091 21218
rect 85771 20898 85813 21134
rect 86049 20898 86091 21134
rect 85771 20866 86091 20898
rect 100910 21454 101230 21486
rect 100910 21218 100952 21454
rect 101188 21218 101230 21454
rect 100910 21134 101230 21218
rect 100910 20898 100952 21134
rect 101188 20898 101230 21134
rect 100910 20866 101230 20898
rect 106840 21454 107160 21486
rect 106840 21218 106882 21454
rect 107118 21218 107160 21454
rect 106840 21134 107160 21218
rect 106840 20898 106882 21134
rect 107118 20898 107160 21134
rect 106840 20866 107160 20898
rect 112771 21454 113091 21486
rect 112771 21218 112813 21454
rect 113049 21218 113091 21454
rect 112771 21134 113091 21218
rect 112771 20898 112813 21134
rect 113049 20898 113091 21134
rect 112771 20866 113091 20898
rect 127910 21454 128230 21486
rect 127910 21218 127952 21454
rect 128188 21218 128230 21454
rect 127910 21134 128230 21218
rect 127910 20898 127952 21134
rect 128188 20898 128230 21134
rect 127910 20866 128230 20898
rect 133840 21454 134160 21486
rect 133840 21218 133882 21454
rect 134118 21218 134160 21454
rect 133840 21134 134160 21218
rect 133840 20898 133882 21134
rect 134118 20898 134160 21134
rect 133840 20866 134160 20898
rect 139771 21454 140091 21486
rect 139771 21218 139813 21454
rect 140049 21218 140091 21454
rect 139771 21134 140091 21218
rect 139771 20898 139813 21134
rect 140049 20898 140091 21134
rect 139771 20866 140091 20898
rect 154910 21454 155230 21486
rect 154910 21218 154952 21454
rect 155188 21218 155230 21454
rect 154910 21134 155230 21218
rect 154910 20898 154952 21134
rect 155188 20898 155230 21134
rect 154910 20866 155230 20898
rect 160840 21454 161160 21486
rect 160840 21218 160882 21454
rect 161118 21218 161160 21454
rect 160840 21134 161160 21218
rect 160840 20898 160882 21134
rect 161118 20898 161160 21134
rect 160840 20866 161160 20898
rect 166771 21454 167091 21486
rect 166771 21218 166813 21454
rect 167049 21218 167091 21454
rect 166771 21134 167091 21218
rect 166771 20898 166813 21134
rect 167049 20898 167091 21134
rect 166771 20866 167091 20898
rect 181910 21454 182230 21486
rect 181910 21218 181952 21454
rect 182188 21218 182230 21454
rect 181910 21134 182230 21218
rect 181910 20898 181952 21134
rect 182188 20898 182230 21134
rect 181910 20866 182230 20898
rect 187840 21454 188160 21486
rect 187840 21218 187882 21454
rect 188118 21218 188160 21454
rect 187840 21134 188160 21218
rect 187840 20898 187882 21134
rect 188118 20898 188160 21134
rect 187840 20866 188160 20898
rect 193771 21454 194091 21486
rect 193771 21218 193813 21454
rect 194049 21218 194091 21454
rect 193771 21134 194091 21218
rect 193771 20898 193813 21134
rect 194049 20898 194091 21134
rect 193771 20866 194091 20898
rect 208910 21454 209230 21486
rect 208910 21218 208952 21454
rect 209188 21218 209230 21454
rect 208910 21134 209230 21218
rect 208910 20898 208952 21134
rect 209188 20898 209230 21134
rect 208910 20866 209230 20898
rect 214840 21454 215160 21486
rect 214840 21218 214882 21454
rect 215118 21218 215160 21454
rect 214840 21134 215160 21218
rect 214840 20898 214882 21134
rect 215118 20898 215160 21134
rect 214840 20866 215160 20898
rect 220771 21454 221091 21486
rect 220771 21218 220813 21454
rect 221049 21218 221091 21454
rect 220771 21134 221091 21218
rect 220771 20898 220813 21134
rect 221049 20898 221091 21134
rect 220771 20866 221091 20898
rect 235910 21454 236230 21486
rect 235910 21218 235952 21454
rect 236188 21218 236230 21454
rect 235910 21134 236230 21218
rect 235910 20898 235952 21134
rect 236188 20898 236230 21134
rect 235910 20866 236230 20898
rect 241840 21454 242160 21486
rect 241840 21218 241882 21454
rect 242118 21218 242160 21454
rect 241840 21134 242160 21218
rect 241840 20898 241882 21134
rect 242118 20898 242160 21134
rect 241840 20866 242160 20898
rect 247771 21454 248091 21486
rect 247771 21218 247813 21454
rect 248049 21218 248091 21454
rect 247771 21134 248091 21218
rect 247771 20898 247813 21134
rect 248049 20898 248091 21134
rect 247771 20866 248091 20898
rect 262910 21454 263230 21486
rect 262910 21218 262952 21454
rect 263188 21218 263230 21454
rect 262910 21134 263230 21218
rect 262910 20898 262952 21134
rect 263188 20898 263230 21134
rect 262910 20866 263230 20898
rect 268840 21454 269160 21486
rect 268840 21218 268882 21454
rect 269118 21218 269160 21454
rect 268840 21134 269160 21218
rect 268840 20898 268882 21134
rect 269118 20898 269160 21134
rect 268840 20866 269160 20898
rect 274771 21454 275091 21486
rect 274771 21218 274813 21454
rect 275049 21218 275091 21454
rect 274771 21134 275091 21218
rect 274771 20898 274813 21134
rect 275049 20898 275091 21134
rect 274771 20866 275091 20898
rect 289910 21454 290230 21486
rect 289910 21218 289952 21454
rect 290188 21218 290230 21454
rect 289910 21134 290230 21218
rect 289910 20898 289952 21134
rect 290188 20898 290230 21134
rect 289910 20866 290230 20898
rect 295840 21454 296160 21486
rect 295840 21218 295882 21454
rect 296118 21218 296160 21454
rect 295840 21134 296160 21218
rect 295840 20898 295882 21134
rect 296118 20898 296160 21134
rect 295840 20866 296160 20898
rect 301771 21454 302091 21486
rect 301771 21218 301813 21454
rect 302049 21218 302091 21454
rect 301771 21134 302091 21218
rect 301771 20898 301813 21134
rect 302049 20898 302091 21134
rect 301771 20866 302091 20898
rect 316910 21454 317230 21486
rect 316910 21218 316952 21454
rect 317188 21218 317230 21454
rect 316910 21134 317230 21218
rect 316910 20898 316952 21134
rect 317188 20898 317230 21134
rect 316910 20866 317230 20898
rect 322840 21454 323160 21486
rect 322840 21218 322882 21454
rect 323118 21218 323160 21454
rect 322840 21134 323160 21218
rect 322840 20898 322882 21134
rect 323118 20898 323160 21134
rect 322840 20866 323160 20898
rect 328771 21454 329091 21486
rect 328771 21218 328813 21454
rect 329049 21218 329091 21454
rect 328771 21134 329091 21218
rect 328771 20898 328813 21134
rect 329049 20898 329091 21134
rect 328771 20866 329091 20898
rect 343910 21454 344230 21486
rect 343910 21218 343952 21454
rect 344188 21218 344230 21454
rect 343910 21134 344230 21218
rect 343910 20898 343952 21134
rect 344188 20898 344230 21134
rect 343910 20866 344230 20898
rect 349840 21454 350160 21486
rect 349840 21218 349882 21454
rect 350118 21218 350160 21454
rect 349840 21134 350160 21218
rect 349840 20898 349882 21134
rect 350118 20898 350160 21134
rect 349840 20866 350160 20898
rect 355771 21454 356091 21486
rect 355771 21218 355813 21454
rect 356049 21218 356091 21454
rect 355771 21134 356091 21218
rect 355771 20898 355813 21134
rect 356049 20898 356091 21134
rect 355771 20866 356091 20898
rect 370910 21454 371230 21486
rect 370910 21218 370952 21454
rect 371188 21218 371230 21454
rect 370910 21134 371230 21218
rect 370910 20898 370952 21134
rect 371188 20898 371230 21134
rect 370910 20866 371230 20898
rect 376840 21454 377160 21486
rect 376840 21218 376882 21454
rect 377118 21218 377160 21454
rect 376840 21134 377160 21218
rect 376840 20898 376882 21134
rect 377118 20898 377160 21134
rect 376840 20866 377160 20898
rect 382771 21454 383091 21486
rect 382771 21218 382813 21454
rect 383049 21218 383091 21454
rect 382771 21134 383091 21218
rect 382771 20898 382813 21134
rect 383049 20898 383091 21134
rect 382771 20866 383091 20898
rect 397910 21454 398230 21486
rect 397910 21218 397952 21454
rect 398188 21218 398230 21454
rect 397910 21134 398230 21218
rect 397910 20898 397952 21134
rect 398188 20898 398230 21134
rect 397910 20866 398230 20898
rect 403840 21454 404160 21486
rect 403840 21218 403882 21454
rect 404118 21218 404160 21454
rect 403840 21134 404160 21218
rect 403840 20898 403882 21134
rect 404118 20898 404160 21134
rect 403840 20866 404160 20898
rect 409771 21454 410091 21486
rect 409771 21218 409813 21454
rect 410049 21218 410091 21454
rect 409771 21134 410091 21218
rect 409771 20898 409813 21134
rect 410049 20898 410091 21134
rect 409771 20866 410091 20898
rect 424910 21454 425230 21486
rect 424910 21218 424952 21454
rect 425188 21218 425230 21454
rect 424910 21134 425230 21218
rect 424910 20898 424952 21134
rect 425188 20898 425230 21134
rect 424910 20866 425230 20898
rect 430840 21454 431160 21486
rect 430840 21218 430882 21454
rect 431118 21218 431160 21454
rect 430840 21134 431160 21218
rect 430840 20898 430882 21134
rect 431118 20898 431160 21134
rect 430840 20866 431160 20898
rect 436771 21454 437091 21486
rect 436771 21218 436813 21454
rect 437049 21218 437091 21454
rect 436771 21134 437091 21218
rect 436771 20898 436813 21134
rect 437049 20898 437091 21134
rect 436771 20866 437091 20898
rect 451910 21454 452230 21486
rect 451910 21218 451952 21454
rect 452188 21218 452230 21454
rect 451910 21134 452230 21218
rect 451910 20898 451952 21134
rect 452188 20898 452230 21134
rect 451910 20866 452230 20898
rect 457840 21454 458160 21486
rect 457840 21218 457882 21454
rect 458118 21218 458160 21454
rect 457840 21134 458160 21218
rect 457840 20898 457882 21134
rect 458118 20898 458160 21134
rect 457840 20866 458160 20898
rect 463771 21454 464091 21486
rect 463771 21218 463813 21454
rect 464049 21218 464091 21454
rect 463771 21134 464091 21218
rect 463771 20898 463813 21134
rect 464049 20898 464091 21134
rect 463771 20866 464091 20898
rect 478910 21454 479230 21486
rect 478910 21218 478952 21454
rect 479188 21218 479230 21454
rect 478910 21134 479230 21218
rect 478910 20898 478952 21134
rect 479188 20898 479230 21134
rect 478910 20866 479230 20898
rect 484840 21454 485160 21486
rect 484840 21218 484882 21454
rect 485118 21218 485160 21454
rect 484840 21134 485160 21218
rect 484840 20898 484882 21134
rect 485118 20898 485160 21134
rect 484840 20866 485160 20898
rect 490771 21454 491091 21486
rect 490771 21218 490813 21454
rect 491049 21218 491091 21454
rect 490771 21134 491091 21218
rect 490771 20898 490813 21134
rect 491049 20898 491091 21134
rect 490771 20866 491091 20898
rect 505910 21454 506230 21486
rect 505910 21218 505952 21454
rect 506188 21218 506230 21454
rect 505910 21134 506230 21218
rect 505910 20898 505952 21134
rect 506188 20898 506230 21134
rect 505910 20866 506230 20898
rect 511840 21454 512160 21486
rect 511840 21218 511882 21454
rect 512118 21218 512160 21454
rect 511840 21134 512160 21218
rect 511840 20898 511882 21134
rect 512118 20898 512160 21134
rect 511840 20866 512160 20898
rect 517771 21454 518091 21486
rect 517771 21218 517813 21454
rect 518049 21218 518091 21454
rect 517771 21134 518091 21218
rect 517771 20898 517813 21134
rect 518049 20898 518091 21134
rect 517771 20866 518091 20898
rect 532910 21454 533230 21486
rect 532910 21218 532952 21454
rect 533188 21218 533230 21454
rect 532910 21134 533230 21218
rect 532910 20898 532952 21134
rect 533188 20898 533230 21134
rect 532910 20866 533230 20898
rect 538840 21454 539160 21486
rect 538840 21218 538882 21454
rect 539118 21218 539160 21454
rect 538840 21134 539160 21218
rect 538840 20898 538882 21134
rect 539118 20898 539160 21134
rect 538840 20866 539160 20898
rect 544771 21454 545091 21486
rect 544771 21218 544813 21454
rect 545049 21218 545091 21454
rect 544771 21134 545091 21218
rect 544771 20898 544813 21134
rect 545049 20898 545091 21134
rect 544771 20866 545091 20898
rect 559794 21454 560414 38898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -1306 11414 11898
rect 10794 -1542 10826 -1306
rect 11062 -1542 11146 -1306
rect 11382 -1542 11414 -1306
rect 10794 -1626 11414 -1542
rect 10794 -1862 10826 -1626
rect 11062 -1862 11146 -1626
rect 11382 -1862 11414 -1626
rect 10794 -1894 11414 -1862
rect 19794 3454 20414 14000
rect 19794 3218 19826 3454
rect 20062 3218 20146 3454
rect 20382 3218 20414 3454
rect 19794 3134 20414 3218
rect 19794 2898 19826 3134
rect 20062 2898 20146 3134
rect 20382 2898 20414 3134
rect 19794 -346 20414 2898
rect 19794 -582 19826 -346
rect 20062 -582 20146 -346
rect 20382 -582 20414 -346
rect 19794 -666 20414 -582
rect 19794 -902 19826 -666
rect 20062 -902 20146 -666
rect 20382 -902 20414 -666
rect 19794 -1894 20414 -902
rect 28794 12454 29414 14000
rect 28794 12218 28826 12454
rect 29062 12218 29146 12454
rect 29382 12218 29414 12454
rect 28794 12134 29414 12218
rect 28794 11898 28826 12134
rect 29062 11898 29146 12134
rect 29382 11898 29414 12134
rect 28794 -1306 29414 11898
rect 28794 -1542 28826 -1306
rect 29062 -1542 29146 -1306
rect 29382 -1542 29414 -1306
rect 28794 -1626 29414 -1542
rect 28794 -1862 28826 -1626
rect 29062 -1862 29146 -1626
rect 29382 -1862 29414 -1626
rect 28794 -1894 29414 -1862
rect 37794 3454 38414 14000
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 46794 12454 47414 14000
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -1306 47414 11898
rect 46794 -1542 46826 -1306
rect 47062 -1542 47146 -1306
rect 47382 -1542 47414 -1306
rect 46794 -1626 47414 -1542
rect 46794 -1862 46826 -1626
rect 47062 -1862 47146 -1626
rect 47382 -1862 47414 -1626
rect 46794 -1894 47414 -1862
rect 55794 3454 56414 14000
rect 55794 3218 55826 3454
rect 56062 3218 56146 3454
rect 56382 3218 56414 3454
rect 55794 3134 56414 3218
rect 55794 2898 55826 3134
rect 56062 2898 56146 3134
rect 56382 2898 56414 3134
rect 55794 -346 56414 2898
rect 55794 -582 55826 -346
rect 56062 -582 56146 -346
rect 56382 -582 56414 -346
rect 55794 -666 56414 -582
rect 55794 -902 55826 -666
rect 56062 -902 56146 -666
rect 56382 -902 56414 -666
rect 55794 -1894 56414 -902
rect 64794 12454 65414 14000
rect 64794 12218 64826 12454
rect 65062 12218 65146 12454
rect 65382 12218 65414 12454
rect 64794 12134 65414 12218
rect 64794 11898 64826 12134
rect 65062 11898 65146 12134
rect 65382 11898 65414 12134
rect 64794 -1306 65414 11898
rect 64794 -1542 64826 -1306
rect 65062 -1542 65146 -1306
rect 65382 -1542 65414 -1306
rect 64794 -1626 65414 -1542
rect 64794 -1862 64826 -1626
rect 65062 -1862 65146 -1626
rect 65382 -1862 65414 -1626
rect 64794 -1894 65414 -1862
rect 73794 3454 74414 14000
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 82794 12454 83414 14000
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -1306 83414 11898
rect 82794 -1542 82826 -1306
rect 83062 -1542 83146 -1306
rect 83382 -1542 83414 -1306
rect 82794 -1626 83414 -1542
rect 82794 -1862 82826 -1626
rect 83062 -1862 83146 -1626
rect 83382 -1862 83414 -1626
rect 82794 -1894 83414 -1862
rect 91794 3454 92414 14000
rect 91794 3218 91826 3454
rect 92062 3218 92146 3454
rect 92382 3218 92414 3454
rect 91794 3134 92414 3218
rect 91794 2898 91826 3134
rect 92062 2898 92146 3134
rect 92382 2898 92414 3134
rect 91794 -346 92414 2898
rect 91794 -582 91826 -346
rect 92062 -582 92146 -346
rect 92382 -582 92414 -346
rect 91794 -666 92414 -582
rect 91794 -902 91826 -666
rect 92062 -902 92146 -666
rect 92382 -902 92414 -666
rect 91794 -1894 92414 -902
rect 100794 12454 101414 14000
rect 100794 12218 100826 12454
rect 101062 12218 101146 12454
rect 101382 12218 101414 12454
rect 100794 12134 101414 12218
rect 100794 11898 100826 12134
rect 101062 11898 101146 12134
rect 101382 11898 101414 12134
rect 100794 -1306 101414 11898
rect 100794 -1542 100826 -1306
rect 101062 -1542 101146 -1306
rect 101382 -1542 101414 -1306
rect 100794 -1626 101414 -1542
rect 100794 -1862 100826 -1626
rect 101062 -1862 101146 -1626
rect 101382 -1862 101414 -1626
rect 100794 -1894 101414 -1862
rect 109794 3454 110414 14000
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 118794 12454 119414 14000
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -1306 119414 11898
rect 118794 -1542 118826 -1306
rect 119062 -1542 119146 -1306
rect 119382 -1542 119414 -1306
rect 118794 -1626 119414 -1542
rect 118794 -1862 118826 -1626
rect 119062 -1862 119146 -1626
rect 119382 -1862 119414 -1626
rect 118794 -1894 119414 -1862
rect 127794 3454 128414 14000
rect 127794 3218 127826 3454
rect 128062 3218 128146 3454
rect 128382 3218 128414 3454
rect 127794 3134 128414 3218
rect 127794 2898 127826 3134
rect 128062 2898 128146 3134
rect 128382 2898 128414 3134
rect 127794 -346 128414 2898
rect 127794 -582 127826 -346
rect 128062 -582 128146 -346
rect 128382 -582 128414 -346
rect 127794 -666 128414 -582
rect 127794 -902 127826 -666
rect 128062 -902 128146 -666
rect 128382 -902 128414 -666
rect 127794 -1894 128414 -902
rect 136794 12454 137414 14000
rect 136794 12218 136826 12454
rect 137062 12218 137146 12454
rect 137382 12218 137414 12454
rect 136794 12134 137414 12218
rect 136794 11898 136826 12134
rect 137062 11898 137146 12134
rect 137382 11898 137414 12134
rect 136794 -1306 137414 11898
rect 136794 -1542 136826 -1306
rect 137062 -1542 137146 -1306
rect 137382 -1542 137414 -1306
rect 136794 -1626 137414 -1542
rect 136794 -1862 136826 -1626
rect 137062 -1862 137146 -1626
rect 137382 -1862 137414 -1626
rect 136794 -1894 137414 -1862
rect 145794 3454 146414 14000
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 154794 12454 155414 14000
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -1306 155414 11898
rect 154794 -1542 154826 -1306
rect 155062 -1542 155146 -1306
rect 155382 -1542 155414 -1306
rect 154794 -1626 155414 -1542
rect 154794 -1862 154826 -1626
rect 155062 -1862 155146 -1626
rect 155382 -1862 155414 -1626
rect 154794 -1894 155414 -1862
rect 163794 3454 164414 14000
rect 163794 3218 163826 3454
rect 164062 3218 164146 3454
rect 164382 3218 164414 3454
rect 163794 3134 164414 3218
rect 163794 2898 163826 3134
rect 164062 2898 164146 3134
rect 164382 2898 164414 3134
rect 163794 -346 164414 2898
rect 163794 -582 163826 -346
rect 164062 -582 164146 -346
rect 164382 -582 164414 -346
rect 163794 -666 164414 -582
rect 163794 -902 163826 -666
rect 164062 -902 164146 -666
rect 164382 -902 164414 -666
rect 163794 -1894 164414 -902
rect 172794 12454 173414 14000
rect 172794 12218 172826 12454
rect 173062 12218 173146 12454
rect 173382 12218 173414 12454
rect 172794 12134 173414 12218
rect 172794 11898 172826 12134
rect 173062 11898 173146 12134
rect 173382 11898 173414 12134
rect 172794 -1306 173414 11898
rect 172794 -1542 172826 -1306
rect 173062 -1542 173146 -1306
rect 173382 -1542 173414 -1306
rect 172794 -1626 173414 -1542
rect 172794 -1862 172826 -1626
rect 173062 -1862 173146 -1626
rect 173382 -1862 173414 -1626
rect 172794 -1894 173414 -1862
rect 181794 3454 182414 14000
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 190794 12454 191414 14000
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -1306 191414 11898
rect 190794 -1542 190826 -1306
rect 191062 -1542 191146 -1306
rect 191382 -1542 191414 -1306
rect 190794 -1626 191414 -1542
rect 190794 -1862 190826 -1626
rect 191062 -1862 191146 -1626
rect 191382 -1862 191414 -1626
rect 190794 -1894 191414 -1862
rect 199794 3454 200414 14000
rect 199794 3218 199826 3454
rect 200062 3218 200146 3454
rect 200382 3218 200414 3454
rect 199794 3134 200414 3218
rect 199794 2898 199826 3134
rect 200062 2898 200146 3134
rect 200382 2898 200414 3134
rect 199794 -346 200414 2898
rect 199794 -582 199826 -346
rect 200062 -582 200146 -346
rect 200382 -582 200414 -346
rect 199794 -666 200414 -582
rect 199794 -902 199826 -666
rect 200062 -902 200146 -666
rect 200382 -902 200414 -666
rect 199794 -1894 200414 -902
rect 208794 12454 209414 14000
rect 208794 12218 208826 12454
rect 209062 12218 209146 12454
rect 209382 12218 209414 12454
rect 208794 12134 209414 12218
rect 208794 11898 208826 12134
rect 209062 11898 209146 12134
rect 209382 11898 209414 12134
rect 208794 -1306 209414 11898
rect 208794 -1542 208826 -1306
rect 209062 -1542 209146 -1306
rect 209382 -1542 209414 -1306
rect 208794 -1626 209414 -1542
rect 208794 -1862 208826 -1626
rect 209062 -1862 209146 -1626
rect 209382 -1862 209414 -1626
rect 208794 -1894 209414 -1862
rect 217794 3454 218414 14000
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 226794 12454 227414 14000
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -1306 227414 11898
rect 226794 -1542 226826 -1306
rect 227062 -1542 227146 -1306
rect 227382 -1542 227414 -1306
rect 226794 -1626 227414 -1542
rect 226794 -1862 226826 -1626
rect 227062 -1862 227146 -1626
rect 227382 -1862 227414 -1626
rect 226794 -1894 227414 -1862
rect 235794 3454 236414 14000
rect 235794 3218 235826 3454
rect 236062 3218 236146 3454
rect 236382 3218 236414 3454
rect 235794 3134 236414 3218
rect 235794 2898 235826 3134
rect 236062 2898 236146 3134
rect 236382 2898 236414 3134
rect 235794 -346 236414 2898
rect 235794 -582 235826 -346
rect 236062 -582 236146 -346
rect 236382 -582 236414 -346
rect 235794 -666 236414 -582
rect 235794 -902 235826 -666
rect 236062 -902 236146 -666
rect 236382 -902 236414 -666
rect 235794 -1894 236414 -902
rect 244794 12454 245414 14000
rect 244794 12218 244826 12454
rect 245062 12218 245146 12454
rect 245382 12218 245414 12454
rect 244794 12134 245414 12218
rect 244794 11898 244826 12134
rect 245062 11898 245146 12134
rect 245382 11898 245414 12134
rect 244794 -1306 245414 11898
rect 244794 -1542 244826 -1306
rect 245062 -1542 245146 -1306
rect 245382 -1542 245414 -1306
rect 244794 -1626 245414 -1542
rect 244794 -1862 244826 -1626
rect 245062 -1862 245146 -1626
rect 245382 -1862 245414 -1626
rect 244794 -1894 245414 -1862
rect 253794 3454 254414 14000
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 262794 12454 263414 14000
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -1306 263414 11898
rect 262794 -1542 262826 -1306
rect 263062 -1542 263146 -1306
rect 263382 -1542 263414 -1306
rect 262794 -1626 263414 -1542
rect 262794 -1862 262826 -1626
rect 263062 -1862 263146 -1626
rect 263382 -1862 263414 -1626
rect 262794 -1894 263414 -1862
rect 271794 3454 272414 14000
rect 271794 3218 271826 3454
rect 272062 3218 272146 3454
rect 272382 3218 272414 3454
rect 271794 3134 272414 3218
rect 271794 2898 271826 3134
rect 272062 2898 272146 3134
rect 272382 2898 272414 3134
rect 271794 -346 272414 2898
rect 271794 -582 271826 -346
rect 272062 -582 272146 -346
rect 272382 -582 272414 -346
rect 271794 -666 272414 -582
rect 271794 -902 271826 -666
rect 272062 -902 272146 -666
rect 272382 -902 272414 -666
rect 271794 -1894 272414 -902
rect 280794 12454 281414 14000
rect 280794 12218 280826 12454
rect 281062 12218 281146 12454
rect 281382 12218 281414 12454
rect 280794 12134 281414 12218
rect 280794 11898 280826 12134
rect 281062 11898 281146 12134
rect 281382 11898 281414 12134
rect 280794 -1306 281414 11898
rect 280794 -1542 280826 -1306
rect 281062 -1542 281146 -1306
rect 281382 -1542 281414 -1306
rect 280794 -1626 281414 -1542
rect 280794 -1862 280826 -1626
rect 281062 -1862 281146 -1626
rect 281382 -1862 281414 -1626
rect 280794 -1894 281414 -1862
rect 289794 3454 290414 14000
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 298794 12454 299414 14000
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -1306 299414 11898
rect 298794 -1542 298826 -1306
rect 299062 -1542 299146 -1306
rect 299382 -1542 299414 -1306
rect 298794 -1626 299414 -1542
rect 298794 -1862 298826 -1626
rect 299062 -1862 299146 -1626
rect 299382 -1862 299414 -1626
rect 298794 -1894 299414 -1862
rect 307794 3454 308414 14000
rect 307794 3218 307826 3454
rect 308062 3218 308146 3454
rect 308382 3218 308414 3454
rect 307794 3134 308414 3218
rect 307794 2898 307826 3134
rect 308062 2898 308146 3134
rect 308382 2898 308414 3134
rect 307794 -346 308414 2898
rect 307794 -582 307826 -346
rect 308062 -582 308146 -346
rect 308382 -582 308414 -346
rect 307794 -666 308414 -582
rect 307794 -902 307826 -666
rect 308062 -902 308146 -666
rect 308382 -902 308414 -666
rect 307794 -1894 308414 -902
rect 316794 12454 317414 14000
rect 316794 12218 316826 12454
rect 317062 12218 317146 12454
rect 317382 12218 317414 12454
rect 316794 12134 317414 12218
rect 316794 11898 316826 12134
rect 317062 11898 317146 12134
rect 317382 11898 317414 12134
rect 316794 -1306 317414 11898
rect 316794 -1542 316826 -1306
rect 317062 -1542 317146 -1306
rect 317382 -1542 317414 -1306
rect 316794 -1626 317414 -1542
rect 316794 -1862 316826 -1626
rect 317062 -1862 317146 -1626
rect 317382 -1862 317414 -1626
rect 316794 -1894 317414 -1862
rect 325794 3454 326414 14000
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 334794 12454 335414 14000
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -1306 335414 11898
rect 334794 -1542 334826 -1306
rect 335062 -1542 335146 -1306
rect 335382 -1542 335414 -1306
rect 334794 -1626 335414 -1542
rect 334794 -1862 334826 -1626
rect 335062 -1862 335146 -1626
rect 335382 -1862 335414 -1626
rect 334794 -1894 335414 -1862
rect 343794 3454 344414 14000
rect 343794 3218 343826 3454
rect 344062 3218 344146 3454
rect 344382 3218 344414 3454
rect 343794 3134 344414 3218
rect 343794 2898 343826 3134
rect 344062 2898 344146 3134
rect 344382 2898 344414 3134
rect 343794 -346 344414 2898
rect 343794 -582 343826 -346
rect 344062 -582 344146 -346
rect 344382 -582 344414 -346
rect 343794 -666 344414 -582
rect 343794 -902 343826 -666
rect 344062 -902 344146 -666
rect 344382 -902 344414 -666
rect 343794 -1894 344414 -902
rect 352794 12454 353414 14000
rect 352794 12218 352826 12454
rect 353062 12218 353146 12454
rect 353382 12218 353414 12454
rect 352794 12134 353414 12218
rect 352794 11898 352826 12134
rect 353062 11898 353146 12134
rect 353382 11898 353414 12134
rect 352794 -1306 353414 11898
rect 352794 -1542 352826 -1306
rect 353062 -1542 353146 -1306
rect 353382 -1542 353414 -1306
rect 352794 -1626 353414 -1542
rect 352794 -1862 352826 -1626
rect 353062 -1862 353146 -1626
rect 353382 -1862 353414 -1626
rect 352794 -1894 353414 -1862
rect 361794 3454 362414 14000
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 370794 12454 371414 14000
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -1306 371414 11898
rect 370794 -1542 370826 -1306
rect 371062 -1542 371146 -1306
rect 371382 -1542 371414 -1306
rect 370794 -1626 371414 -1542
rect 370794 -1862 370826 -1626
rect 371062 -1862 371146 -1626
rect 371382 -1862 371414 -1626
rect 370794 -1894 371414 -1862
rect 379794 3454 380414 14000
rect 379794 3218 379826 3454
rect 380062 3218 380146 3454
rect 380382 3218 380414 3454
rect 379794 3134 380414 3218
rect 379794 2898 379826 3134
rect 380062 2898 380146 3134
rect 380382 2898 380414 3134
rect 379794 -346 380414 2898
rect 379794 -582 379826 -346
rect 380062 -582 380146 -346
rect 380382 -582 380414 -346
rect 379794 -666 380414 -582
rect 379794 -902 379826 -666
rect 380062 -902 380146 -666
rect 380382 -902 380414 -666
rect 379794 -1894 380414 -902
rect 388794 12454 389414 14000
rect 388794 12218 388826 12454
rect 389062 12218 389146 12454
rect 389382 12218 389414 12454
rect 388794 12134 389414 12218
rect 388794 11898 388826 12134
rect 389062 11898 389146 12134
rect 389382 11898 389414 12134
rect 388794 -1306 389414 11898
rect 388794 -1542 388826 -1306
rect 389062 -1542 389146 -1306
rect 389382 -1542 389414 -1306
rect 388794 -1626 389414 -1542
rect 388794 -1862 388826 -1626
rect 389062 -1862 389146 -1626
rect 389382 -1862 389414 -1626
rect 388794 -1894 389414 -1862
rect 397794 3454 398414 14000
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 406794 12454 407414 14000
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -1306 407414 11898
rect 406794 -1542 406826 -1306
rect 407062 -1542 407146 -1306
rect 407382 -1542 407414 -1306
rect 406794 -1626 407414 -1542
rect 406794 -1862 406826 -1626
rect 407062 -1862 407146 -1626
rect 407382 -1862 407414 -1626
rect 406794 -1894 407414 -1862
rect 415794 3454 416414 14000
rect 415794 3218 415826 3454
rect 416062 3218 416146 3454
rect 416382 3218 416414 3454
rect 415794 3134 416414 3218
rect 415794 2898 415826 3134
rect 416062 2898 416146 3134
rect 416382 2898 416414 3134
rect 415794 -346 416414 2898
rect 415794 -582 415826 -346
rect 416062 -582 416146 -346
rect 416382 -582 416414 -346
rect 415794 -666 416414 -582
rect 415794 -902 415826 -666
rect 416062 -902 416146 -666
rect 416382 -902 416414 -666
rect 415794 -1894 416414 -902
rect 424794 12454 425414 14000
rect 424794 12218 424826 12454
rect 425062 12218 425146 12454
rect 425382 12218 425414 12454
rect 424794 12134 425414 12218
rect 424794 11898 424826 12134
rect 425062 11898 425146 12134
rect 425382 11898 425414 12134
rect 424794 -1306 425414 11898
rect 424794 -1542 424826 -1306
rect 425062 -1542 425146 -1306
rect 425382 -1542 425414 -1306
rect 424794 -1626 425414 -1542
rect 424794 -1862 424826 -1626
rect 425062 -1862 425146 -1626
rect 425382 -1862 425414 -1626
rect 424794 -1894 425414 -1862
rect 433794 3454 434414 14000
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 442794 12454 443414 14000
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -1306 443414 11898
rect 442794 -1542 442826 -1306
rect 443062 -1542 443146 -1306
rect 443382 -1542 443414 -1306
rect 442794 -1626 443414 -1542
rect 442794 -1862 442826 -1626
rect 443062 -1862 443146 -1626
rect 443382 -1862 443414 -1626
rect 442794 -1894 443414 -1862
rect 451794 3454 452414 14000
rect 451794 3218 451826 3454
rect 452062 3218 452146 3454
rect 452382 3218 452414 3454
rect 451794 3134 452414 3218
rect 451794 2898 451826 3134
rect 452062 2898 452146 3134
rect 452382 2898 452414 3134
rect 451794 -346 452414 2898
rect 451794 -582 451826 -346
rect 452062 -582 452146 -346
rect 452382 -582 452414 -346
rect 451794 -666 452414 -582
rect 451794 -902 451826 -666
rect 452062 -902 452146 -666
rect 452382 -902 452414 -666
rect 451794 -1894 452414 -902
rect 460794 12454 461414 14000
rect 460794 12218 460826 12454
rect 461062 12218 461146 12454
rect 461382 12218 461414 12454
rect 460794 12134 461414 12218
rect 460794 11898 460826 12134
rect 461062 11898 461146 12134
rect 461382 11898 461414 12134
rect 460794 -1306 461414 11898
rect 460794 -1542 460826 -1306
rect 461062 -1542 461146 -1306
rect 461382 -1542 461414 -1306
rect 460794 -1626 461414 -1542
rect 460794 -1862 460826 -1626
rect 461062 -1862 461146 -1626
rect 461382 -1862 461414 -1626
rect 460794 -1894 461414 -1862
rect 469794 3454 470414 14000
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 478794 12454 479414 14000
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -1306 479414 11898
rect 478794 -1542 478826 -1306
rect 479062 -1542 479146 -1306
rect 479382 -1542 479414 -1306
rect 478794 -1626 479414 -1542
rect 478794 -1862 478826 -1626
rect 479062 -1862 479146 -1626
rect 479382 -1862 479414 -1626
rect 478794 -1894 479414 -1862
rect 487794 3454 488414 14000
rect 487794 3218 487826 3454
rect 488062 3218 488146 3454
rect 488382 3218 488414 3454
rect 487794 3134 488414 3218
rect 487794 2898 487826 3134
rect 488062 2898 488146 3134
rect 488382 2898 488414 3134
rect 487794 -346 488414 2898
rect 487794 -582 487826 -346
rect 488062 -582 488146 -346
rect 488382 -582 488414 -346
rect 487794 -666 488414 -582
rect 487794 -902 487826 -666
rect 488062 -902 488146 -666
rect 488382 -902 488414 -666
rect 487794 -1894 488414 -902
rect 496794 12454 497414 14000
rect 496794 12218 496826 12454
rect 497062 12218 497146 12454
rect 497382 12218 497414 12454
rect 496794 12134 497414 12218
rect 496794 11898 496826 12134
rect 497062 11898 497146 12134
rect 497382 11898 497414 12134
rect 496794 -1306 497414 11898
rect 496794 -1542 496826 -1306
rect 497062 -1542 497146 -1306
rect 497382 -1542 497414 -1306
rect 496794 -1626 497414 -1542
rect 496794 -1862 496826 -1626
rect 497062 -1862 497146 -1626
rect 497382 -1862 497414 -1626
rect 496794 -1894 497414 -1862
rect 505794 3454 506414 14000
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 514794 12454 515414 14000
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -1306 515414 11898
rect 514794 -1542 514826 -1306
rect 515062 -1542 515146 -1306
rect 515382 -1542 515414 -1306
rect 514794 -1626 515414 -1542
rect 514794 -1862 514826 -1626
rect 515062 -1862 515146 -1626
rect 515382 -1862 515414 -1626
rect 514794 -1894 515414 -1862
rect 523794 3454 524414 14000
rect 523794 3218 523826 3454
rect 524062 3218 524146 3454
rect 524382 3218 524414 3454
rect 523794 3134 524414 3218
rect 523794 2898 523826 3134
rect 524062 2898 524146 3134
rect 524382 2898 524414 3134
rect 523794 -346 524414 2898
rect 523794 -582 523826 -346
rect 524062 -582 524146 -346
rect 524382 -582 524414 -346
rect 523794 -666 524414 -582
rect 523794 -902 523826 -666
rect 524062 -902 524146 -666
rect 524382 -902 524414 -666
rect 523794 -1894 524414 -902
rect 532794 12454 533414 14000
rect 532794 12218 532826 12454
rect 533062 12218 533146 12454
rect 533382 12218 533414 12454
rect 532794 12134 533414 12218
rect 532794 11898 532826 12134
rect 533062 11898 533146 12134
rect 533382 11898 533414 12134
rect 532794 -1306 533414 11898
rect 532794 -1542 532826 -1306
rect 533062 -1542 533146 -1306
rect 533382 -1542 533414 -1306
rect 532794 -1626 533414 -1542
rect 532794 -1862 532826 -1626
rect 533062 -1862 533146 -1626
rect 533382 -1862 533414 -1626
rect 532794 -1894 533414 -1862
rect 541794 3454 542414 14000
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 550794 12454 551414 14000
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -1306 551414 11898
rect 550794 -1542 550826 -1306
rect 551062 -1542 551146 -1306
rect 551382 -1542 551414 -1306
rect 550794 -1626 551414 -1542
rect 550794 -1862 550826 -1626
rect 551062 -1862 551146 -1626
rect 551382 -1862 551414 -1626
rect 550794 -1894 551414 -1862
rect 559794 3454 560414 20898
rect 559794 3218 559826 3454
rect 560062 3218 560146 3454
rect 560382 3218 560414 3454
rect 559794 3134 560414 3218
rect 559794 2898 559826 3134
rect 560062 2898 560146 3134
rect 560382 2898 560414 3134
rect 559794 -346 560414 2898
rect 559794 -582 559826 -346
rect 560062 -582 560146 -346
rect 560382 -582 560414 -346
rect 559794 -666 560414 -582
rect 559794 -902 559826 -666
rect 560062 -902 560146 -666
rect 560382 -902 560414 -666
rect 559794 -1894 560414 -902
rect 568794 705798 569414 705830
rect 568794 705562 568826 705798
rect 569062 705562 569146 705798
rect 569382 705562 569414 705798
rect 568794 705478 569414 705562
rect 568794 705242 568826 705478
rect 569062 705242 569146 705478
rect 569382 705242 569414 705478
rect 568794 696454 569414 705242
rect 568794 696218 568826 696454
rect 569062 696218 569146 696454
rect 569382 696218 569414 696454
rect 568794 696134 569414 696218
rect 568794 695898 568826 696134
rect 569062 695898 569146 696134
rect 569382 695898 569414 696134
rect 568794 678454 569414 695898
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 660454 569414 677898
rect 568794 660218 568826 660454
rect 569062 660218 569146 660454
rect 569382 660218 569414 660454
rect 568794 660134 569414 660218
rect 568794 659898 568826 660134
rect 569062 659898 569146 660134
rect 569382 659898 569414 660134
rect 568794 642454 569414 659898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 624454 569414 641898
rect 568794 624218 568826 624454
rect 569062 624218 569146 624454
rect 569382 624218 569414 624454
rect 568794 624134 569414 624218
rect 568794 623898 568826 624134
rect 569062 623898 569146 624134
rect 569382 623898 569414 624134
rect 568794 606454 569414 623898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 588454 569414 605898
rect 568794 588218 568826 588454
rect 569062 588218 569146 588454
rect 569382 588218 569414 588454
rect 568794 588134 569414 588218
rect 568794 587898 568826 588134
rect 569062 587898 569146 588134
rect 569382 587898 569414 588134
rect 568794 570454 569414 587898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 552454 569414 569898
rect 568794 552218 568826 552454
rect 569062 552218 569146 552454
rect 569382 552218 569414 552454
rect 568794 552134 569414 552218
rect 568794 551898 568826 552134
rect 569062 551898 569146 552134
rect 569382 551898 569414 552134
rect 568794 534454 569414 551898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 516454 569414 533898
rect 568794 516218 568826 516454
rect 569062 516218 569146 516454
rect 569382 516218 569414 516454
rect 568794 516134 569414 516218
rect 568794 515898 568826 516134
rect 569062 515898 569146 516134
rect 569382 515898 569414 516134
rect 568794 498454 569414 515898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 480454 569414 497898
rect 568794 480218 568826 480454
rect 569062 480218 569146 480454
rect 569382 480218 569414 480454
rect 568794 480134 569414 480218
rect 568794 479898 568826 480134
rect 569062 479898 569146 480134
rect 569382 479898 569414 480134
rect 568794 462454 569414 479898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 444454 569414 461898
rect 568794 444218 568826 444454
rect 569062 444218 569146 444454
rect 569382 444218 569414 444454
rect 568794 444134 569414 444218
rect 568794 443898 568826 444134
rect 569062 443898 569146 444134
rect 569382 443898 569414 444134
rect 568794 426454 569414 443898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 408454 569414 425898
rect 568794 408218 568826 408454
rect 569062 408218 569146 408454
rect 569382 408218 569414 408454
rect 568794 408134 569414 408218
rect 568794 407898 568826 408134
rect 569062 407898 569146 408134
rect 569382 407898 569414 408134
rect 568794 390454 569414 407898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 372454 569414 389898
rect 568794 372218 568826 372454
rect 569062 372218 569146 372454
rect 569382 372218 569414 372454
rect 568794 372134 569414 372218
rect 568794 371898 568826 372134
rect 569062 371898 569146 372134
rect 569382 371898 569414 372134
rect 568794 354454 569414 371898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 336454 569414 353898
rect 568794 336218 568826 336454
rect 569062 336218 569146 336454
rect 569382 336218 569414 336454
rect 568794 336134 569414 336218
rect 568794 335898 568826 336134
rect 569062 335898 569146 336134
rect 569382 335898 569414 336134
rect 568794 318454 569414 335898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 300454 569414 317898
rect 568794 300218 568826 300454
rect 569062 300218 569146 300454
rect 569382 300218 569414 300454
rect 568794 300134 569414 300218
rect 568794 299898 568826 300134
rect 569062 299898 569146 300134
rect 569382 299898 569414 300134
rect 568794 282454 569414 299898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 264454 569414 281898
rect 568794 264218 568826 264454
rect 569062 264218 569146 264454
rect 569382 264218 569414 264454
rect 568794 264134 569414 264218
rect 568794 263898 568826 264134
rect 569062 263898 569146 264134
rect 569382 263898 569414 264134
rect 568794 246454 569414 263898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 228454 569414 245898
rect 568794 228218 568826 228454
rect 569062 228218 569146 228454
rect 569382 228218 569414 228454
rect 568794 228134 569414 228218
rect 568794 227898 568826 228134
rect 569062 227898 569146 228134
rect 569382 227898 569414 228134
rect 568794 210454 569414 227898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 192454 569414 209898
rect 568794 192218 568826 192454
rect 569062 192218 569146 192454
rect 569382 192218 569414 192454
rect 568794 192134 569414 192218
rect 568794 191898 568826 192134
rect 569062 191898 569146 192134
rect 569382 191898 569414 192134
rect 568794 174454 569414 191898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 156454 569414 173898
rect 568794 156218 568826 156454
rect 569062 156218 569146 156454
rect 569382 156218 569414 156454
rect 568794 156134 569414 156218
rect 568794 155898 568826 156134
rect 569062 155898 569146 156134
rect 569382 155898 569414 156134
rect 568794 138454 569414 155898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 120454 569414 137898
rect 568794 120218 568826 120454
rect 569062 120218 569146 120454
rect 569382 120218 569414 120454
rect 568794 120134 569414 120218
rect 568794 119898 568826 120134
rect 569062 119898 569146 120134
rect 569382 119898 569414 120134
rect 568794 102454 569414 119898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 84454 569414 101898
rect 568794 84218 568826 84454
rect 569062 84218 569146 84454
rect 569382 84218 569414 84454
rect 568794 84134 569414 84218
rect 568794 83898 568826 84134
rect 569062 83898 569146 84134
rect 569382 83898 569414 84134
rect 568794 66454 569414 83898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 48454 569414 65898
rect 568794 48218 568826 48454
rect 569062 48218 569146 48454
rect 569382 48218 569414 48454
rect 568794 48134 569414 48218
rect 568794 47898 568826 48134
rect 569062 47898 569146 48134
rect 569382 47898 569414 48134
rect 568794 30454 569414 47898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 12454 569414 29898
rect 568794 12218 568826 12454
rect 569062 12218 569146 12454
rect 569382 12218 569414 12454
rect 568794 12134 569414 12218
rect 568794 11898 568826 12134
rect 569062 11898 569146 12134
rect 569382 11898 569414 12134
rect 568794 -1306 569414 11898
rect 568794 -1542 568826 -1306
rect 569062 -1542 569146 -1306
rect 569382 -1542 569414 -1306
rect 568794 -1626 569414 -1542
rect 568794 -1862 568826 -1626
rect 569062 -1862 569146 -1626
rect 569382 -1862 569414 -1626
rect 568794 -1894 569414 -1862
rect 577794 704838 578414 705830
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 669454 578414 686898
rect 577794 669218 577826 669454
rect 578062 669218 578146 669454
rect 578382 669218 578414 669454
rect 577794 669134 578414 669218
rect 577794 668898 577826 669134
rect 578062 668898 578146 669134
rect 578382 668898 578414 669134
rect 577794 651454 578414 668898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 633454 578414 650898
rect 577794 633218 577826 633454
rect 578062 633218 578146 633454
rect 578382 633218 578414 633454
rect 577794 633134 578414 633218
rect 577794 632898 577826 633134
rect 578062 632898 578146 633134
rect 578382 632898 578414 633134
rect 577794 615454 578414 632898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 597454 578414 614898
rect 577794 597218 577826 597454
rect 578062 597218 578146 597454
rect 578382 597218 578414 597454
rect 577794 597134 578414 597218
rect 577794 596898 577826 597134
rect 578062 596898 578146 597134
rect 578382 596898 578414 597134
rect 577794 579454 578414 596898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 561454 578414 578898
rect 577794 561218 577826 561454
rect 578062 561218 578146 561454
rect 578382 561218 578414 561454
rect 577794 561134 578414 561218
rect 577794 560898 577826 561134
rect 578062 560898 578146 561134
rect 578382 560898 578414 561134
rect 577794 543454 578414 560898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 525454 578414 542898
rect 577794 525218 577826 525454
rect 578062 525218 578146 525454
rect 578382 525218 578414 525454
rect 577794 525134 578414 525218
rect 577794 524898 577826 525134
rect 578062 524898 578146 525134
rect 578382 524898 578414 525134
rect 577794 507454 578414 524898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 489454 578414 506898
rect 577794 489218 577826 489454
rect 578062 489218 578146 489454
rect 578382 489218 578414 489454
rect 577794 489134 578414 489218
rect 577794 488898 577826 489134
rect 578062 488898 578146 489134
rect 578382 488898 578414 489134
rect 577794 471454 578414 488898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 453454 578414 470898
rect 577794 453218 577826 453454
rect 578062 453218 578146 453454
rect 578382 453218 578414 453454
rect 577794 453134 578414 453218
rect 577794 452898 577826 453134
rect 578062 452898 578146 453134
rect 578382 452898 578414 453134
rect 577794 435454 578414 452898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 417454 578414 434898
rect 577794 417218 577826 417454
rect 578062 417218 578146 417454
rect 578382 417218 578414 417454
rect 577794 417134 578414 417218
rect 577794 416898 577826 417134
rect 578062 416898 578146 417134
rect 578382 416898 578414 417134
rect 577794 399454 578414 416898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 381454 578414 398898
rect 577794 381218 577826 381454
rect 578062 381218 578146 381454
rect 578382 381218 578414 381454
rect 577794 381134 578414 381218
rect 577794 380898 577826 381134
rect 578062 380898 578146 381134
rect 578382 380898 578414 381134
rect 577794 363454 578414 380898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 345454 578414 362898
rect 577794 345218 577826 345454
rect 578062 345218 578146 345454
rect 578382 345218 578414 345454
rect 577794 345134 578414 345218
rect 577794 344898 577826 345134
rect 578062 344898 578146 345134
rect 578382 344898 578414 345134
rect 577794 327454 578414 344898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 309454 578414 326898
rect 577794 309218 577826 309454
rect 578062 309218 578146 309454
rect 578382 309218 578414 309454
rect 577794 309134 578414 309218
rect 577794 308898 577826 309134
rect 578062 308898 578146 309134
rect 578382 308898 578414 309134
rect 577794 291454 578414 308898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 273454 578414 290898
rect 577794 273218 577826 273454
rect 578062 273218 578146 273454
rect 578382 273218 578414 273454
rect 577794 273134 578414 273218
rect 577794 272898 577826 273134
rect 578062 272898 578146 273134
rect 578382 272898 578414 273134
rect 577794 255454 578414 272898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 237454 578414 254898
rect 577794 237218 577826 237454
rect 578062 237218 578146 237454
rect 578382 237218 578414 237454
rect 577794 237134 578414 237218
rect 577794 236898 577826 237134
rect 578062 236898 578146 237134
rect 578382 236898 578414 237134
rect 577794 219454 578414 236898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 201454 578414 218898
rect 577794 201218 577826 201454
rect 578062 201218 578146 201454
rect 578382 201218 578414 201454
rect 577794 201134 578414 201218
rect 577794 200898 577826 201134
rect 578062 200898 578146 201134
rect 578382 200898 578414 201134
rect 577794 183454 578414 200898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 165454 578414 182898
rect 577794 165218 577826 165454
rect 578062 165218 578146 165454
rect 578382 165218 578414 165454
rect 577794 165134 578414 165218
rect 577794 164898 577826 165134
rect 578062 164898 578146 165134
rect 578382 164898 578414 165134
rect 577794 147454 578414 164898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 129454 578414 146898
rect 577794 129218 577826 129454
rect 578062 129218 578146 129454
rect 578382 129218 578414 129454
rect 577794 129134 578414 129218
rect 577794 128898 577826 129134
rect 578062 128898 578146 129134
rect 578382 128898 578414 129134
rect 577794 111454 578414 128898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 93454 578414 110898
rect 577794 93218 577826 93454
rect 578062 93218 578146 93454
rect 578382 93218 578414 93454
rect 577794 93134 578414 93218
rect 577794 92898 577826 93134
rect 578062 92898 578146 93134
rect 578382 92898 578414 93134
rect 577794 75454 578414 92898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 57454 578414 74898
rect 577794 57218 577826 57454
rect 578062 57218 578146 57454
rect 578382 57218 578414 57454
rect 577794 57134 578414 57218
rect 577794 56898 577826 57134
rect 578062 56898 578146 57134
rect 578382 56898 578414 57134
rect 577794 39454 578414 56898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 21454 578414 38898
rect 577794 21218 577826 21454
rect 578062 21218 578146 21454
rect 578382 21218 578414 21454
rect 577794 21134 578414 21218
rect 577794 20898 577826 21134
rect 578062 20898 578146 21134
rect 578382 20898 578414 21134
rect 577794 3454 578414 20898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 669454 585930 686898
rect 585310 669218 585342 669454
rect 585578 669218 585662 669454
rect 585898 669218 585930 669454
rect 585310 669134 585930 669218
rect 585310 668898 585342 669134
rect 585578 668898 585662 669134
rect 585898 668898 585930 669134
rect 585310 651454 585930 668898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 633454 585930 650898
rect 585310 633218 585342 633454
rect 585578 633218 585662 633454
rect 585898 633218 585930 633454
rect 585310 633134 585930 633218
rect 585310 632898 585342 633134
rect 585578 632898 585662 633134
rect 585898 632898 585930 633134
rect 585310 615454 585930 632898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 597454 585930 614898
rect 585310 597218 585342 597454
rect 585578 597218 585662 597454
rect 585898 597218 585930 597454
rect 585310 597134 585930 597218
rect 585310 596898 585342 597134
rect 585578 596898 585662 597134
rect 585898 596898 585930 597134
rect 585310 579454 585930 596898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 561454 585930 578898
rect 585310 561218 585342 561454
rect 585578 561218 585662 561454
rect 585898 561218 585930 561454
rect 585310 561134 585930 561218
rect 585310 560898 585342 561134
rect 585578 560898 585662 561134
rect 585898 560898 585930 561134
rect 585310 543454 585930 560898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 525454 585930 542898
rect 585310 525218 585342 525454
rect 585578 525218 585662 525454
rect 585898 525218 585930 525454
rect 585310 525134 585930 525218
rect 585310 524898 585342 525134
rect 585578 524898 585662 525134
rect 585898 524898 585930 525134
rect 585310 507454 585930 524898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 489454 585930 506898
rect 585310 489218 585342 489454
rect 585578 489218 585662 489454
rect 585898 489218 585930 489454
rect 585310 489134 585930 489218
rect 585310 488898 585342 489134
rect 585578 488898 585662 489134
rect 585898 488898 585930 489134
rect 585310 471454 585930 488898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 453454 585930 470898
rect 585310 453218 585342 453454
rect 585578 453218 585662 453454
rect 585898 453218 585930 453454
rect 585310 453134 585930 453218
rect 585310 452898 585342 453134
rect 585578 452898 585662 453134
rect 585898 452898 585930 453134
rect 585310 435454 585930 452898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 417454 585930 434898
rect 585310 417218 585342 417454
rect 585578 417218 585662 417454
rect 585898 417218 585930 417454
rect 585310 417134 585930 417218
rect 585310 416898 585342 417134
rect 585578 416898 585662 417134
rect 585898 416898 585930 417134
rect 585310 399454 585930 416898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 381454 585930 398898
rect 585310 381218 585342 381454
rect 585578 381218 585662 381454
rect 585898 381218 585930 381454
rect 585310 381134 585930 381218
rect 585310 380898 585342 381134
rect 585578 380898 585662 381134
rect 585898 380898 585930 381134
rect 585310 363454 585930 380898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 345454 585930 362898
rect 585310 345218 585342 345454
rect 585578 345218 585662 345454
rect 585898 345218 585930 345454
rect 585310 345134 585930 345218
rect 585310 344898 585342 345134
rect 585578 344898 585662 345134
rect 585898 344898 585930 345134
rect 585310 327454 585930 344898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 309454 585930 326898
rect 585310 309218 585342 309454
rect 585578 309218 585662 309454
rect 585898 309218 585930 309454
rect 585310 309134 585930 309218
rect 585310 308898 585342 309134
rect 585578 308898 585662 309134
rect 585898 308898 585930 309134
rect 585310 291454 585930 308898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 273454 585930 290898
rect 585310 273218 585342 273454
rect 585578 273218 585662 273454
rect 585898 273218 585930 273454
rect 585310 273134 585930 273218
rect 585310 272898 585342 273134
rect 585578 272898 585662 273134
rect 585898 272898 585930 273134
rect 585310 255454 585930 272898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 237454 585930 254898
rect 585310 237218 585342 237454
rect 585578 237218 585662 237454
rect 585898 237218 585930 237454
rect 585310 237134 585930 237218
rect 585310 236898 585342 237134
rect 585578 236898 585662 237134
rect 585898 236898 585930 237134
rect 585310 219454 585930 236898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 201454 585930 218898
rect 585310 201218 585342 201454
rect 585578 201218 585662 201454
rect 585898 201218 585930 201454
rect 585310 201134 585930 201218
rect 585310 200898 585342 201134
rect 585578 200898 585662 201134
rect 585898 200898 585930 201134
rect 585310 183454 585930 200898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 165454 585930 182898
rect 585310 165218 585342 165454
rect 585578 165218 585662 165454
rect 585898 165218 585930 165454
rect 585310 165134 585930 165218
rect 585310 164898 585342 165134
rect 585578 164898 585662 165134
rect 585898 164898 585930 165134
rect 585310 147454 585930 164898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 129454 585930 146898
rect 585310 129218 585342 129454
rect 585578 129218 585662 129454
rect 585898 129218 585930 129454
rect 585310 129134 585930 129218
rect 585310 128898 585342 129134
rect 585578 128898 585662 129134
rect 585898 128898 585930 129134
rect 585310 111454 585930 128898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 93454 585930 110898
rect 585310 93218 585342 93454
rect 585578 93218 585662 93454
rect 585898 93218 585930 93454
rect 585310 93134 585930 93218
rect 585310 92898 585342 93134
rect 585578 92898 585662 93134
rect 585898 92898 585930 93134
rect 585310 75454 585930 92898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 57454 585930 74898
rect 585310 57218 585342 57454
rect 585578 57218 585662 57454
rect 585898 57218 585930 57454
rect 585310 57134 585930 57218
rect 585310 56898 585342 57134
rect 585578 56898 585662 57134
rect 585898 56898 585930 57134
rect 585310 39454 585930 56898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 21454 585930 38898
rect 585310 21218 585342 21454
rect 585578 21218 585662 21454
rect 585898 21218 585930 21454
rect 585310 21134 585930 21218
rect 585310 20898 585342 21134
rect 585578 20898 585662 21134
rect 585898 20898 585930 21134
rect 585310 3454 585930 20898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 696454 586890 705242
rect 586270 696218 586302 696454
rect 586538 696218 586622 696454
rect 586858 696218 586890 696454
rect 586270 696134 586890 696218
rect 586270 695898 586302 696134
rect 586538 695898 586622 696134
rect 586858 695898 586890 696134
rect 586270 678454 586890 695898
rect 586270 678218 586302 678454
rect 586538 678218 586622 678454
rect 586858 678218 586890 678454
rect 586270 678134 586890 678218
rect 586270 677898 586302 678134
rect 586538 677898 586622 678134
rect 586858 677898 586890 678134
rect 586270 660454 586890 677898
rect 586270 660218 586302 660454
rect 586538 660218 586622 660454
rect 586858 660218 586890 660454
rect 586270 660134 586890 660218
rect 586270 659898 586302 660134
rect 586538 659898 586622 660134
rect 586858 659898 586890 660134
rect 586270 642454 586890 659898
rect 586270 642218 586302 642454
rect 586538 642218 586622 642454
rect 586858 642218 586890 642454
rect 586270 642134 586890 642218
rect 586270 641898 586302 642134
rect 586538 641898 586622 642134
rect 586858 641898 586890 642134
rect 586270 624454 586890 641898
rect 586270 624218 586302 624454
rect 586538 624218 586622 624454
rect 586858 624218 586890 624454
rect 586270 624134 586890 624218
rect 586270 623898 586302 624134
rect 586538 623898 586622 624134
rect 586858 623898 586890 624134
rect 586270 606454 586890 623898
rect 586270 606218 586302 606454
rect 586538 606218 586622 606454
rect 586858 606218 586890 606454
rect 586270 606134 586890 606218
rect 586270 605898 586302 606134
rect 586538 605898 586622 606134
rect 586858 605898 586890 606134
rect 586270 588454 586890 605898
rect 586270 588218 586302 588454
rect 586538 588218 586622 588454
rect 586858 588218 586890 588454
rect 586270 588134 586890 588218
rect 586270 587898 586302 588134
rect 586538 587898 586622 588134
rect 586858 587898 586890 588134
rect 586270 570454 586890 587898
rect 586270 570218 586302 570454
rect 586538 570218 586622 570454
rect 586858 570218 586890 570454
rect 586270 570134 586890 570218
rect 586270 569898 586302 570134
rect 586538 569898 586622 570134
rect 586858 569898 586890 570134
rect 586270 552454 586890 569898
rect 586270 552218 586302 552454
rect 586538 552218 586622 552454
rect 586858 552218 586890 552454
rect 586270 552134 586890 552218
rect 586270 551898 586302 552134
rect 586538 551898 586622 552134
rect 586858 551898 586890 552134
rect 586270 534454 586890 551898
rect 586270 534218 586302 534454
rect 586538 534218 586622 534454
rect 586858 534218 586890 534454
rect 586270 534134 586890 534218
rect 586270 533898 586302 534134
rect 586538 533898 586622 534134
rect 586858 533898 586890 534134
rect 586270 516454 586890 533898
rect 586270 516218 586302 516454
rect 586538 516218 586622 516454
rect 586858 516218 586890 516454
rect 586270 516134 586890 516218
rect 586270 515898 586302 516134
rect 586538 515898 586622 516134
rect 586858 515898 586890 516134
rect 586270 498454 586890 515898
rect 586270 498218 586302 498454
rect 586538 498218 586622 498454
rect 586858 498218 586890 498454
rect 586270 498134 586890 498218
rect 586270 497898 586302 498134
rect 586538 497898 586622 498134
rect 586858 497898 586890 498134
rect 586270 480454 586890 497898
rect 586270 480218 586302 480454
rect 586538 480218 586622 480454
rect 586858 480218 586890 480454
rect 586270 480134 586890 480218
rect 586270 479898 586302 480134
rect 586538 479898 586622 480134
rect 586858 479898 586890 480134
rect 586270 462454 586890 479898
rect 586270 462218 586302 462454
rect 586538 462218 586622 462454
rect 586858 462218 586890 462454
rect 586270 462134 586890 462218
rect 586270 461898 586302 462134
rect 586538 461898 586622 462134
rect 586858 461898 586890 462134
rect 586270 444454 586890 461898
rect 586270 444218 586302 444454
rect 586538 444218 586622 444454
rect 586858 444218 586890 444454
rect 586270 444134 586890 444218
rect 586270 443898 586302 444134
rect 586538 443898 586622 444134
rect 586858 443898 586890 444134
rect 586270 426454 586890 443898
rect 586270 426218 586302 426454
rect 586538 426218 586622 426454
rect 586858 426218 586890 426454
rect 586270 426134 586890 426218
rect 586270 425898 586302 426134
rect 586538 425898 586622 426134
rect 586858 425898 586890 426134
rect 586270 408454 586890 425898
rect 586270 408218 586302 408454
rect 586538 408218 586622 408454
rect 586858 408218 586890 408454
rect 586270 408134 586890 408218
rect 586270 407898 586302 408134
rect 586538 407898 586622 408134
rect 586858 407898 586890 408134
rect 586270 390454 586890 407898
rect 586270 390218 586302 390454
rect 586538 390218 586622 390454
rect 586858 390218 586890 390454
rect 586270 390134 586890 390218
rect 586270 389898 586302 390134
rect 586538 389898 586622 390134
rect 586858 389898 586890 390134
rect 586270 372454 586890 389898
rect 586270 372218 586302 372454
rect 586538 372218 586622 372454
rect 586858 372218 586890 372454
rect 586270 372134 586890 372218
rect 586270 371898 586302 372134
rect 586538 371898 586622 372134
rect 586858 371898 586890 372134
rect 586270 354454 586890 371898
rect 586270 354218 586302 354454
rect 586538 354218 586622 354454
rect 586858 354218 586890 354454
rect 586270 354134 586890 354218
rect 586270 353898 586302 354134
rect 586538 353898 586622 354134
rect 586858 353898 586890 354134
rect 586270 336454 586890 353898
rect 586270 336218 586302 336454
rect 586538 336218 586622 336454
rect 586858 336218 586890 336454
rect 586270 336134 586890 336218
rect 586270 335898 586302 336134
rect 586538 335898 586622 336134
rect 586858 335898 586890 336134
rect 586270 318454 586890 335898
rect 586270 318218 586302 318454
rect 586538 318218 586622 318454
rect 586858 318218 586890 318454
rect 586270 318134 586890 318218
rect 586270 317898 586302 318134
rect 586538 317898 586622 318134
rect 586858 317898 586890 318134
rect 586270 300454 586890 317898
rect 586270 300218 586302 300454
rect 586538 300218 586622 300454
rect 586858 300218 586890 300454
rect 586270 300134 586890 300218
rect 586270 299898 586302 300134
rect 586538 299898 586622 300134
rect 586858 299898 586890 300134
rect 586270 282454 586890 299898
rect 586270 282218 586302 282454
rect 586538 282218 586622 282454
rect 586858 282218 586890 282454
rect 586270 282134 586890 282218
rect 586270 281898 586302 282134
rect 586538 281898 586622 282134
rect 586858 281898 586890 282134
rect 586270 264454 586890 281898
rect 586270 264218 586302 264454
rect 586538 264218 586622 264454
rect 586858 264218 586890 264454
rect 586270 264134 586890 264218
rect 586270 263898 586302 264134
rect 586538 263898 586622 264134
rect 586858 263898 586890 264134
rect 586270 246454 586890 263898
rect 586270 246218 586302 246454
rect 586538 246218 586622 246454
rect 586858 246218 586890 246454
rect 586270 246134 586890 246218
rect 586270 245898 586302 246134
rect 586538 245898 586622 246134
rect 586858 245898 586890 246134
rect 586270 228454 586890 245898
rect 586270 228218 586302 228454
rect 586538 228218 586622 228454
rect 586858 228218 586890 228454
rect 586270 228134 586890 228218
rect 586270 227898 586302 228134
rect 586538 227898 586622 228134
rect 586858 227898 586890 228134
rect 586270 210454 586890 227898
rect 586270 210218 586302 210454
rect 586538 210218 586622 210454
rect 586858 210218 586890 210454
rect 586270 210134 586890 210218
rect 586270 209898 586302 210134
rect 586538 209898 586622 210134
rect 586858 209898 586890 210134
rect 586270 192454 586890 209898
rect 586270 192218 586302 192454
rect 586538 192218 586622 192454
rect 586858 192218 586890 192454
rect 586270 192134 586890 192218
rect 586270 191898 586302 192134
rect 586538 191898 586622 192134
rect 586858 191898 586890 192134
rect 586270 174454 586890 191898
rect 586270 174218 586302 174454
rect 586538 174218 586622 174454
rect 586858 174218 586890 174454
rect 586270 174134 586890 174218
rect 586270 173898 586302 174134
rect 586538 173898 586622 174134
rect 586858 173898 586890 174134
rect 586270 156454 586890 173898
rect 586270 156218 586302 156454
rect 586538 156218 586622 156454
rect 586858 156218 586890 156454
rect 586270 156134 586890 156218
rect 586270 155898 586302 156134
rect 586538 155898 586622 156134
rect 586858 155898 586890 156134
rect 586270 138454 586890 155898
rect 586270 138218 586302 138454
rect 586538 138218 586622 138454
rect 586858 138218 586890 138454
rect 586270 138134 586890 138218
rect 586270 137898 586302 138134
rect 586538 137898 586622 138134
rect 586858 137898 586890 138134
rect 586270 120454 586890 137898
rect 586270 120218 586302 120454
rect 586538 120218 586622 120454
rect 586858 120218 586890 120454
rect 586270 120134 586890 120218
rect 586270 119898 586302 120134
rect 586538 119898 586622 120134
rect 586858 119898 586890 120134
rect 586270 102454 586890 119898
rect 586270 102218 586302 102454
rect 586538 102218 586622 102454
rect 586858 102218 586890 102454
rect 586270 102134 586890 102218
rect 586270 101898 586302 102134
rect 586538 101898 586622 102134
rect 586858 101898 586890 102134
rect 586270 84454 586890 101898
rect 586270 84218 586302 84454
rect 586538 84218 586622 84454
rect 586858 84218 586890 84454
rect 586270 84134 586890 84218
rect 586270 83898 586302 84134
rect 586538 83898 586622 84134
rect 586858 83898 586890 84134
rect 586270 66454 586890 83898
rect 586270 66218 586302 66454
rect 586538 66218 586622 66454
rect 586858 66218 586890 66454
rect 586270 66134 586890 66218
rect 586270 65898 586302 66134
rect 586538 65898 586622 66134
rect 586858 65898 586890 66134
rect 586270 48454 586890 65898
rect 586270 48218 586302 48454
rect 586538 48218 586622 48454
rect 586858 48218 586890 48454
rect 586270 48134 586890 48218
rect 586270 47898 586302 48134
rect 586538 47898 586622 48134
rect 586858 47898 586890 48134
rect 586270 30454 586890 47898
rect 586270 30218 586302 30454
rect 586538 30218 586622 30454
rect 586858 30218 586890 30454
rect 586270 30134 586890 30218
rect 586270 29898 586302 30134
rect 586538 29898 586622 30134
rect 586858 29898 586890 30134
rect 586270 12454 586890 29898
rect 586270 12218 586302 12454
rect 586538 12218 586622 12454
rect 586858 12218 586890 12454
rect 586270 12134 586890 12218
rect 586270 11898 586302 12134
rect 586538 11898 586622 12134
rect 586858 11898 586890 12134
rect 586270 -1306 586890 11898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
<< via4 >>
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 696218 -2698 696454
rect -2614 696218 -2378 696454
rect -2934 695898 -2698 696134
rect -2614 695898 -2378 696134
rect -2934 678218 -2698 678454
rect -2614 678218 -2378 678454
rect -2934 677898 -2698 678134
rect -2614 677898 -2378 678134
rect -2934 660218 -2698 660454
rect -2614 660218 -2378 660454
rect -2934 659898 -2698 660134
rect -2614 659898 -2378 660134
rect -2934 642218 -2698 642454
rect -2614 642218 -2378 642454
rect -2934 641898 -2698 642134
rect -2614 641898 -2378 642134
rect -2934 624218 -2698 624454
rect -2614 624218 -2378 624454
rect -2934 623898 -2698 624134
rect -2614 623898 -2378 624134
rect -2934 606218 -2698 606454
rect -2614 606218 -2378 606454
rect -2934 605898 -2698 606134
rect -2614 605898 -2378 606134
rect -2934 588218 -2698 588454
rect -2614 588218 -2378 588454
rect -2934 587898 -2698 588134
rect -2614 587898 -2378 588134
rect -2934 570218 -2698 570454
rect -2614 570218 -2378 570454
rect -2934 569898 -2698 570134
rect -2614 569898 -2378 570134
rect -2934 552218 -2698 552454
rect -2614 552218 -2378 552454
rect -2934 551898 -2698 552134
rect -2614 551898 -2378 552134
rect -2934 534218 -2698 534454
rect -2614 534218 -2378 534454
rect -2934 533898 -2698 534134
rect -2614 533898 -2378 534134
rect -2934 516218 -2698 516454
rect -2614 516218 -2378 516454
rect -2934 515898 -2698 516134
rect -2614 515898 -2378 516134
rect -2934 498218 -2698 498454
rect -2614 498218 -2378 498454
rect -2934 497898 -2698 498134
rect -2614 497898 -2378 498134
rect -2934 480218 -2698 480454
rect -2614 480218 -2378 480454
rect -2934 479898 -2698 480134
rect -2614 479898 -2378 480134
rect -2934 462218 -2698 462454
rect -2614 462218 -2378 462454
rect -2934 461898 -2698 462134
rect -2614 461898 -2378 462134
rect -2934 444218 -2698 444454
rect -2614 444218 -2378 444454
rect -2934 443898 -2698 444134
rect -2614 443898 -2378 444134
rect -2934 426218 -2698 426454
rect -2614 426218 -2378 426454
rect -2934 425898 -2698 426134
rect -2614 425898 -2378 426134
rect -2934 408218 -2698 408454
rect -2614 408218 -2378 408454
rect -2934 407898 -2698 408134
rect -2614 407898 -2378 408134
rect -2934 390218 -2698 390454
rect -2614 390218 -2378 390454
rect -2934 389898 -2698 390134
rect -2614 389898 -2378 390134
rect -2934 372218 -2698 372454
rect -2614 372218 -2378 372454
rect -2934 371898 -2698 372134
rect -2614 371898 -2378 372134
rect -2934 354218 -2698 354454
rect -2614 354218 -2378 354454
rect -2934 353898 -2698 354134
rect -2614 353898 -2378 354134
rect -2934 336218 -2698 336454
rect -2614 336218 -2378 336454
rect -2934 335898 -2698 336134
rect -2614 335898 -2378 336134
rect -2934 318218 -2698 318454
rect -2614 318218 -2378 318454
rect -2934 317898 -2698 318134
rect -2614 317898 -2378 318134
rect -2934 300218 -2698 300454
rect -2614 300218 -2378 300454
rect -2934 299898 -2698 300134
rect -2614 299898 -2378 300134
rect -2934 282218 -2698 282454
rect -2614 282218 -2378 282454
rect -2934 281898 -2698 282134
rect -2614 281898 -2378 282134
rect -2934 264218 -2698 264454
rect -2614 264218 -2378 264454
rect -2934 263898 -2698 264134
rect -2614 263898 -2378 264134
rect -2934 246218 -2698 246454
rect -2614 246218 -2378 246454
rect -2934 245898 -2698 246134
rect -2614 245898 -2378 246134
rect -2934 228218 -2698 228454
rect -2614 228218 -2378 228454
rect -2934 227898 -2698 228134
rect -2614 227898 -2378 228134
rect -2934 210218 -2698 210454
rect -2614 210218 -2378 210454
rect -2934 209898 -2698 210134
rect -2614 209898 -2378 210134
rect -2934 192218 -2698 192454
rect -2614 192218 -2378 192454
rect -2934 191898 -2698 192134
rect -2614 191898 -2378 192134
rect -2934 174218 -2698 174454
rect -2614 174218 -2378 174454
rect -2934 173898 -2698 174134
rect -2614 173898 -2378 174134
rect -2934 156218 -2698 156454
rect -2614 156218 -2378 156454
rect -2934 155898 -2698 156134
rect -2614 155898 -2378 156134
rect -2934 138218 -2698 138454
rect -2614 138218 -2378 138454
rect -2934 137898 -2698 138134
rect -2614 137898 -2378 138134
rect -2934 120218 -2698 120454
rect -2614 120218 -2378 120454
rect -2934 119898 -2698 120134
rect -2614 119898 -2378 120134
rect -2934 102218 -2698 102454
rect -2614 102218 -2378 102454
rect -2934 101898 -2698 102134
rect -2614 101898 -2378 102134
rect -2934 84218 -2698 84454
rect -2614 84218 -2378 84454
rect -2934 83898 -2698 84134
rect -2614 83898 -2378 84134
rect -2934 66218 -2698 66454
rect -2614 66218 -2378 66454
rect -2934 65898 -2698 66134
rect -2614 65898 -2378 66134
rect -2934 48218 -2698 48454
rect -2614 48218 -2378 48454
rect -2934 47898 -2698 48134
rect -2614 47898 -2378 48134
rect -2934 30218 -2698 30454
rect -2614 30218 -2378 30454
rect -2934 29898 -2698 30134
rect -2614 29898 -2378 30134
rect -2934 12218 -2698 12454
rect -2614 12218 -2378 12454
rect -2934 11898 -2698 12134
rect -2614 11898 -2378 12134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 669218 -1738 669454
rect -1654 669218 -1418 669454
rect -1974 668898 -1738 669134
rect -1654 668898 -1418 669134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 633218 -1738 633454
rect -1654 633218 -1418 633454
rect -1974 632898 -1738 633134
rect -1654 632898 -1418 633134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 597218 -1738 597454
rect -1654 597218 -1418 597454
rect -1974 596898 -1738 597134
rect -1654 596898 -1418 597134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 561218 -1738 561454
rect -1654 561218 -1418 561454
rect -1974 560898 -1738 561134
rect -1654 560898 -1418 561134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 525218 -1738 525454
rect -1654 525218 -1418 525454
rect -1974 524898 -1738 525134
rect -1654 524898 -1418 525134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 489218 -1738 489454
rect -1654 489218 -1418 489454
rect -1974 488898 -1738 489134
rect -1654 488898 -1418 489134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 453218 -1738 453454
rect -1654 453218 -1418 453454
rect -1974 452898 -1738 453134
rect -1654 452898 -1418 453134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 417218 -1738 417454
rect -1654 417218 -1418 417454
rect -1974 416898 -1738 417134
rect -1654 416898 -1418 417134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 381218 -1738 381454
rect -1654 381218 -1418 381454
rect -1974 380898 -1738 381134
rect -1654 380898 -1418 381134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 345218 -1738 345454
rect -1654 345218 -1418 345454
rect -1974 344898 -1738 345134
rect -1654 344898 -1418 345134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 309218 -1738 309454
rect -1654 309218 -1418 309454
rect -1974 308898 -1738 309134
rect -1654 308898 -1418 309134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 273218 -1738 273454
rect -1654 273218 -1418 273454
rect -1974 272898 -1738 273134
rect -1654 272898 -1418 273134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 237218 -1738 237454
rect -1654 237218 -1418 237454
rect -1974 236898 -1738 237134
rect -1654 236898 -1418 237134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 201218 -1738 201454
rect -1654 201218 -1418 201454
rect -1974 200898 -1738 201134
rect -1654 200898 -1418 201134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 165218 -1738 165454
rect -1654 165218 -1418 165454
rect -1974 164898 -1738 165134
rect -1654 164898 -1418 165134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 129218 -1738 129454
rect -1654 129218 -1418 129454
rect -1974 128898 -1738 129134
rect -1654 128898 -1418 129134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 93218 -1738 93454
rect -1654 93218 -1418 93454
rect -1974 92898 -1738 93134
rect -1654 92898 -1418 93134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 57218 -1738 57454
rect -1654 57218 -1418 57454
rect -1974 56898 -1738 57134
rect -1654 56898 -1418 57134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 21218 -1738 21454
rect -1654 21218 -1418 21454
rect -1974 20898 -1738 21134
rect -1654 20898 -1418 21134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 669218 2062 669454
rect 2146 669218 2382 669454
rect 1826 668898 2062 669134
rect 2146 668898 2382 669134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 633218 2062 633454
rect 2146 633218 2382 633454
rect 1826 632898 2062 633134
rect 2146 632898 2382 633134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 597218 2062 597454
rect 2146 597218 2382 597454
rect 1826 596898 2062 597134
rect 2146 596898 2382 597134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 561218 2062 561454
rect 2146 561218 2382 561454
rect 1826 560898 2062 561134
rect 2146 560898 2382 561134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 525218 2062 525454
rect 2146 525218 2382 525454
rect 1826 524898 2062 525134
rect 2146 524898 2382 525134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 489218 2062 489454
rect 2146 489218 2382 489454
rect 1826 488898 2062 489134
rect 2146 488898 2382 489134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 453218 2062 453454
rect 2146 453218 2382 453454
rect 1826 452898 2062 453134
rect 2146 452898 2382 453134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 417218 2062 417454
rect 2146 417218 2382 417454
rect 1826 416898 2062 417134
rect 2146 416898 2382 417134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 381218 2062 381454
rect 2146 381218 2382 381454
rect 1826 380898 2062 381134
rect 2146 380898 2382 381134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 345218 2062 345454
rect 2146 345218 2382 345454
rect 1826 344898 2062 345134
rect 2146 344898 2382 345134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 309218 2062 309454
rect 2146 309218 2382 309454
rect 1826 308898 2062 309134
rect 2146 308898 2382 309134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 273218 2062 273454
rect 2146 273218 2382 273454
rect 1826 272898 2062 273134
rect 2146 272898 2382 273134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 237218 2062 237454
rect 2146 237218 2382 237454
rect 1826 236898 2062 237134
rect 2146 236898 2382 237134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 201218 2062 201454
rect 2146 201218 2382 201454
rect 1826 200898 2062 201134
rect 2146 200898 2382 201134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 165218 2062 165454
rect 2146 165218 2382 165454
rect 1826 164898 2062 165134
rect 2146 164898 2382 165134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 129218 2062 129454
rect 2146 129218 2382 129454
rect 1826 128898 2062 129134
rect 2146 128898 2382 129134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 93218 2062 93454
rect 2146 93218 2382 93454
rect 1826 92898 2062 93134
rect 2146 92898 2382 93134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 57218 2062 57454
rect 2146 57218 2382 57454
rect 1826 56898 2062 57134
rect 2146 56898 2382 57134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 21218 2062 21454
rect 2146 21218 2382 21454
rect 1826 20898 2062 21134
rect 2146 20898 2382 21134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 10826 705562 11062 705798
rect 11146 705562 11382 705798
rect 10826 705242 11062 705478
rect 11146 705242 11382 705478
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 19826 704602 20062 704838
rect 20146 704602 20382 704838
rect 19826 704282 20062 704518
rect 20146 704282 20382 704518
rect 19826 687218 20062 687454
rect 20146 687218 20382 687454
rect 19826 686898 20062 687134
rect 20146 686898 20382 687134
rect 28826 705562 29062 705798
rect 29146 705562 29382 705798
rect 28826 705242 29062 705478
rect 29146 705242 29382 705478
rect 28826 696218 29062 696454
rect 29146 696218 29382 696454
rect 28826 695898 29062 696134
rect 29146 695898 29382 696134
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 46826 705562 47062 705798
rect 47146 705562 47382 705798
rect 46826 705242 47062 705478
rect 47146 705242 47382 705478
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 55826 704602 56062 704838
rect 56146 704602 56382 704838
rect 55826 704282 56062 704518
rect 56146 704282 56382 704518
rect 55826 687218 56062 687454
rect 56146 687218 56382 687454
rect 55826 686898 56062 687134
rect 56146 686898 56382 687134
rect 64826 705562 65062 705798
rect 65146 705562 65382 705798
rect 64826 705242 65062 705478
rect 65146 705242 65382 705478
rect 64826 696218 65062 696454
rect 65146 696218 65382 696454
rect 64826 695898 65062 696134
rect 65146 695898 65382 696134
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 82826 705562 83062 705798
rect 83146 705562 83382 705798
rect 82826 705242 83062 705478
rect 83146 705242 83382 705478
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 91826 704602 92062 704838
rect 92146 704602 92382 704838
rect 91826 704282 92062 704518
rect 92146 704282 92382 704518
rect 91826 687218 92062 687454
rect 92146 687218 92382 687454
rect 91826 686898 92062 687134
rect 92146 686898 92382 687134
rect 100826 705562 101062 705798
rect 101146 705562 101382 705798
rect 100826 705242 101062 705478
rect 101146 705242 101382 705478
rect 100826 696218 101062 696454
rect 101146 696218 101382 696454
rect 100826 695898 101062 696134
rect 101146 695898 101382 696134
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 118826 705562 119062 705798
rect 119146 705562 119382 705798
rect 118826 705242 119062 705478
rect 119146 705242 119382 705478
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 127826 704602 128062 704838
rect 128146 704602 128382 704838
rect 127826 704282 128062 704518
rect 128146 704282 128382 704518
rect 127826 687218 128062 687454
rect 128146 687218 128382 687454
rect 127826 686898 128062 687134
rect 128146 686898 128382 687134
rect 136826 705562 137062 705798
rect 137146 705562 137382 705798
rect 136826 705242 137062 705478
rect 137146 705242 137382 705478
rect 136826 696218 137062 696454
rect 137146 696218 137382 696454
rect 136826 695898 137062 696134
rect 137146 695898 137382 696134
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 154826 705562 155062 705798
rect 155146 705562 155382 705798
rect 154826 705242 155062 705478
rect 155146 705242 155382 705478
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 163826 704602 164062 704838
rect 164146 704602 164382 704838
rect 163826 704282 164062 704518
rect 164146 704282 164382 704518
rect 163826 687218 164062 687454
rect 164146 687218 164382 687454
rect 163826 686898 164062 687134
rect 164146 686898 164382 687134
rect 172826 705562 173062 705798
rect 173146 705562 173382 705798
rect 172826 705242 173062 705478
rect 173146 705242 173382 705478
rect 172826 696218 173062 696454
rect 173146 696218 173382 696454
rect 172826 695898 173062 696134
rect 173146 695898 173382 696134
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 190826 705562 191062 705798
rect 191146 705562 191382 705798
rect 190826 705242 191062 705478
rect 191146 705242 191382 705478
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 199826 704602 200062 704838
rect 200146 704602 200382 704838
rect 199826 704282 200062 704518
rect 200146 704282 200382 704518
rect 199826 687218 200062 687454
rect 200146 687218 200382 687454
rect 199826 686898 200062 687134
rect 200146 686898 200382 687134
rect 208826 705562 209062 705798
rect 209146 705562 209382 705798
rect 208826 705242 209062 705478
rect 209146 705242 209382 705478
rect 208826 696218 209062 696454
rect 209146 696218 209382 696454
rect 208826 695898 209062 696134
rect 209146 695898 209382 696134
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 226826 705562 227062 705798
rect 227146 705562 227382 705798
rect 226826 705242 227062 705478
rect 227146 705242 227382 705478
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 235826 704602 236062 704838
rect 236146 704602 236382 704838
rect 235826 704282 236062 704518
rect 236146 704282 236382 704518
rect 235826 687218 236062 687454
rect 236146 687218 236382 687454
rect 235826 686898 236062 687134
rect 236146 686898 236382 687134
rect 244826 705562 245062 705798
rect 245146 705562 245382 705798
rect 244826 705242 245062 705478
rect 245146 705242 245382 705478
rect 244826 696218 245062 696454
rect 245146 696218 245382 696454
rect 244826 695898 245062 696134
rect 245146 695898 245382 696134
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 262826 705562 263062 705798
rect 263146 705562 263382 705798
rect 262826 705242 263062 705478
rect 263146 705242 263382 705478
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 271826 704602 272062 704838
rect 272146 704602 272382 704838
rect 271826 704282 272062 704518
rect 272146 704282 272382 704518
rect 271826 687218 272062 687454
rect 272146 687218 272382 687454
rect 271826 686898 272062 687134
rect 272146 686898 272382 687134
rect 280826 705562 281062 705798
rect 281146 705562 281382 705798
rect 280826 705242 281062 705478
rect 281146 705242 281382 705478
rect 280826 696218 281062 696454
rect 281146 696218 281382 696454
rect 280826 695898 281062 696134
rect 281146 695898 281382 696134
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 298826 705562 299062 705798
rect 299146 705562 299382 705798
rect 298826 705242 299062 705478
rect 299146 705242 299382 705478
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 307826 704602 308062 704838
rect 308146 704602 308382 704838
rect 307826 704282 308062 704518
rect 308146 704282 308382 704518
rect 307826 687218 308062 687454
rect 308146 687218 308382 687454
rect 307826 686898 308062 687134
rect 308146 686898 308382 687134
rect 316826 705562 317062 705798
rect 317146 705562 317382 705798
rect 316826 705242 317062 705478
rect 317146 705242 317382 705478
rect 316826 696218 317062 696454
rect 317146 696218 317382 696454
rect 316826 695898 317062 696134
rect 317146 695898 317382 696134
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 334826 705562 335062 705798
rect 335146 705562 335382 705798
rect 334826 705242 335062 705478
rect 335146 705242 335382 705478
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 343826 704602 344062 704838
rect 344146 704602 344382 704838
rect 343826 704282 344062 704518
rect 344146 704282 344382 704518
rect 343826 687218 344062 687454
rect 344146 687218 344382 687454
rect 343826 686898 344062 687134
rect 344146 686898 344382 687134
rect 352826 705562 353062 705798
rect 353146 705562 353382 705798
rect 352826 705242 353062 705478
rect 353146 705242 353382 705478
rect 352826 696218 353062 696454
rect 353146 696218 353382 696454
rect 352826 695898 353062 696134
rect 353146 695898 353382 696134
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 370826 705562 371062 705798
rect 371146 705562 371382 705798
rect 370826 705242 371062 705478
rect 371146 705242 371382 705478
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 379826 704602 380062 704838
rect 380146 704602 380382 704838
rect 379826 704282 380062 704518
rect 380146 704282 380382 704518
rect 379826 687218 380062 687454
rect 380146 687218 380382 687454
rect 379826 686898 380062 687134
rect 380146 686898 380382 687134
rect 388826 705562 389062 705798
rect 389146 705562 389382 705798
rect 388826 705242 389062 705478
rect 389146 705242 389382 705478
rect 388826 696218 389062 696454
rect 389146 696218 389382 696454
rect 388826 695898 389062 696134
rect 389146 695898 389382 696134
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 406826 705562 407062 705798
rect 407146 705562 407382 705798
rect 406826 705242 407062 705478
rect 407146 705242 407382 705478
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 415826 704602 416062 704838
rect 416146 704602 416382 704838
rect 415826 704282 416062 704518
rect 416146 704282 416382 704518
rect 415826 687218 416062 687454
rect 416146 687218 416382 687454
rect 415826 686898 416062 687134
rect 416146 686898 416382 687134
rect 424826 705562 425062 705798
rect 425146 705562 425382 705798
rect 424826 705242 425062 705478
rect 425146 705242 425382 705478
rect 424826 696218 425062 696454
rect 425146 696218 425382 696454
rect 424826 695898 425062 696134
rect 425146 695898 425382 696134
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 442826 705562 443062 705798
rect 443146 705562 443382 705798
rect 442826 705242 443062 705478
rect 443146 705242 443382 705478
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 451826 704602 452062 704838
rect 452146 704602 452382 704838
rect 451826 704282 452062 704518
rect 452146 704282 452382 704518
rect 451826 687218 452062 687454
rect 452146 687218 452382 687454
rect 451826 686898 452062 687134
rect 452146 686898 452382 687134
rect 460826 705562 461062 705798
rect 461146 705562 461382 705798
rect 460826 705242 461062 705478
rect 461146 705242 461382 705478
rect 460826 696218 461062 696454
rect 461146 696218 461382 696454
rect 460826 695898 461062 696134
rect 461146 695898 461382 696134
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 478826 705562 479062 705798
rect 479146 705562 479382 705798
rect 478826 705242 479062 705478
rect 479146 705242 479382 705478
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 487826 704602 488062 704838
rect 488146 704602 488382 704838
rect 487826 704282 488062 704518
rect 488146 704282 488382 704518
rect 487826 687218 488062 687454
rect 488146 687218 488382 687454
rect 487826 686898 488062 687134
rect 488146 686898 488382 687134
rect 496826 705562 497062 705798
rect 497146 705562 497382 705798
rect 496826 705242 497062 705478
rect 497146 705242 497382 705478
rect 496826 696218 497062 696454
rect 497146 696218 497382 696454
rect 496826 695898 497062 696134
rect 497146 695898 497382 696134
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 514826 705562 515062 705798
rect 515146 705562 515382 705798
rect 514826 705242 515062 705478
rect 515146 705242 515382 705478
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 523826 704602 524062 704838
rect 524146 704602 524382 704838
rect 523826 704282 524062 704518
rect 524146 704282 524382 704518
rect 523826 687218 524062 687454
rect 524146 687218 524382 687454
rect 523826 686898 524062 687134
rect 524146 686898 524382 687134
rect 532826 705562 533062 705798
rect 533146 705562 533382 705798
rect 532826 705242 533062 705478
rect 533146 705242 533382 705478
rect 532826 696218 533062 696454
rect 533146 696218 533382 696454
rect 532826 695898 533062 696134
rect 533146 695898 533382 696134
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 550826 705562 551062 705798
rect 551146 705562 551382 705798
rect 550826 705242 551062 705478
rect 551146 705242 551382 705478
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 559826 704602 560062 704838
rect 560146 704602 560382 704838
rect 559826 704282 560062 704518
rect 560146 704282 560382 704518
rect 559826 687218 560062 687454
rect 560146 687218 560382 687454
rect 559826 686898 560062 687134
rect 560146 686898 560382 687134
rect 10826 678218 11062 678454
rect 11146 678218 11382 678454
rect 10826 677898 11062 678134
rect 11146 677898 11382 678134
rect 22916 678218 23152 678454
rect 22916 677898 23152 678134
rect 28847 678218 29083 678454
rect 28847 677898 29083 678134
rect 49916 678218 50152 678454
rect 49916 677898 50152 678134
rect 55847 678218 56083 678454
rect 55847 677898 56083 678134
rect 76916 678218 77152 678454
rect 76916 677898 77152 678134
rect 82847 678218 83083 678454
rect 82847 677898 83083 678134
rect 103916 678218 104152 678454
rect 103916 677898 104152 678134
rect 109847 678218 110083 678454
rect 109847 677898 110083 678134
rect 130916 678218 131152 678454
rect 130916 677898 131152 678134
rect 136847 678218 137083 678454
rect 136847 677898 137083 678134
rect 157916 678218 158152 678454
rect 157916 677898 158152 678134
rect 163847 678218 164083 678454
rect 163847 677898 164083 678134
rect 184916 678218 185152 678454
rect 184916 677898 185152 678134
rect 190847 678218 191083 678454
rect 190847 677898 191083 678134
rect 211916 678218 212152 678454
rect 211916 677898 212152 678134
rect 217847 678218 218083 678454
rect 217847 677898 218083 678134
rect 238916 678218 239152 678454
rect 238916 677898 239152 678134
rect 244847 678218 245083 678454
rect 244847 677898 245083 678134
rect 265916 678218 266152 678454
rect 265916 677898 266152 678134
rect 271847 678218 272083 678454
rect 271847 677898 272083 678134
rect 292916 678218 293152 678454
rect 292916 677898 293152 678134
rect 298847 678218 299083 678454
rect 298847 677898 299083 678134
rect 319916 678218 320152 678454
rect 319916 677898 320152 678134
rect 325847 678218 326083 678454
rect 325847 677898 326083 678134
rect 346916 678218 347152 678454
rect 346916 677898 347152 678134
rect 352847 678218 353083 678454
rect 352847 677898 353083 678134
rect 373916 678218 374152 678454
rect 373916 677898 374152 678134
rect 379847 678218 380083 678454
rect 379847 677898 380083 678134
rect 400916 678218 401152 678454
rect 400916 677898 401152 678134
rect 406847 678218 407083 678454
rect 406847 677898 407083 678134
rect 427916 678218 428152 678454
rect 427916 677898 428152 678134
rect 433847 678218 434083 678454
rect 433847 677898 434083 678134
rect 454916 678218 455152 678454
rect 454916 677898 455152 678134
rect 460847 678218 461083 678454
rect 460847 677898 461083 678134
rect 481916 678218 482152 678454
rect 481916 677898 482152 678134
rect 487847 678218 488083 678454
rect 487847 677898 488083 678134
rect 508916 678218 509152 678454
rect 508916 677898 509152 678134
rect 514847 678218 515083 678454
rect 514847 677898 515083 678134
rect 535916 678218 536152 678454
rect 535916 677898 536152 678134
rect 541847 678218 542083 678454
rect 541847 677898 542083 678134
rect 19952 669218 20188 669454
rect 19952 668898 20188 669134
rect 25882 669218 26118 669454
rect 25882 668898 26118 669134
rect 31813 669218 32049 669454
rect 31813 668898 32049 669134
rect 46952 669218 47188 669454
rect 46952 668898 47188 669134
rect 52882 669218 53118 669454
rect 52882 668898 53118 669134
rect 58813 669218 59049 669454
rect 58813 668898 59049 669134
rect 73952 669218 74188 669454
rect 73952 668898 74188 669134
rect 79882 669218 80118 669454
rect 79882 668898 80118 669134
rect 85813 669218 86049 669454
rect 85813 668898 86049 669134
rect 100952 669218 101188 669454
rect 100952 668898 101188 669134
rect 106882 669218 107118 669454
rect 106882 668898 107118 669134
rect 112813 669218 113049 669454
rect 112813 668898 113049 669134
rect 127952 669218 128188 669454
rect 127952 668898 128188 669134
rect 133882 669218 134118 669454
rect 133882 668898 134118 669134
rect 139813 669218 140049 669454
rect 139813 668898 140049 669134
rect 154952 669218 155188 669454
rect 154952 668898 155188 669134
rect 160882 669218 161118 669454
rect 160882 668898 161118 669134
rect 166813 669218 167049 669454
rect 166813 668898 167049 669134
rect 181952 669218 182188 669454
rect 181952 668898 182188 669134
rect 187882 669218 188118 669454
rect 187882 668898 188118 669134
rect 193813 669218 194049 669454
rect 193813 668898 194049 669134
rect 208952 669218 209188 669454
rect 208952 668898 209188 669134
rect 214882 669218 215118 669454
rect 214882 668898 215118 669134
rect 220813 669218 221049 669454
rect 220813 668898 221049 669134
rect 235952 669218 236188 669454
rect 235952 668898 236188 669134
rect 241882 669218 242118 669454
rect 241882 668898 242118 669134
rect 247813 669218 248049 669454
rect 247813 668898 248049 669134
rect 262952 669218 263188 669454
rect 262952 668898 263188 669134
rect 268882 669218 269118 669454
rect 268882 668898 269118 669134
rect 274813 669218 275049 669454
rect 274813 668898 275049 669134
rect 289952 669218 290188 669454
rect 289952 668898 290188 669134
rect 295882 669218 296118 669454
rect 295882 668898 296118 669134
rect 301813 669218 302049 669454
rect 301813 668898 302049 669134
rect 316952 669218 317188 669454
rect 316952 668898 317188 669134
rect 322882 669218 323118 669454
rect 322882 668898 323118 669134
rect 328813 669218 329049 669454
rect 328813 668898 329049 669134
rect 343952 669218 344188 669454
rect 343952 668898 344188 669134
rect 349882 669218 350118 669454
rect 349882 668898 350118 669134
rect 355813 669218 356049 669454
rect 355813 668898 356049 669134
rect 370952 669218 371188 669454
rect 370952 668898 371188 669134
rect 376882 669218 377118 669454
rect 376882 668898 377118 669134
rect 382813 669218 383049 669454
rect 382813 668898 383049 669134
rect 397952 669218 398188 669454
rect 397952 668898 398188 669134
rect 403882 669218 404118 669454
rect 403882 668898 404118 669134
rect 409813 669218 410049 669454
rect 409813 668898 410049 669134
rect 424952 669218 425188 669454
rect 424952 668898 425188 669134
rect 430882 669218 431118 669454
rect 430882 668898 431118 669134
rect 436813 669218 437049 669454
rect 436813 668898 437049 669134
rect 451952 669218 452188 669454
rect 451952 668898 452188 669134
rect 457882 669218 458118 669454
rect 457882 668898 458118 669134
rect 463813 669218 464049 669454
rect 463813 668898 464049 669134
rect 478952 669218 479188 669454
rect 478952 668898 479188 669134
rect 484882 669218 485118 669454
rect 484882 668898 485118 669134
rect 490813 669218 491049 669454
rect 490813 668898 491049 669134
rect 505952 669218 506188 669454
rect 505952 668898 506188 669134
rect 511882 669218 512118 669454
rect 511882 668898 512118 669134
rect 517813 669218 518049 669454
rect 517813 668898 518049 669134
rect 532952 669218 533188 669454
rect 532952 668898 533188 669134
rect 538882 669218 539118 669454
rect 538882 668898 539118 669134
rect 544813 669218 545049 669454
rect 544813 668898 545049 669134
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 19826 661158 20062 661394
rect 20146 661158 20382 661394
rect 19826 660838 20062 661074
rect 20146 660838 20382 661074
rect 28826 660218 29062 660454
rect 29146 660218 29382 660454
rect 28826 659898 29062 660134
rect 29146 659898 29382 660134
rect 37826 661158 38062 661394
rect 38146 661158 38382 661394
rect 37826 660838 38062 661074
rect 38146 660838 38382 661074
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 55826 661158 56062 661394
rect 56146 661158 56382 661394
rect 55826 660838 56062 661074
rect 56146 660838 56382 661074
rect 64826 660218 65062 660454
rect 65146 660218 65382 660454
rect 64826 659898 65062 660134
rect 65146 659898 65382 660134
rect 73826 661158 74062 661394
rect 74146 661158 74382 661394
rect 73826 660838 74062 661074
rect 74146 660838 74382 661074
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 91826 661158 92062 661394
rect 92146 661158 92382 661394
rect 91826 660838 92062 661074
rect 92146 660838 92382 661074
rect 100826 660218 101062 660454
rect 101146 660218 101382 660454
rect 100826 659898 101062 660134
rect 101146 659898 101382 660134
rect 109826 661158 110062 661394
rect 110146 661158 110382 661394
rect 109826 660838 110062 661074
rect 110146 660838 110382 661074
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 127826 661158 128062 661394
rect 128146 661158 128382 661394
rect 127826 660838 128062 661074
rect 128146 660838 128382 661074
rect 136826 660218 137062 660454
rect 137146 660218 137382 660454
rect 136826 659898 137062 660134
rect 137146 659898 137382 660134
rect 145826 661158 146062 661394
rect 146146 661158 146382 661394
rect 145826 660838 146062 661074
rect 146146 660838 146382 661074
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 163826 661158 164062 661394
rect 164146 661158 164382 661394
rect 163826 660838 164062 661074
rect 164146 660838 164382 661074
rect 172826 660218 173062 660454
rect 173146 660218 173382 660454
rect 172826 659898 173062 660134
rect 173146 659898 173382 660134
rect 181826 661158 182062 661394
rect 182146 661158 182382 661394
rect 181826 660838 182062 661074
rect 182146 660838 182382 661074
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 199826 661158 200062 661394
rect 200146 661158 200382 661394
rect 199826 660838 200062 661074
rect 200146 660838 200382 661074
rect 208826 660218 209062 660454
rect 209146 660218 209382 660454
rect 208826 659898 209062 660134
rect 209146 659898 209382 660134
rect 217826 661158 218062 661394
rect 218146 661158 218382 661394
rect 217826 660838 218062 661074
rect 218146 660838 218382 661074
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 235826 661158 236062 661394
rect 236146 661158 236382 661394
rect 235826 660838 236062 661074
rect 236146 660838 236382 661074
rect 244826 660218 245062 660454
rect 245146 660218 245382 660454
rect 244826 659898 245062 660134
rect 245146 659898 245382 660134
rect 253826 661158 254062 661394
rect 254146 661158 254382 661394
rect 253826 660838 254062 661074
rect 254146 660838 254382 661074
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 271826 661158 272062 661394
rect 272146 661158 272382 661394
rect 271826 660838 272062 661074
rect 272146 660838 272382 661074
rect 280826 660218 281062 660454
rect 281146 660218 281382 660454
rect 280826 659898 281062 660134
rect 281146 659898 281382 660134
rect 289826 661158 290062 661394
rect 290146 661158 290382 661394
rect 289826 660838 290062 661074
rect 290146 660838 290382 661074
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 307826 661158 308062 661394
rect 308146 661158 308382 661394
rect 307826 660838 308062 661074
rect 308146 660838 308382 661074
rect 316826 660218 317062 660454
rect 317146 660218 317382 660454
rect 316826 659898 317062 660134
rect 317146 659898 317382 660134
rect 325826 661158 326062 661394
rect 326146 661158 326382 661394
rect 325826 660838 326062 661074
rect 326146 660838 326382 661074
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 343826 661158 344062 661394
rect 344146 661158 344382 661394
rect 343826 660838 344062 661074
rect 344146 660838 344382 661074
rect 352826 660218 353062 660454
rect 353146 660218 353382 660454
rect 352826 659898 353062 660134
rect 353146 659898 353382 660134
rect 361826 661158 362062 661394
rect 362146 661158 362382 661394
rect 361826 660838 362062 661074
rect 362146 660838 362382 661074
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 379826 661158 380062 661394
rect 380146 661158 380382 661394
rect 379826 660838 380062 661074
rect 380146 660838 380382 661074
rect 388826 660218 389062 660454
rect 389146 660218 389382 660454
rect 388826 659898 389062 660134
rect 389146 659898 389382 660134
rect 397826 661158 398062 661394
rect 398146 661158 398382 661394
rect 397826 660838 398062 661074
rect 398146 660838 398382 661074
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 415826 661158 416062 661394
rect 416146 661158 416382 661394
rect 415826 660838 416062 661074
rect 416146 660838 416382 661074
rect 424826 660218 425062 660454
rect 425146 660218 425382 660454
rect 424826 659898 425062 660134
rect 425146 659898 425382 660134
rect 433826 661158 434062 661394
rect 434146 661158 434382 661394
rect 433826 660838 434062 661074
rect 434146 660838 434382 661074
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 451826 661158 452062 661394
rect 452146 661158 452382 661394
rect 451826 660838 452062 661074
rect 452146 660838 452382 661074
rect 460826 660218 461062 660454
rect 461146 660218 461382 660454
rect 460826 659898 461062 660134
rect 461146 659898 461382 660134
rect 469826 661158 470062 661394
rect 470146 661158 470382 661394
rect 469826 660838 470062 661074
rect 470146 660838 470382 661074
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 487826 661158 488062 661394
rect 488146 661158 488382 661394
rect 487826 660838 488062 661074
rect 488146 660838 488382 661074
rect 496826 660218 497062 660454
rect 497146 660218 497382 660454
rect 496826 659898 497062 660134
rect 497146 659898 497382 660134
rect 505826 661158 506062 661394
rect 506146 661158 506382 661394
rect 505826 660838 506062 661074
rect 506146 660838 506382 661074
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 523826 661158 524062 661394
rect 524146 661158 524382 661394
rect 523826 660838 524062 661074
rect 524146 660838 524382 661074
rect 532826 660218 533062 660454
rect 533146 660218 533382 660454
rect 532826 659898 533062 660134
rect 533146 659898 533382 660134
rect 541826 661158 542062 661394
rect 542146 661158 542382 661394
rect 541826 660838 542062 661074
rect 542146 660838 542382 661074
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 19952 651218 20188 651454
rect 19952 650898 20188 651134
rect 25882 651218 26118 651454
rect 25882 650898 26118 651134
rect 31813 651218 32049 651454
rect 31813 650898 32049 651134
rect 46952 651218 47188 651454
rect 46952 650898 47188 651134
rect 52882 651218 53118 651454
rect 52882 650898 53118 651134
rect 58813 651218 59049 651454
rect 58813 650898 59049 651134
rect 73952 651218 74188 651454
rect 73952 650898 74188 651134
rect 79882 651218 80118 651454
rect 79882 650898 80118 651134
rect 85813 651218 86049 651454
rect 85813 650898 86049 651134
rect 100952 651218 101188 651454
rect 100952 650898 101188 651134
rect 106882 651218 107118 651454
rect 106882 650898 107118 651134
rect 112813 651218 113049 651454
rect 112813 650898 113049 651134
rect 127952 651218 128188 651454
rect 127952 650898 128188 651134
rect 133882 651218 134118 651454
rect 133882 650898 134118 651134
rect 139813 651218 140049 651454
rect 139813 650898 140049 651134
rect 154952 651218 155188 651454
rect 154952 650898 155188 651134
rect 160882 651218 161118 651454
rect 160882 650898 161118 651134
rect 166813 651218 167049 651454
rect 166813 650898 167049 651134
rect 181952 651218 182188 651454
rect 181952 650898 182188 651134
rect 187882 651218 188118 651454
rect 187882 650898 188118 651134
rect 193813 651218 194049 651454
rect 193813 650898 194049 651134
rect 208952 651218 209188 651454
rect 208952 650898 209188 651134
rect 214882 651218 215118 651454
rect 214882 650898 215118 651134
rect 220813 651218 221049 651454
rect 220813 650898 221049 651134
rect 235952 651218 236188 651454
rect 235952 650898 236188 651134
rect 241882 651218 242118 651454
rect 241882 650898 242118 651134
rect 247813 651218 248049 651454
rect 247813 650898 248049 651134
rect 262952 651218 263188 651454
rect 262952 650898 263188 651134
rect 268882 651218 269118 651454
rect 268882 650898 269118 651134
rect 274813 651218 275049 651454
rect 274813 650898 275049 651134
rect 289952 651218 290188 651454
rect 289952 650898 290188 651134
rect 295882 651218 296118 651454
rect 295882 650898 296118 651134
rect 301813 651218 302049 651454
rect 301813 650898 302049 651134
rect 316952 651218 317188 651454
rect 316952 650898 317188 651134
rect 322882 651218 323118 651454
rect 322882 650898 323118 651134
rect 328813 651218 329049 651454
rect 328813 650898 329049 651134
rect 343952 651218 344188 651454
rect 343952 650898 344188 651134
rect 349882 651218 350118 651454
rect 349882 650898 350118 651134
rect 355813 651218 356049 651454
rect 355813 650898 356049 651134
rect 370952 651218 371188 651454
rect 370952 650898 371188 651134
rect 376882 651218 377118 651454
rect 376882 650898 377118 651134
rect 382813 651218 383049 651454
rect 382813 650898 383049 651134
rect 397952 651218 398188 651454
rect 397952 650898 398188 651134
rect 403882 651218 404118 651454
rect 403882 650898 404118 651134
rect 409813 651218 410049 651454
rect 409813 650898 410049 651134
rect 424952 651218 425188 651454
rect 424952 650898 425188 651134
rect 430882 651218 431118 651454
rect 430882 650898 431118 651134
rect 436813 651218 437049 651454
rect 436813 650898 437049 651134
rect 451952 651218 452188 651454
rect 451952 650898 452188 651134
rect 457882 651218 458118 651454
rect 457882 650898 458118 651134
rect 463813 651218 464049 651454
rect 463813 650898 464049 651134
rect 478952 651218 479188 651454
rect 478952 650898 479188 651134
rect 484882 651218 485118 651454
rect 484882 650898 485118 651134
rect 490813 651218 491049 651454
rect 490813 650898 491049 651134
rect 505952 651218 506188 651454
rect 505952 650898 506188 651134
rect 511882 651218 512118 651454
rect 511882 650898 512118 651134
rect 517813 651218 518049 651454
rect 517813 650898 518049 651134
rect 532952 651218 533188 651454
rect 532952 650898 533188 651134
rect 538882 651218 539118 651454
rect 538882 650898 539118 651134
rect 544813 651218 545049 651454
rect 544813 650898 545049 651134
rect 559826 651218 560062 651454
rect 560146 651218 560382 651454
rect 559826 650898 560062 651134
rect 560146 650898 560382 651134
rect 10826 642218 11062 642454
rect 11146 642218 11382 642454
rect 10826 641898 11062 642134
rect 11146 641898 11382 642134
rect 22916 642218 23152 642454
rect 22916 641898 23152 642134
rect 28847 642218 29083 642454
rect 28847 641898 29083 642134
rect 49916 642218 50152 642454
rect 49916 641898 50152 642134
rect 55847 642218 56083 642454
rect 55847 641898 56083 642134
rect 76916 642218 77152 642454
rect 76916 641898 77152 642134
rect 82847 642218 83083 642454
rect 82847 641898 83083 642134
rect 103916 642218 104152 642454
rect 103916 641898 104152 642134
rect 109847 642218 110083 642454
rect 109847 641898 110083 642134
rect 130916 642218 131152 642454
rect 130916 641898 131152 642134
rect 136847 642218 137083 642454
rect 136847 641898 137083 642134
rect 157916 642218 158152 642454
rect 157916 641898 158152 642134
rect 163847 642218 164083 642454
rect 163847 641898 164083 642134
rect 184916 642218 185152 642454
rect 184916 641898 185152 642134
rect 190847 642218 191083 642454
rect 190847 641898 191083 642134
rect 211916 642218 212152 642454
rect 211916 641898 212152 642134
rect 217847 642218 218083 642454
rect 217847 641898 218083 642134
rect 238916 642218 239152 642454
rect 238916 641898 239152 642134
rect 244847 642218 245083 642454
rect 244847 641898 245083 642134
rect 265916 642218 266152 642454
rect 265916 641898 266152 642134
rect 271847 642218 272083 642454
rect 271847 641898 272083 642134
rect 292916 642218 293152 642454
rect 292916 641898 293152 642134
rect 298847 642218 299083 642454
rect 298847 641898 299083 642134
rect 319916 642218 320152 642454
rect 319916 641898 320152 642134
rect 325847 642218 326083 642454
rect 325847 641898 326083 642134
rect 346916 642218 347152 642454
rect 346916 641898 347152 642134
rect 352847 642218 353083 642454
rect 352847 641898 353083 642134
rect 373916 642218 374152 642454
rect 373916 641898 374152 642134
rect 379847 642218 380083 642454
rect 379847 641898 380083 642134
rect 400916 642218 401152 642454
rect 400916 641898 401152 642134
rect 406847 642218 407083 642454
rect 406847 641898 407083 642134
rect 427916 642218 428152 642454
rect 427916 641898 428152 642134
rect 433847 642218 434083 642454
rect 433847 641898 434083 642134
rect 454916 642218 455152 642454
rect 454916 641898 455152 642134
rect 460847 642218 461083 642454
rect 460847 641898 461083 642134
rect 481916 642218 482152 642454
rect 481916 641898 482152 642134
rect 487847 642218 488083 642454
rect 487847 641898 488083 642134
rect 508916 642218 509152 642454
rect 508916 641898 509152 642134
rect 514847 642218 515083 642454
rect 514847 641898 515083 642134
rect 535916 642218 536152 642454
rect 535916 641898 536152 642134
rect 541847 642218 542083 642454
rect 541847 641898 542083 642134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 28826 634158 29062 634394
rect 29146 634158 29382 634394
rect 28826 633838 29062 634074
rect 29146 633838 29382 634074
rect 37826 633218 38062 633454
rect 38146 633218 38382 633454
rect 37826 632898 38062 633134
rect 38146 632898 38382 633134
rect 46826 634158 47062 634394
rect 47146 634158 47382 634394
rect 46826 633838 47062 634074
rect 47146 633838 47382 634074
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 64826 634158 65062 634394
rect 65146 634158 65382 634394
rect 64826 633838 65062 634074
rect 65146 633838 65382 634074
rect 73826 633218 74062 633454
rect 74146 633218 74382 633454
rect 73826 632898 74062 633134
rect 74146 632898 74382 633134
rect 82826 634158 83062 634394
rect 83146 634158 83382 634394
rect 82826 633838 83062 634074
rect 83146 633838 83382 634074
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 100826 634158 101062 634394
rect 101146 634158 101382 634394
rect 100826 633838 101062 634074
rect 101146 633838 101382 634074
rect 109826 633218 110062 633454
rect 110146 633218 110382 633454
rect 109826 632898 110062 633134
rect 110146 632898 110382 633134
rect 118826 634158 119062 634394
rect 119146 634158 119382 634394
rect 118826 633838 119062 634074
rect 119146 633838 119382 634074
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 136826 634158 137062 634394
rect 137146 634158 137382 634394
rect 136826 633838 137062 634074
rect 137146 633838 137382 634074
rect 145826 633218 146062 633454
rect 146146 633218 146382 633454
rect 145826 632898 146062 633134
rect 146146 632898 146382 633134
rect 154826 634158 155062 634394
rect 155146 634158 155382 634394
rect 154826 633838 155062 634074
rect 155146 633838 155382 634074
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 172826 634158 173062 634394
rect 173146 634158 173382 634394
rect 172826 633838 173062 634074
rect 173146 633838 173382 634074
rect 181826 633218 182062 633454
rect 182146 633218 182382 633454
rect 181826 632898 182062 633134
rect 182146 632898 182382 633134
rect 190826 634158 191062 634394
rect 191146 634158 191382 634394
rect 190826 633838 191062 634074
rect 191146 633838 191382 634074
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 208826 634158 209062 634394
rect 209146 634158 209382 634394
rect 208826 633838 209062 634074
rect 209146 633838 209382 634074
rect 217826 633218 218062 633454
rect 218146 633218 218382 633454
rect 217826 632898 218062 633134
rect 218146 632898 218382 633134
rect 226826 634158 227062 634394
rect 227146 634158 227382 634394
rect 226826 633838 227062 634074
rect 227146 633838 227382 634074
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 244826 634158 245062 634394
rect 245146 634158 245382 634394
rect 244826 633838 245062 634074
rect 245146 633838 245382 634074
rect 253826 633218 254062 633454
rect 254146 633218 254382 633454
rect 253826 632898 254062 633134
rect 254146 632898 254382 633134
rect 262826 634158 263062 634394
rect 263146 634158 263382 634394
rect 262826 633838 263062 634074
rect 263146 633838 263382 634074
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 280826 634158 281062 634394
rect 281146 634158 281382 634394
rect 280826 633838 281062 634074
rect 281146 633838 281382 634074
rect 289826 633218 290062 633454
rect 290146 633218 290382 633454
rect 289826 632898 290062 633134
rect 290146 632898 290382 633134
rect 298826 634158 299062 634394
rect 299146 634158 299382 634394
rect 298826 633838 299062 634074
rect 299146 633838 299382 634074
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 316826 634158 317062 634394
rect 317146 634158 317382 634394
rect 316826 633838 317062 634074
rect 317146 633838 317382 634074
rect 325826 633218 326062 633454
rect 326146 633218 326382 633454
rect 325826 632898 326062 633134
rect 326146 632898 326382 633134
rect 334826 634158 335062 634394
rect 335146 634158 335382 634394
rect 334826 633838 335062 634074
rect 335146 633838 335382 634074
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 352826 634158 353062 634394
rect 353146 634158 353382 634394
rect 352826 633838 353062 634074
rect 353146 633838 353382 634074
rect 361826 633218 362062 633454
rect 362146 633218 362382 633454
rect 361826 632898 362062 633134
rect 362146 632898 362382 633134
rect 370826 634158 371062 634394
rect 371146 634158 371382 634394
rect 370826 633838 371062 634074
rect 371146 633838 371382 634074
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 388826 634158 389062 634394
rect 389146 634158 389382 634394
rect 388826 633838 389062 634074
rect 389146 633838 389382 634074
rect 397826 633218 398062 633454
rect 398146 633218 398382 633454
rect 397826 632898 398062 633134
rect 398146 632898 398382 633134
rect 406826 634158 407062 634394
rect 407146 634158 407382 634394
rect 406826 633838 407062 634074
rect 407146 633838 407382 634074
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 424826 634158 425062 634394
rect 425146 634158 425382 634394
rect 424826 633838 425062 634074
rect 425146 633838 425382 634074
rect 433826 633218 434062 633454
rect 434146 633218 434382 633454
rect 433826 632898 434062 633134
rect 434146 632898 434382 633134
rect 442826 634158 443062 634394
rect 443146 634158 443382 634394
rect 442826 633838 443062 634074
rect 443146 633838 443382 634074
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 460826 634158 461062 634394
rect 461146 634158 461382 634394
rect 460826 633838 461062 634074
rect 461146 633838 461382 634074
rect 469826 633218 470062 633454
rect 470146 633218 470382 633454
rect 469826 632898 470062 633134
rect 470146 632898 470382 633134
rect 478826 634158 479062 634394
rect 479146 634158 479382 634394
rect 478826 633838 479062 634074
rect 479146 633838 479382 634074
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 496826 634158 497062 634394
rect 497146 634158 497382 634394
rect 496826 633838 497062 634074
rect 497146 633838 497382 634074
rect 505826 633218 506062 633454
rect 506146 633218 506382 633454
rect 505826 632898 506062 633134
rect 506146 632898 506382 633134
rect 514826 634158 515062 634394
rect 515146 634158 515382 634394
rect 514826 633838 515062 634074
rect 515146 633838 515382 634074
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 532826 634158 533062 634394
rect 533146 634158 533382 634394
rect 532826 633838 533062 634074
rect 533146 633838 533382 634074
rect 541826 633218 542062 633454
rect 542146 633218 542382 633454
rect 541826 632898 542062 633134
rect 542146 632898 542382 633134
rect 550826 634158 551062 634394
rect 551146 634158 551382 634394
rect 550826 633838 551062 634074
rect 551146 633838 551382 634074
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 22916 624218 23152 624454
rect 22916 623898 23152 624134
rect 28847 624218 29083 624454
rect 28847 623898 29083 624134
rect 49916 624218 50152 624454
rect 49916 623898 50152 624134
rect 55847 624218 56083 624454
rect 55847 623898 56083 624134
rect 76916 624218 77152 624454
rect 76916 623898 77152 624134
rect 82847 624218 83083 624454
rect 82847 623898 83083 624134
rect 103916 624218 104152 624454
rect 103916 623898 104152 624134
rect 109847 624218 110083 624454
rect 109847 623898 110083 624134
rect 130916 624218 131152 624454
rect 130916 623898 131152 624134
rect 136847 624218 137083 624454
rect 136847 623898 137083 624134
rect 157916 624218 158152 624454
rect 157916 623898 158152 624134
rect 163847 624218 164083 624454
rect 163847 623898 164083 624134
rect 184916 624218 185152 624454
rect 184916 623898 185152 624134
rect 190847 624218 191083 624454
rect 190847 623898 191083 624134
rect 211916 624218 212152 624454
rect 211916 623898 212152 624134
rect 217847 624218 218083 624454
rect 217847 623898 218083 624134
rect 238916 624218 239152 624454
rect 238916 623898 239152 624134
rect 244847 624218 245083 624454
rect 244847 623898 245083 624134
rect 265916 624218 266152 624454
rect 265916 623898 266152 624134
rect 271847 624218 272083 624454
rect 271847 623898 272083 624134
rect 292916 624218 293152 624454
rect 292916 623898 293152 624134
rect 298847 624218 299083 624454
rect 298847 623898 299083 624134
rect 319916 624218 320152 624454
rect 319916 623898 320152 624134
rect 325847 624218 326083 624454
rect 325847 623898 326083 624134
rect 346916 624218 347152 624454
rect 346916 623898 347152 624134
rect 352847 624218 353083 624454
rect 352847 623898 353083 624134
rect 373916 624218 374152 624454
rect 373916 623898 374152 624134
rect 379847 624218 380083 624454
rect 379847 623898 380083 624134
rect 400916 624218 401152 624454
rect 400916 623898 401152 624134
rect 406847 624218 407083 624454
rect 406847 623898 407083 624134
rect 427916 624218 428152 624454
rect 427916 623898 428152 624134
rect 433847 624218 434083 624454
rect 433847 623898 434083 624134
rect 454916 624218 455152 624454
rect 454916 623898 455152 624134
rect 460847 624218 461083 624454
rect 460847 623898 461083 624134
rect 481916 624218 482152 624454
rect 481916 623898 482152 624134
rect 487847 624218 488083 624454
rect 487847 623898 488083 624134
rect 508916 624218 509152 624454
rect 508916 623898 509152 624134
rect 514847 624218 515083 624454
rect 514847 623898 515083 624134
rect 535916 624218 536152 624454
rect 535916 623898 536152 624134
rect 541847 624218 542083 624454
rect 541847 623898 542083 624134
rect 19952 615218 20188 615454
rect 19952 614898 20188 615134
rect 25882 615218 26118 615454
rect 25882 614898 26118 615134
rect 31813 615218 32049 615454
rect 31813 614898 32049 615134
rect 46952 615218 47188 615454
rect 46952 614898 47188 615134
rect 52882 615218 53118 615454
rect 52882 614898 53118 615134
rect 58813 615218 59049 615454
rect 58813 614898 59049 615134
rect 73952 615218 74188 615454
rect 73952 614898 74188 615134
rect 79882 615218 80118 615454
rect 79882 614898 80118 615134
rect 85813 615218 86049 615454
rect 85813 614898 86049 615134
rect 100952 615218 101188 615454
rect 100952 614898 101188 615134
rect 106882 615218 107118 615454
rect 106882 614898 107118 615134
rect 112813 615218 113049 615454
rect 112813 614898 113049 615134
rect 127952 615218 128188 615454
rect 127952 614898 128188 615134
rect 133882 615218 134118 615454
rect 133882 614898 134118 615134
rect 139813 615218 140049 615454
rect 139813 614898 140049 615134
rect 154952 615218 155188 615454
rect 154952 614898 155188 615134
rect 160882 615218 161118 615454
rect 160882 614898 161118 615134
rect 166813 615218 167049 615454
rect 166813 614898 167049 615134
rect 181952 615218 182188 615454
rect 181952 614898 182188 615134
rect 187882 615218 188118 615454
rect 187882 614898 188118 615134
rect 193813 615218 194049 615454
rect 193813 614898 194049 615134
rect 208952 615218 209188 615454
rect 208952 614898 209188 615134
rect 214882 615218 215118 615454
rect 214882 614898 215118 615134
rect 220813 615218 221049 615454
rect 220813 614898 221049 615134
rect 235952 615218 236188 615454
rect 235952 614898 236188 615134
rect 241882 615218 242118 615454
rect 241882 614898 242118 615134
rect 247813 615218 248049 615454
rect 247813 614898 248049 615134
rect 262952 615218 263188 615454
rect 262952 614898 263188 615134
rect 268882 615218 269118 615454
rect 268882 614898 269118 615134
rect 274813 615218 275049 615454
rect 274813 614898 275049 615134
rect 289952 615218 290188 615454
rect 289952 614898 290188 615134
rect 295882 615218 296118 615454
rect 295882 614898 296118 615134
rect 301813 615218 302049 615454
rect 301813 614898 302049 615134
rect 316952 615218 317188 615454
rect 316952 614898 317188 615134
rect 322882 615218 323118 615454
rect 322882 614898 323118 615134
rect 328813 615218 329049 615454
rect 328813 614898 329049 615134
rect 343952 615218 344188 615454
rect 343952 614898 344188 615134
rect 349882 615218 350118 615454
rect 349882 614898 350118 615134
rect 355813 615218 356049 615454
rect 355813 614898 356049 615134
rect 370952 615218 371188 615454
rect 370952 614898 371188 615134
rect 376882 615218 377118 615454
rect 376882 614898 377118 615134
rect 382813 615218 383049 615454
rect 382813 614898 383049 615134
rect 397952 615218 398188 615454
rect 397952 614898 398188 615134
rect 403882 615218 404118 615454
rect 403882 614898 404118 615134
rect 409813 615218 410049 615454
rect 409813 614898 410049 615134
rect 424952 615218 425188 615454
rect 424952 614898 425188 615134
rect 430882 615218 431118 615454
rect 430882 614898 431118 615134
rect 436813 615218 437049 615454
rect 436813 614898 437049 615134
rect 451952 615218 452188 615454
rect 451952 614898 452188 615134
rect 457882 615218 458118 615454
rect 457882 614898 458118 615134
rect 463813 615218 464049 615454
rect 463813 614898 464049 615134
rect 478952 615218 479188 615454
rect 478952 614898 479188 615134
rect 484882 615218 485118 615454
rect 484882 614898 485118 615134
rect 490813 615218 491049 615454
rect 490813 614898 491049 615134
rect 505952 615218 506188 615454
rect 505952 614898 506188 615134
rect 511882 615218 512118 615454
rect 511882 614898 512118 615134
rect 517813 615218 518049 615454
rect 517813 614898 518049 615134
rect 532952 615218 533188 615454
rect 532952 614898 533188 615134
rect 538882 615218 539118 615454
rect 538882 614898 539118 615134
rect 544813 615218 545049 615454
rect 544813 614898 545049 615134
rect 559826 615218 560062 615454
rect 560146 615218 560382 615454
rect 559826 614898 560062 615134
rect 560146 614898 560382 615134
rect 10826 606218 11062 606454
rect 11146 606218 11382 606454
rect 10826 605898 11062 606134
rect 11146 605898 11382 606134
rect 19826 607158 20062 607394
rect 20146 607158 20382 607394
rect 19826 606838 20062 607074
rect 20146 606838 20382 607074
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 37826 607158 38062 607394
rect 38146 607158 38382 607394
rect 37826 606838 38062 607074
rect 38146 606838 38382 607074
rect 46826 606218 47062 606454
rect 47146 606218 47382 606454
rect 46826 605898 47062 606134
rect 47146 605898 47382 606134
rect 55826 607158 56062 607394
rect 56146 607158 56382 607394
rect 55826 606838 56062 607074
rect 56146 606838 56382 607074
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 73826 607158 74062 607394
rect 74146 607158 74382 607394
rect 73826 606838 74062 607074
rect 74146 606838 74382 607074
rect 82826 606218 83062 606454
rect 83146 606218 83382 606454
rect 82826 605898 83062 606134
rect 83146 605898 83382 606134
rect 91826 607158 92062 607394
rect 92146 607158 92382 607394
rect 91826 606838 92062 607074
rect 92146 606838 92382 607074
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 109826 607158 110062 607394
rect 110146 607158 110382 607394
rect 109826 606838 110062 607074
rect 110146 606838 110382 607074
rect 118826 606218 119062 606454
rect 119146 606218 119382 606454
rect 118826 605898 119062 606134
rect 119146 605898 119382 606134
rect 127826 607158 128062 607394
rect 128146 607158 128382 607394
rect 127826 606838 128062 607074
rect 128146 606838 128382 607074
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 145826 607158 146062 607394
rect 146146 607158 146382 607394
rect 145826 606838 146062 607074
rect 146146 606838 146382 607074
rect 154826 606218 155062 606454
rect 155146 606218 155382 606454
rect 154826 605898 155062 606134
rect 155146 605898 155382 606134
rect 163826 607158 164062 607394
rect 164146 607158 164382 607394
rect 163826 606838 164062 607074
rect 164146 606838 164382 607074
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 181826 607158 182062 607394
rect 182146 607158 182382 607394
rect 181826 606838 182062 607074
rect 182146 606838 182382 607074
rect 190826 606218 191062 606454
rect 191146 606218 191382 606454
rect 190826 605898 191062 606134
rect 191146 605898 191382 606134
rect 199826 607158 200062 607394
rect 200146 607158 200382 607394
rect 199826 606838 200062 607074
rect 200146 606838 200382 607074
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 217826 607158 218062 607394
rect 218146 607158 218382 607394
rect 217826 606838 218062 607074
rect 218146 606838 218382 607074
rect 226826 606218 227062 606454
rect 227146 606218 227382 606454
rect 226826 605898 227062 606134
rect 227146 605898 227382 606134
rect 235826 607158 236062 607394
rect 236146 607158 236382 607394
rect 235826 606838 236062 607074
rect 236146 606838 236382 607074
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 253826 607158 254062 607394
rect 254146 607158 254382 607394
rect 253826 606838 254062 607074
rect 254146 606838 254382 607074
rect 262826 606218 263062 606454
rect 263146 606218 263382 606454
rect 262826 605898 263062 606134
rect 263146 605898 263382 606134
rect 271826 607158 272062 607394
rect 272146 607158 272382 607394
rect 271826 606838 272062 607074
rect 272146 606838 272382 607074
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 289826 607158 290062 607394
rect 290146 607158 290382 607394
rect 289826 606838 290062 607074
rect 290146 606838 290382 607074
rect 298826 606218 299062 606454
rect 299146 606218 299382 606454
rect 298826 605898 299062 606134
rect 299146 605898 299382 606134
rect 307826 607158 308062 607394
rect 308146 607158 308382 607394
rect 307826 606838 308062 607074
rect 308146 606838 308382 607074
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 325826 607158 326062 607394
rect 326146 607158 326382 607394
rect 325826 606838 326062 607074
rect 326146 606838 326382 607074
rect 334826 606218 335062 606454
rect 335146 606218 335382 606454
rect 334826 605898 335062 606134
rect 335146 605898 335382 606134
rect 343826 607158 344062 607394
rect 344146 607158 344382 607394
rect 343826 606838 344062 607074
rect 344146 606838 344382 607074
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 361826 607158 362062 607394
rect 362146 607158 362382 607394
rect 361826 606838 362062 607074
rect 362146 606838 362382 607074
rect 370826 606218 371062 606454
rect 371146 606218 371382 606454
rect 370826 605898 371062 606134
rect 371146 605898 371382 606134
rect 379826 607158 380062 607394
rect 380146 607158 380382 607394
rect 379826 606838 380062 607074
rect 380146 606838 380382 607074
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 397826 607158 398062 607394
rect 398146 607158 398382 607394
rect 397826 606838 398062 607074
rect 398146 606838 398382 607074
rect 406826 606218 407062 606454
rect 407146 606218 407382 606454
rect 406826 605898 407062 606134
rect 407146 605898 407382 606134
rect 415826 607158 416062 607394
rect 416146 607158 416382 607394
rect 415826 606838 416062 607074
rect 416146 606838 416382 607074
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 433826 607158 434062 607394
rect 434146 607158 434382 607394
rect 433826 606838 434062 607074
rect 434146 606838 434382 607074
rect 442826 606218 443062 606454
rect 443146 606218 443382 606454
rect 442826 605898 443062 606134
rect 443146 605898 443382 606134
rect 451826 607158 452062 607394
rect 452146 607158 452382 607394
rect 451826 606838 452062 607074
rect 452146 606838 452382 607074
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 469826 607158 470062 607394
rect 470146 607158 470382 607394
rect 469826 606838 470062 607074
rect 470146 606838 470382 607074
rect 478826 606218 479062 606454
rect 479146 606218 479382 606454
rect 478826 605898 479062 606134
rect 479146 605898 479382 606134
rect 487826 607158 488062 607394
rect 488146 607158 488382 607394
rect 487826 606838 488062 607074
rect 488146 606838 488382 607074
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 505826 607158 506062 607394
rect 506146 607158 506382 607394
rect 505826 606838 506062 607074
rect 506146 606838 506382 607074
rect 514826 606218 515062 606454
rect 515146 606218 515382 606454
rect 514826 605898 515062 606134
rect 515146 605898 515382 606134
rect 523826 607158 524062 607394
rect 524146 607158 524382 607394
rect 523826 606838 524062 607074
rect 524146 606838 524382 607074
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 541826 607158 542062 607394
rect 542146 607158 542382 607394
rect 541826 606838 542062 607074
rect 542146 606838 542382 607074
rect 550826 606218 551062 606454
rect 551146 606218 551382 606454
rect 550826 605898 551062 606134
rect 551146 605898 551382 606134
rect 19952 597218 20188 597454
rect 19952 596898 20188 597134
rect 25882 597218 26118 597454
rect 25882 596898 26118 597134
rect 31813 597218 32049 597454
rect 31813 596898 32049 597134
rect 46952 597218 47188 597454
rect 46952 596898 47188 597134
rect 52882 597218 53118 597454
rect 52882 596898 53118 597134
rect 58813 597218 59049 597454
rect 58813 596898 59049 597134
rect 73952 597218 74188 597454
rect 73952 596898 74188 597134
rect 79882 597218 80118 597454
rect 79882 596898 80118 597134
rect 85813 597218 86049 597454
rect 85813 596898 86049 597134
rect 100952 597218 101188 597454
rect 100952 596898 101188 597134
rect 106882 597218 107118 597454
rect 106882 596898 107118 597134
rect 112813 597218 113049 597454
rect 112813 596898 113049 597134
rect 127952 597218 128188 597454
rect 127952 596898 128188 597134
rect 133882 597218 134118 597454
rect 133882 596898 134118 597134
rect 139813 597218 140049 597454
rect 139813 596898 140049 597134
rect 154952 597218 155188 597454
rect 154952 596898 155188 597134
rect 160882 597218 161118 597454
rect 160882 596898 161118 597134
rect 166813 597218 167049 597454
rect 166813 596898 167049 597134
rect 181952 597218 182188 597454
rect 181952 596898 182188 597134
rect 187882 597218 188118 597454
rect 187882 596898 188118 597134
rect 193813 597218 194049 597454
rect 193813 596898 194049 597134
rect 208952 597218 209188 597454
rect 208952 596898 209188 597134
rect 214882 597218 215118 597454
rect 214882 596898 215118 597134
rect 220813 597218 221049 597454
rect 220813 596898 221049 597134
rect 235952 597218 236188 597454
rect 235952 596898 236188 597134
rect 241882 597218 242118 597454
rect 241882 596898 242118 597134
rect 247813 597218 248049 597454
rect 247813 596898 248049 597134
rect 262952 597218 263188 597454
rect 262952 596898 263188 597134
rect 268882 597218 269118 597454
rect 268882 596898 269118 597134
rect 274813 597218 275049 597454
rect 274813 596898 275049 597134
rect 289952 597218 290188 597454
rect 289952 596898 290188 597134
rect 295882 597218 296118 597454
rect 295882 596898 296118 597134
rect 301813 597218 302049 597454
rect 301813 596898 302049 597134
rect 316952 597218 317188 597454
rect 316952 596898 317188 597134
rect 322882 597218 323118 597454
rect 322882 596898 323118 597134
rect 328813 597218 329049 597454
rect 328813 596898 329049 597134
rect 343952 597218 344188 597454
rect 343952 596898 344188 597134
rect 349882 597218 350118 597454
rect 349882 596898 350118 597134
rect 355813 597218 356049 597454
rect 355813 596898 356049 597134
rect 370952 597218 371188 597454
rect 370952 596898 371188 597134
rect 376882 597218 377118 597454
rect 376882 596898 377118 597134
rect 382813 597218 383049 597454
rect 382813 596898 383049 597134
rect 397952 597218 398188 597454
rect 397952 596898 398188 597134
rect 403882 597218 404118 597454
rect 403882 596898 404118 597134
rect 409813 597218 410049 597454
rect 409813 596898 410049 597134
rect 424952 597218 425188 597454
rect 424952 596898 425188 597134
rect 430882 597218 431118 597454
rect 430882 596898 431118 597134
rect 436813 597218 437049 597454
rect 436813 596898 437049 597134
rect 451952 597218 452188 597454
rect 451952 596898 452188 597134
rect 457882 597218 458118 597454
rect 457882 596898 458118 597134
rect 463813 597218 464049 597454
rect 463813 596898 464049 597134
rect 478952 597218 479188 597454
rect 478952 596898 479188 597134
rect 484882 597218 485118 597454
rect 484882 596898 485118 597134
rect 490813 597218 491049 597454
rect 490813 596898 491049 597134
rect 505952 597218 506188 597454
rect 505952 596898 506188 597134
rect 511882 597218 512118 597454
rect 511882 596898 512118 597134
rect 517813 597218 518049 597454
rect 517813 596898 518049 597134
rect 532952 597218 533188 597454
rect 532952 596898 533188 597134
rect 538882 597218 539118 597454
rect 538882 596898 539118 597134
rect 544813 597218 545049 597454
rect 544813 596898 545049 597134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 22916 588218 23152 588454
rect 22916 587898 23152 588134
rect 28847 588218 29083 588454
rect 28847 587898 29083 588134
rect 49916 588218 50152 588454
rect 49916 587898 50152 588134
rect 55847 588218 56083 588454
rect 55847 587898 56083 588134
rect 76916 588218 77152 588454
rect 76916 587898 77152 588134
rect 82847 588218 83083 588454
rect 82847 587898 83083 588134
rect 103916 588218 104152 588454
rect 103916 587898 104152 588134
rect 109847 588218 110083 588454
rect 109847 587898 110083 588134
rect 130916 588218 131152 588454
rect 130916 587898 131152 588134
rect 136847 588218 137083 588454
rect 136847 587898 137083 588134
rect 157916 588218 158152 588454
rect 157916 587898 158152 588134
rect 163847 588218 164083 588454
rect 163847 587898 164083 588134
rect 184916 588218 185152 588454
rect 184916 587898 185152 588134
rect 190847 588218 191083 588454
rect 190847 587898 191083 588134
rect 211916 588218 212152 588454
rect 211916 587898 212152 588134
rect 217847 588218 218083 588454
rect 217847 587898 218083 588134
rect 238916 588218 239152 588454
rect 238916 587898 239152 588134
rect 244847 588218 245083 588454
rect 244847 587898 245083 588134
rect 265916 588218 266152 588454
rect 265916 587898 266152 588134
rect 271847 588218 272083 588454
rect 271847 587898 272083 588134
rect 292916 588218 293152 588454
rect 292916 587898 293152 588134
rect 298847 588218 299083 588454
rect 298847 587898 299083 588134
rect 319916 588218 320152 588454
rect 319916 587898 320152 588134
rect 325847 588218 326083 588454
rect 325847 587898 326083 588134
rect 346916 588218 347152 588454
rect 346916 587898 347152 588134
rect 352847 588218 353083 588454
rect 352847 587898 353083 588134
rect 373916 588218 374152 588454
rect 373916 587898 374152 588134
rect 379847 588218 380083 588454
rect 379847 587898 380083 588134
rect 400916 588218 401152 588454
rect 400916 587898 401152 588134
rect 406847 588218 407083 588454
rect 406847 587898 407083 588134
rect 427916 588218 428152 588454
rect 427916 587898 428152 588134
rect 433847 588218 434083 588454
rect 433847 587898 434083 588134
rect 454916 588218 455152 588454
rect 454916 587898 455152 588134
rect 460847 588218 461083 588454
rect 460847 587898 461083 588134
rect 481916 588218 482152 588454
rect 481916 587898 482152 588134
rect 487847 588218 488083 588454
rect 487847 587898 488083 588134
rect 508916 588218 509152 588454
rect 508916 587898 509152 588134
rect 514847 588218 515083 588454
rect 514847 587898 515083 588134
rect 535916 588218 536152 588454
rect 535916 587898 536152 588134
rect 541847 588218 542083 588454
rect 541847 587898 542083 588134
rect 19826 579218 20062 579454
rect 20146 579218 20382 579454
rect 19826 578898 20062 579134
rect 20146 578898 20382 579134
rect 28826 580158 29062 580394
rect 29146 580158 29382 580394
rect 28826 579838 29062 580074
rect 29146 579838 29382 580074
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 46826 580158 47062 580394
rect 47146 580158 47382 580394
rect 46826 579838 47062 580074
rect 47146 579838 47382 580074
rect 55826 579218 56062 579454
rect 56146 579218 56382 579454
rect 55826 578898 56062 579134
rect 56146 578898 56382 579134
rect 64826 580158 65062 580394
rect 65146 580158 65382 580394
rect 64826 579838 65062 580074
rect 65146 579838 65382 580074
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 82826 580158 83062 580394
rect 83146 580158 83382 580394
rect 82826 579838 83062 580074
rect 83146 579838 83382 580074
rect 91826 579218 92062 579454
rect 92146 579218 92382 579454
rect 91826 578898 92062 579134
rect 92146 578898 92382 579134
rect 100826 580158 101062 580394
rect 101146 580158 101382 580394
rect 100826 579838 101062 580074
rect 101146 579838 101382 580074
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 118826 580158 119062 580394
rect 119146 580158 119382 580394
rect 118826 579838 119062 580074
rect 119146 579838 119382 580074
rect 127826 579218 128062 579454
rect 128146 579218 128382 579454
rect 127826 578898 128062 579134
rect 128146 578898 128382 579134
rect 136826 580158 137062 580394
rect 137146 580158 137382 580394
rect 136826 579838 137062 580074
rect 137146 579838 137382 580074
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 154826 580158 155062 580394
rect 155146 580158 155382 580394
rect 154826 579838 155062 580074
rect 155146 579838 155382 580074
rect 163826 579218 164062 579454
rect 164146 579218 164382 579454
rect 163826 578898 164062 579134
rect 164146 578898 164382 579134
rect 172826 580158 173062 580394
rect 173146 580158 173382 580394
rect 172826 579838 173062 580074
rect 173146 579838 173382 580074
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 190826 580158 191062 580394
rect 191146 580158 191382 580394
rect 190826 579838 191062 580074
rect 191146 579838 191382 580074
rect 199826 579218 200062 579454
rect 200146 579218 200382 579454
rect 199826 578898 200062 579134
rect 200146 578898 200382 579134
rect 208826 580158 209062 580394
rect 209146 580158 209382 580394
rect 208826 579838 209062 580074
rect 209146 579838 209382 580074
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 226826 580158 227062 580394
rect 227146 580158 227382 580394
rect 226826 579838 227062 580074
rect 227146 579838 227382 580074
rect 235826 579218 236062 579454
rect 236146 579218 236382 579454
rect 235826 578898 236062 579134
rect 236146 578898 236382 579134
rect 244826 580158 245062 580394
rect 245146 580158 245382 580394
rect 244826 579838 245062 580074
rect 245146 579838 245382 580074
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 262826 580158 263062 580394
rect 263146 580158 263382 580394
rect 262826 579838 263062 580074
rect 263146 579838 263382 580074
rect 271826 579218 272062 579454
rect 272146 579218 272382 579454
rect 271826 578898 272062 579134
rect 272146 578898 272382 579134
rect 280826 580158 281062 580394
rect 281146 580158 281382 580394
rect 280826 579838 281062 580074
rect 281146 579838 281382 580074
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 298826 580158 299062 580394
rect 299146 580158 299382 580394
rect 298826 579838 299062 580074
rect 299146 579838 299382 580074
rect 307826 579218 308062 579454
rect 308146 579218 308382 579454
rect 307826 578898 308062 579134
rect 308146 578898 308382 579134
rect 316826 580158 317062 580394
rect 317146 580158 317382 580394
rect 316826 579838 317062 580074
rect 317146 579838 317382 580074
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 334826 580158 335062 580394
rect 335146 580158 335382 580394
rect 334826 579838 335062 580074
rect 335146 579838 335382 580074
rect 343826 579218 344062 579454
rect 344146 579218 344382 579454
rect 343826 578898 344062 579134
rect 344146 578898 344382 579134
rect 352826 580158 353062 580394
rect 353146 580158 353382 580394
rect 352826 579838 353062 580074
rect 353146 579838 353382 580074
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 370826 580158 371062 580394
rect 371146 580158 371382 580394
rect 370826 579838 371062 580074
rect 371146 579838 371382 580074
rect 379826 579218 380062 579454
rect 380146 579218 380382 579454
rect 379826 578898 380062 579134
rect 380146 578898 380382 579134
rect 388826 580158 389062 580394
rect 389146 580158 389382 580394
rect 388826 579838 389062 580074
rect 389146 579838 389382 580074
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 406826 580158 407062 580394
rect 407146 580158 407382 580394
rect 406826 579838 407062 580074
rect 407146 579838 407382 580074
rect 415826 579218 416062 579454
rect 416146 579218 416382 579454
rect 415826 578898 416062 579134
rect 416146 578898 416382 579134
rect 424826 580158 425062 580394
rect 425146 580158 425382 580394
rect 424826 579838 425062 580074
rect 425146 579838 425382 580074
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 442826 580158 443062 580394
rect 443146 580158 443382 580394
rect 442826 579838 443062 580074
rect 443146 579838 443382 580074
rect 451826 579218 452062 579454
rect 452146 579218 452382 579454
rect 451826 578898 452062 579134
rect 452146 578898 452382 579134
rect 460826 580158 461062 580394
rect 461146 580158 461382 580394
rect 460826 579838 461062 580074
rect 461146 579838 461382 580074
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 478826 580158 479062 580394
rect 479146 580158 479382 580394
rect 478826 579838 479062 580074
rect 479146 579838 479382 580074
rect 487826 579218 488062 579454
rect 488146 579218 488382 579454
rect 487826 578898 488062 579134
rect 488146 578898 488382 579134
rect 496826 580158 497062 580394
rect 497146 580158 497382 580394
rect 496826 579838 497062 580074
rect 497146 579838 497382 580074
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 514826 580158 515062 580394
rect 515146 580158 515382 580394
rect 514826 579838 515062 580074
rect 515146 579838 515382 580074
rect 523826 579218 524062 579454
rect 524146 579218 524382 579454
rect 523826 578898 524062 579134
rect 524146 578898 524382 579134
rect 532826 580158 533062 580394
rect 533146 580158 533382 580394
rect 532826 579838 533062 580074
rect 533146 579838 533382 580074
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 550826 580158 551062 580394
rect 551146 580158 551382 580394
rect 550826 579838 551062 580074
rect 551146 579838 551382 580074
rect 559826 579218 560062 579454
rect 560146 579218 560382 579454
rect 559826 578898 560062 579134
rect 560146 578898 560382 579134
rect 10826 570218 11062 570454
rect 11146 570218 11382 570454
rect 10826 569898 11062 570134
rect 11146 569898 11382 570134
rect 22916 570218 23152 570454
rect 22916 569898 23152 570134
rect 28847 570218 29083 570454
rect 28847 569898 29083 570134
rect 49916 570218 50152 570454
rect 49916 569898 50152 570134
rect 55847 570218 56083 570454
rect 55847 569898 56083 570134
rect 76916 570218 77152 570454
rect 76916 569898 77152 570134
rect 82847 570218 83083 570454
rect 82847 569898 83083 570134
rect 103916 570218 104152 570454
rect 103916 569898 104152 570134
rect 109847 570218 110083 570454
rect 109847 569898 110083 570134
rect 130916 570218 131152 570454
rect 130916 569898 131152 570134
rect 136847 570218 137083 570454
rect 136847 569898 137083 570134
rect 157916 570218 158152 570454
rect 157916 569898 158152 570134
rect 163847 570218 164083 570454
rect 163847 569898 164083 570134
rect 184916 570218 185152 570454
rect 184916 569898 185152 570134
rect 190847 570218 191083 570454
rect 190847 569898 191083 570134
rect 211916 570218 212152 570454
rect 211916 569898 212152 570134
rect 217847 570218 218083 570454
rect 217847 569898 218083 570134
rect 238916 570218 239152 570454
rect 238916 569898 239152 570134
rect 244847 570218 245083 570454
rect 244847 569898 245083 570134
rect 265916 570218 266152 570454
rect 265916 569898 266152 570134
rect 271847 570218 272083 570454
rect 271847 569898 272083 570134
rect 292916 570218 293152 570454
rect 292916 569898 293152 570134
rect 298847 570218 299083 570454
rect 298847 569898 299083 570134
rect 319916 570218 320152 570454
rect 319916 569898 320152 570134
rect 325847 570218 326083 570454
rect 325847 569898 326083 570134
rect 346916 570218 347152 570454
rect 346916 569898 347152 570134
rect 352847 570218 353083 570454
rect 352847 569898 353083 570134
rect 373916 570218 374152 570454
rect 373916 569898 374152 570134
rect 379847 570218 380083 570454
rect 379847 569898 380083 570134
rect 400916 570218 401152 570454
rect 400916 569898 401152 570134
rect 406847 570218 407083 570454
rect 406847 569898 407083 570134
rect 427916 570218 428152 570454
rect 427916 569898 428152 570134
rect 433847 570218 434083 570454
rect 433847 569898 434083 570134
rect 454916 570218 455152 570454
rect 454916 569898 455152 570134
rect 460847 570218 461083 570454
rect 460847 569898 461083 570134
rect 481916 570218 482152 570454
rect 481916 569898 482152 570134
rect 487847 570218 488083 570454
rect 487847 569898 488083 570134
rect 508916 570218 509152 570454
rect 508916 569898 509152 570134
rect 514847 570218 515083 570454
rect 514847 569898 515083 570134
rect 535916 570218 536152 570454
rect 535916 569898 536152 570134
rect 541847 570218 542083 570454
rect 541847 569898 542083 570134
rect 19952 561218 20188 561454
rect 19952 560898 20188 561134
rect 25882 561218 26118 561454
rect 25882 560898 26118 561134
rect 31813 561218 32049 561454
rect 31813 560898 32049 561134
rect 46952 561218 47188 561454
rect 46952 560898 47188 561134
rect 52882 561218 53118 561454
rect 52882 560898 53118 561134
rect 58813 561218 59049 561454
rect 58813 560898 59049 561134
rect 73952 561218 74188 561454
rect 73952 560898 74188 561134
rect 79882 561218 80118 561454
rect 79882 560898 80118 561134
rect 85813 561218 86049 561454
rect 85813 560898 86049 561134
rect 100952 561218 101188 561454
rect 100952 560898 101188 561134
rect 106882 561218 107118 561454
rect 106882 560898 107118 561134
rect 112813 561218 113049 561454
rect 112813 560898 113049 561134
rect 127952 561218 128188 561454
rect 127952 560898 128188 561134
rect 133882 561218 134118 561454
rect 133882 560898 134118 561134
rect 139813 561218 140049 561454
rect 139813 560898 140049 561134
rect 154952 561218 155188 561454
rect 154952 560898 155188 561134
rect 160882 561218 161118 561454
rect 160882 560898 161118 561134
rect 166813 561218 167049 561454
rect 166813 560898 167049 561134
rect 181952 561218 182188 561454
rect 181952 560898 182188 561134
rect 187882 561218 188118 561454
rect 187882 560898 188118 561134
rect 193813 561218 194049 561454
rect 193813 560898 194049 561134
rect 208952 561218 209188 561454
rect 208952 560898 209188 561134
rect 214882 561218 215118 561454
rect 214882 560898 215118 561134
rect 220813 561218 221049 561454
rect 220813 560898 221049 561134
rect 235952 561218 236188 561454
rect 235952 560898 236188 561134
rect 241882 561218 242118 561454
rect 241882 560898 242118 561134
rect 247813 561218 248049 561454
rect 247813 560898 248049 561134
rect 262952 561218 263188 561454
rect 262952 560898 263188 561134
rect 268882 561218 269118 561454
rect 268882 560898 269118 561134
rect 274813 561218 275049 561454
rect 274813 560898 275049 561134
rect 289952 561218 290188 561454
rect 289952 560898 290188 561134
rect 295882 561218 296118 561454
rect 295882 560898 296118 561134
rect 301813 561218 302049 561454
rect 301813 560898 302049 561134
rect 316952 561218 317188 561454
rect 316952 560898 317188 561134
rect 322882 561218 323118 561454
rect 322882 560898 323118 561134
rect 328813 561218 329049 561454
rect 328813 560898 329049 561134
rect 343952 561218 344188 561454
rect 343952 560898 344188 561134
rect 349882 561218 350118 561454
rect 349882 560898 350118 561134
rect 355813 561218 356049 561454
rect 355813 560898 356049 561134
rect 370952 561218 371188 561454
rect 370952 560898 371188 561134
rect 376882 561218 377118 561454
rect 376882 560898 377118 561134
rect 382813 561218 383049 561454
rect 382813 560898 383049 561134
rect 397952 561218 398188 561454
rect 397952 560898 398188 561134
rect 403882 561218 404118 561454
rect 403882 560898 404118 561134
rect 409813 561218 410049 561454
rect 409813 560898 410049 561134
rect 424952 561218 425188 561454
rect 424952 560898 425188 561134
rect 430882 561218 431118 561454
rect 430882 560898 431118 561134
rect 436813 561218 437049 561454
rect 436813 560898 437049 561134
rect 451952 561218 452188 561454
rect 451952 560898 452188 561134
rect 457882 561218 458118 561454
rect 457882 560898 458118 561134
rect 463813 561218 464049 561454
rect 463813 560898 464049 561134
rect 478952 561218 479188 561454
rect 478952 560898 479188 561134
rect 484882 561218 485118 561454
rect 484882 560898 485118 561134
rect 490813 561218 491049 561454
rect 490813 560898 491049 561134
rect 505952 561218 506188 561454
rect 505952 560898 506188 561134
rect 511882 561218 512118 561454
rect 511882 560898 512118 561134
rect 517813 561218 518049 561454
rect 517813 560898 518049 561134
rect 532952 561218 533188 561454
rect 532952 560898 533188 561134
rect 538882 561218 539118 561454
rect 538882 560898 539118 561134
rect 544813 561218 545049 561454
rect 544813 560898 545049 561134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 19826 553158 20062 553394
rect 20146 553158 20382 553394
rect 19826 552838 20062 553074
rect 20146 552838 20382 553074
rect 28826 552218 29062 552454
rect 29146 552218 29382 552454
rect 28826 551898 29062 552134
rect 29146 551898 29382 552134
rect 37826 553158 38062 553394
rect 38146 553158 38382 553394
rect 37826 552838 38062 553074
rect 38146 552838 38382 553074
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 55826 553158 56062 553394
rect 56146 553158 56382 553394
rect 55826 552838 56062 553074
rect 56146 552838 56382 553074
rect 64826 552218 65062 552454
rect 65146 552218 65382 552454
rect 64826 551898 65062 552134
rect 65146 551898 65382 552134
rect 73826 553158 74062 553394
rect 74146 553158 74382 553394
rect 73826 552838 74062 553074
rect 74146 552838 74382 553074
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 91826 553158 92062 553394
rect 92146 553158 92382 553394
rect 91826 552838 92062 553074
rect 92146 552838 92382 553074
rect 100826 552218 101062 552454
rect 101146 552218 101382 552454
rect 100826 551898 101062 552134
rect 101146 551898 101382 552134
rect 109826 553158 110062 553394
rect 110146 553158 110382 553394
rect 109826 552838 110062 553074
rect 110146 552838 110382 553074
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 127826 553158 128062 553394
rect 128146 553158 128382 553394
rect 127826 552838 128062 553074
rect 128146 552838 128382 553074
rect 136826 552218 137062 552454
rect 137146 552218 137382 552454
rect 136826 551898 137062 552134
rect 137146 551898 137382 552134
rect 145826 553158 146062 553394
rect 146146 553158 146382 553394
rect 145826 552838 146062 553074
rect 146146 552838 146382 553074
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 163826 553158 164062 553394
rect 164146 553158 164382 553394
rect 163826 552838 164062 553074
rect 164146 552838 164382 553074
rect 172826 552218 173062 552454
rect 173146 552218 173382 552454
rect 172826 551898 173062 552134
rect 173146 551898 173382 552134
rect 181826 553158 182062 553394
rect 182146 553158 182382 553394
rect 181826 552838 182062 553074
rect 182146 552838 182382 553074
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 199826 553158 200062 553394
rect 200146 553158 200382 553394
rect 199826 552838 200062 553074
rect 200146 552838 200382 553074
rect 208826 552218 209062 552454
rect 209146 552218 209382 552454
rect 208826 551898 209062 552134
rect 209146 551898 209382 552134
rect 217826 553158 218062 553394
rect 218146 553158 218382 553394
rect 217826 552838 218062 553074
rect 218146 552838 218382 553074
rect 226826 552218 227062 552454
rect 227146 552218 227382 552454
rect 226826 551898 227062 552134
rect 227146 551898 227382 552134
rect 235826 553158 236062 553394
rect 236146 553158 236382 553394
rect 235826 552838 236062 553074
rect 236146 552838 236382 553074
rect 244826 552218 245062 552454
rect 245146 552218 245382 552454
rect 244826 551898 245062 552134
rect 245146 551898 245382 552134
rect 253826 553158 254062 553394
rect 254146 553158 254382 553394
rect 253826 552838 254062 553074
rect 254146 552838 254382 553074
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 271826 553158 272062 553394
rect 272146 553158 272382 553394
rect 271826 552838 272062 553074
rect 272146 552838 272382 553074
rect 280826 552218 281062 552454
rect 281146 552218 281382 552454
rect 280826 551898 281062 552134
rect 281146 551898 281382 552134
rect 289826 553158 290062 553394
rect 290146 553158 290382 553394
rect 289826 552838 290062 553074
rect 290146 552838 290382 553074
rect 298826 552218 299062 552454
rect 299146 552218 299382 552454
rect 298826 551898 299062 552134
rect 299146 551898 299382 552134
rect 307826 553158 308062 553394
rect 308146 553158 308382 553394
rect 307826 552838 308062 553074
rect 308146 552838 308382 553074
rect 316826 552218 317062 552454
rect 317146 552218 317382 552454
rect 316826 551898 317062 552134
rect 317146 551898 317382 552134
rect 325826 553158 326062 553394
rect 326146 553158 326382 553394
rect 325826 552838 326062 553074
rect 326146 552838 326382 553074
rect 334826 552218 335062 552454
rect 335146 552218 335382 552454
rect 334826 551898 335062 552134
rect 335146 551898 335382 552134
rect 343826 553158 344062 553394
rect 344146 553158 344382 553394
rect 343826 552838 344062 553074
rect 344146 552838 344382 553074
rect 352826 552218 353062 552454
rect 353146 552218 353382 552454
rect 352826 551898 353062 552134
rect 353146 551898 353382 552134
rect 361826 553158 362062 553394
rect 362146 553158 362382 553394
rect 361826 552838 362062 553074
rect 362146 552838 362382 553074
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 379826 553158 380062 553394
rect 380146 553158 380382 553394
rect 379826 552838 380062 553074
rect 380146 552838 380382 553074
rect 388826 552218 389062 552454
rect 389146 552218 389382 552454
rect 388826 551898 389062 552134
rect 389146 551898 389382 552134
rect 397826 553158 398062 553394
rect 398146 553158 398382 553394
rect 397826 552838 398062 553074
rect 398146 552838 398382 553074
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 415826 553158 416062 553394
rect 416146 553158 416382 553394
rect 415826 552838 416062 553074
rect 416146 552838 416382 553074
rect 424826 552218 425062 552454
rect 425146 552218 425382 552454
rect 424826 551898 425062 552134
rect 425146 551898 425382 552134
rect 433826 553158 434062 553394
rect 434146 553158 434382 553394
rect 433826 552838 434062 553074
rect 434146 552838 434382 553074
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 451826 553158 452062 553394
rect 452146 553158 452382 553394
rect 451826 552838 452062 553074
rect 452146 552838 452382 553074
rect 460826 552218 461062 552454
rect 461146 552218 461382 552454
rect 460826 551898 461062 552134
rect 461146 551898 461382 552134
rect 469826 553158 470062 553394
rect 470146 553158 470382 553394
rect 469826 552838 470062 553074
rect 470146 552838 470382 553074
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 487826 553158 488062 553394
rect 488146 553158 488382 553394
rect 487826 552838 488062 553074
rect 488146 552838 488382 553074
rect 496826 552218 497062 552454
rect 497146 552218 497382 552454
rect 496826 551898 497062 552134
rect 497146 551898 497382 552134
rect 505826 553158 506062 553394
rect 506146 553158 506382 553394
rect 505826 552838 506062 553074
rect 506146 552838 506382 553074
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 523826 553158 524062 553394
rect 524146 553158 524382 553394
rect 523826 552838 524062 553074
rect 524146 552838 524382 553074
rect 532826 552218 533062 552454
rect 533146 552218 533382 552454
rect 532826 551898 533062 552134
rect 533146 551898 533382 552134
rect 541826 553158 542062 553394
rect 542146 553158 542382 553394
rect 541826 552838 542062 553074
rect 542146 552838 542382 553074
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 19952 543218 20188 543454
rect 19952 542898 20188 543134
rect 25882 543218 26118 543454
rect 25882 542898 26118 543134
rect 31813 543218 32049 543454
rect 31813 542898 32049 543134
rect 46952 543218 47188 543454
rect 46952 542898 47188 543134
rect 52882 543218 53118 543454
rect 52882 542898 53118 543134
rect 58813 543218 59049 543454
rect 58813 542898 59049 543134
rect 73952 543218 74188 543454
rect 73952 542898 74188 543134
rect 79882 543218 80118 543454
rect 79882 542898 80118 543134
rect 85813 543218 86049 543454
rect 85813 542898 86049 543134
rect 100952 543218 101188 543454
rect 100952 542898 101188 543134
rect 106882 543218 107118 543454
rect 106882 542898 107118 543134
rect 112813 543218 113049 543454
rect 112813 542898 113049 543134
rect 127952 543218 128188 543454
rect 127952 542898 128188 543134
rect 133882 543218 134118 543454
rect 133882 542898 134118 543134
rect 139813 543218 140049 543454
rect 139813 542898 140049 543134
rect 154952 543218 155188 543454
rect 154952 542898 155188 543134
rect 160882 543218 161118 543454
rect 160882 542898 161118 543134
rect 166813 543218 167049 543454
rect 166813 542898 167049 543134
rect 181952 543218 182188 543454
rect 181952 542898 182188 543134
rect 187882 543218 188118 543454
rect 187882 542898 188118 543134
rect 193813 543218 194049 543454
rect 193813 542898 194049 543134
rect 208952 543218 209188 543454
rect 208952 542898 209188 543134
rect 214882 543218 215118 543454
rect 214882 542898 215118 543134
rect 220813 543218 221049 543454
rect 220813 542898 221049 543134
rect 235952 543218 236188 543454
rect 235952 542898 236188 543134
rect 241882 543218 242118 543454
rect 241882 542898 242118 543134
rect 247813 543218 248049 543454
rect 247813 542898 248049 543134
rect 262952 543218 263188 543454
rect 262952 542898 263188 543134
rect 268882 543218 269118 543454
rect 268882 542898 269118 543134
rect 274813 543218 275049 543454
rect 274813 542898 275049 543134
rect 289952 543218 290188 543454
rect 289952 542898 290188 543134
rect 295882 543218 296118 543454
rect 295882 542898 296118 543134
rect 301813 543218 302049 543454
rect 301813 542898 302049 543134
rect 316952 543218 317188 543454
rect 316952 542898 317188 543134
rect 322882 543218 323118 543454
rect 322882 542898 323118 543134
rect 328813 543218 329049 543454
rect 328813 542898 329049 543134
rect 343952 543218 344188 543454
rect 343952 542898 344188 543134
rect 349882 543218 350118 543454
rect 349882 542898 350118 543134
rect 355813 543218 356049 543454
rect 355813 542898 356049 543134
rect 370952 543218 371188 543454
rect 370952 542898 371188 543134
rect 376882 543218 377118 543454
rect 376882 542898 377118 543134
rect 382813 543218 383049 543454
rect 382813 542898 383049 543134
rect 397952 543218 398188 543454
rect 397952 542898 398188 543134
rect 403882 543218 404118 543454
rect 403882 542898 404118 543134
rect 409813 543218 410049 543454
rect 409813 542898 410049 543134
rect 424952 543218 425188 543454
rect 424952 542898 425188 543134
rect 430882 543218 431118 543454
rect 430882 542898 431118 543134
rect 436813 543218 437049 543454
rect 436813 542898 437049 543134
rect 451952 543218 452188 543454
rect 451952 542898 452188 543134
rect 457882 543218 458118 543454
rect 457882 542898 458118 543134
rect 463813 543218 464049 543454
rect 463813 542898 464049 543134
rect 478952 543218 479188 543454
rect 478952 542898 479188 543134
rect 484882 543218 485118 543454
rect 484882 542898 485118 543134
rect 490813 543218 491049 543454
rect 490813 542898 491049 543134
rect 505952 543218 506188 543454
rect 505952 542898 506188 543134
rect 511882 543218 512118 543454
rect 511882 542898 512118 543134
rect 517813 543218 518049 543454
rect 517813 542898 518049 543134
rect 532952 543218 533188 543454
rect 532952 542898 533188 543134
rect 538882 543218 539118 543454
rect 538882 542898 539118 543134
rect 544813 543218 545049 543454
rect 544813 542898 545049 543134
rect 559826 543218 560062 543454
rect 560146 543218 560382 543454
rect 559826 542898 560062 543134
rect 560146 542898 560382 543134
rect 10826 534218 11062 534454
rect 11146 534218 11382 534454
rect 10826 533898 11062 534134
rect 11146 533898 11382 534134
rect 22916 534218 23152 534454
rect 22916 533898 23152 534134
rect 28847 534218 29083 534454
rect 28847 533898 29083 534134
rect 49916 534218 50152 534454
rect 49916 533898 50152 534134
rect 55847 534218 56083 534454
rect 55847 533898 56083 534134
rect 76916 534218 77152 534454
rect 76916 533898 77152 534134
rect 82847 534218 83083 534454
rect 82847 533898 83083 534134
rect 103916 534218 104152 534454
rect 103916 533898 104152 534134
rect 109847 534218 110083 534454
rect 109847 533898 110083 534134
rect 130916 534218 131152 534454
rect 130916 533898 131152 534134
rect 136847 534218 137083 534454
rect 136847 533898 137083 534134
rect 157916 534218 158152 534454
rect 157916 533898 158152 534134
rect 163847 534218 164083 534454
rect 163847 533898 164083 534134
rect 184916 534218 185152 534454
rect 184916 533898 185152 534134
rect 190847 534218 191083 534454
rect 190847 533898 191083 534134
rect 211916 534218 212152 534454
rect 211916 533898 212152 534134
rect 217847 534218 218083 534454
rect 217847 533898 218083 534134
rect 238916 534218 239152 534454
rect 238916 533898 239152 534134
rect 244847 534218 245083 534454
rect 244847 533898 245083 534134
rect 265916 534218 266152 534454
rect 265916 533898 266152 534134
rect 271847 534218 272083 534454
rect 271847 533898 272083 534134
rect 292916 534218 293152 534454
rect 292916 533898 293152 534134
rect 298847 534218 299083 534454
rect 298847 533898 299083 534134
rect 319916 534218 320152 534454
rect 319916 533898 320152 534134
rect 325847 534218 326083 534454
rect 325847 533898 326083 534134
rect 346916 534218 347152 534454
rect 346916 533898 347152 534134
rect 352847 534218 353083 534454
rect 352847 533898 353083 534134
rect 373916 534218 374152 534454
rect 373916 533898 374152 534134
rect 379847 534218 380083 534454
rect 379847 533898 380083 534134
rect 400916 534218 401152 534454
rect 400916 533898 401152 534134
rect 406847 534218 407083 534454
rect 406847 533898 407083 534134
rect 427916 534218 428152 534454
rect 427916 533898 428152 534134
rect 433847 534218 434083 534454
rect 433847 533898 434083 534134
rect 454916 534218 455152 534454
rect 454916 533898 455152 534134
rect 460847 534218 461083 534454
rect 460847 533898 461083 534134
rect 481916 534218 482152 534454
rect 481916 533898 482152 534134
rect 487847 534218 488083 534454
rect 487847 533898 488083 534134
rect 508916 534218 509152 534454
rect 508916 533898 509152 534134
rect 514847 534218 515083 534454
rect 514847 533898 515083 534134
rect 535916 534218 536152 534454
rect 535916 533898 536152 534134
rect 541847 534218 542083 534454
rect 541847 533898 542083 534134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 28826 526158 29062 526394
rect 29146 526158 29382 526394
rect 28826 525838 29062 526074
rect 29146 525838 29382 526074
rect 37826 525218 38062 525454
rect 38146 525218 38382 525454
rect 37826 524898 38062 525134
rect 38146 524898 38382 525134
rect 46826 526158 47062 526394
rect 47146 526158 47382 526394
rect 46826 525838 47062 526074
rect 47146 525838 47382 526074
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 64826 526158 65062 526394
rect 65146 526158 65382 526394
rect 64826 525838 65062 526074
rect 65146 525838 65382 526074
rect 73826 525218 74062 525454
rect 74146 525218 74382 525454
rect 73826 524898 74062 525134
rect 74146 524898 74382 525134
rect 82826 526158 83062 526394
rect 83146 526158 83382 526394
rect 82826 525838 83062 526074
rect 83146 525838 83382 526074
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 100826 526158 101062 526394
rect 101146 526158 101382 526394
rect 100826 525838 101062 526074
rect 101146 525838 101382 526074
rect 109826 525218 110062 525454
rect 110146 525218 110382 525454
rect 109826 524898 110062 525134
rect 110146 524898 110382 525134
rect 118826 526158 119062 526394
rect 119146 526158 119382 526394
rect 118826 525838 119062 526074
rect 119146 525838 119382 526074
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 136826 526158 137062 526394
rect 137146 526158 137382 526394
rect 136826 525838 137062 526074
rect 137146 525838 137382 526074
rect 145826 525218 146062 525454
rect 146146 525218 146382 525454
rect 145826 524898 146062 525134
rect 146146 524898 146382 525134
rect 154826 526158 155062 526394
rect 155146 526158 155382 526394
rect 154826 525838 155062 526074
rect 155146 525838 155382 526074
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 172826 526158 173062 526394
rect 173146 526158 173382 526394
rect 172826 525838 173062 526074
rect 173146 525838 173382 526074
rect 181826 525218 182062 525454
rect 182146 525218 182382 525454
rect 181826 524898 182062 525134
rect 182146 524898 182382 525134
rect 190826 526158 191062 526394
rect 191146 526158 191382 526394
rect 190826 525838 191062 526074
rect 191146 525838 191382 526074
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 208826 526158 209062 526394
rect 209146 526158 209382 526394
rect 208826 525838 209062 526074
rect 209146 525838 209382 526074
rect 217826 525218 218062 525454
rect 218146 525218 218382 525454
rect 217826 524898 218062 525134
rect 218146 524898 218382 525134
rect 226826 526158 227062 526394
rect 227146 526158 227382 526394
rect 226826 525838 227062 526074
rect 227146 525838 227382 526074
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 244826 526158 245062 526394
rect 245146 526158 245382 526394
rect 244826 525838 245062 526074
rect 245146 525838 245382 526074
rect 253826 525218 254062 525454
rect 254146 525218 254382 525454
rect 253826 524898 254062 525134
rect 254146 524898 254382 525134
rect 262826 526158 263062 526394
rect 263146 526158 263382 526394
rect 262826 525838 263062 526074
rect 263146 525838 263382 526074
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 280826 526158 281062 526394
rect 281146 526158 281382 526394
rect 280826 525838 281062 526074
rect 281146 525838 281382 526074
rect 289826 525218 290062 525454
rect 290146 525218 290382 525454
rect 289826 524898 290062 525134
rect 290146 524898 290382 525134
rect 298826 526158 299062 526394
rect 299146 526158 299382 526394
rect 298826 525838 299062 526074
rect 299146 525838 299382 526074
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 316826 526158 317062 526394
rect 317146 526158 317382 526394
rect 316826 525838 317062 526074
rect 317146 525838 317382 526074
rect 325826 525218 326062 525454
rect 326146 525218 326382 525454
rect 325826 524898 326062 525134
rect 326146 524898 326382 525134
rect 334826 526158 335062 526394
rect 335146 526158 335382 526394
rect 334826 525838 335062 526074
rect 335146 525838 335382 526074
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 352826 526158 353062 526394
rect 353146 526158 353382 526394
rect 352826 525838 353062 526074
rect 353146 525838 353382 526074
rect 361826 525218 362062 525454
rect 362146 525218 362382 525454
rect 361826 524898 362062 525134
rect 362146 524898 362382 525134
rect 370826 526158 371062 526394
rect 371146 526158 371382 526394
rect 370826 525838 371062 526074
rect 371146 525838 371382 526074
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 388826 526158 389062 526394
rect 389146 526158 389382 526394
rect 388826 525838 389062 526074
rect 389146 525838 389382 526074
rect 397826 525218 398062 525454
rect 398146 525218 398382 525454
rect 397826 524898 398062 525134
rect 398146 524898 398382 525134
rect 406826 526158 407062 526394
rect 407146 526158 407382 526394
rect 406826 525838 407062 526074
rect 407146 525838 407382 526074
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 424826 526158 425062 526394
rect 425146 526158 425382 526394
rect 424826 525838 425062 526074
rect 425146 525838 425382 526074
rect 433826 525218 434062 525454
rect 434146 525218 434382 525454
rect 433826 524898 434062 525134
rect 434146 524898 434382 525134
rect 442826 526158 443062 526394
rect 443146 526158 443382 526394
rect 442826 525838 443062 526074
rect 443146 525838 443382 526074
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 460826 526158 461062 526394
rect 461146 526158 461382 526394
rect 460826 525838 461062 526074
rect 461146 525838 461382 526074
rect 469826 525218 470062 525454
rect 470146 525218 470382 525454
rect 469826 524898 470062 525134
rect 470146 524898 470382 525134
rect 478826 526158 479062 526394
rect 479146 526158 479382 526394
rect 478826 525838 479062 526074
rect 479146 525838 479382 526074
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 496826 526158 497062 526394
rect 497146 526158 497382 526394
rect 496826 525838 497062 526074
rect 497146 525838 497382 526074
rect 505826 525218 506062 525454
rect 506146 525218 506382 525454
rect 505826 524898 506062 525134
rect 506146 524898 506382 525134
rect 514826 526158 515062 526394
rect 515146 526158 515382 526394
rect 514826 525838 515062 526074
rect 515146 525838 515382 526074
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 532826 526158 533062 526394
rect 533146 526158 533382 526394
rect 532826 525838 533062 526074
rect 533146 525838 533382 526074
rect 541826 525218 542062 525454
rect 542146 525218 542382 525454
rect 541826 524898 542062 525134
rect 542146 524898 542382 525134
rect 550826 526158 551062 526394
rect 551146 526158 551382 526394
rect 550826 525838 551062 526074
rect 551146 525838 551382 526074
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 22916 516218 23152 516454
rect 22916 515898 23152 516134
rect 28847 516218 29083 516454
rect 28847 515898 29083 516134
rect 49916 516218 50152 516454
rect 49916 515898 50152 516134
rect 55847 516218 56083 516454
rect 55847 515898 56083 516134
rect 76916 516218 77152 516454
rect 76916 515898 77152 516134
rect 82847 516218 83083 516454
rect 82847 515898 83083 516134
rect 103916 516218 104152 516454
rect 103916 515898 104152 516134
rect 109847 516218 110083 516454
rect 109847 515898 110083 516134
rect 130916 516218 131152 516454
rect 130916 515898 131152 516134
rect 136847 516218 137083 516454
rect 136847 515898 137083 516134
rect 157916 516218 158152 516454
rect 157916 515898 158152 516134
rect 163847 516218 164083 516454
rect 163847 515898 164083 516134
rect 184916 516218 185152 516454
rect 184916 515898 185152 516134
rect 190847 516218 191083 516454
rect 190847 515898 191083 516134
rect 211916 516218 212152 516454
rect 211916 515898 212152 516134
rect 217847 516218 218083 516454
rect 217847 515898 218083 516134
rect 238916 516218 239152 516454
rect 238916 515898 239152 516134
rect 244847 516218 245083 516454
rect 244847 515898 245083 516134
rect 265916 516218 266152 516454
rect 265916 515898 266152 516134
rect 271847 516218 272083 516454
rect 271847 515898 272083 516134
rect 292916 516218 293152 516454
rect 292916 515898 293152 516134
rect 298847 516218 299083 516454
rect 298847 515898 299083 516134
rect 319916 516218 320152 516454
rect 319916 515898 320152 516134
rect 325847 516218 326083 516454
rect 325847 515898 326083 516134
rect 346916 516218 347152 516454
rect 346916 515898 347152 516134
rect 352847 516218 353083 516454
rect 352847 515898 353083 516134
rect 373916 516218 374152 516454
rect 373916 515898 374152 516134
rect 379847 516218 380083 516454
rect 379847 515898 380083 516134
rect 400916 516218 401152 516454
rect 400916 515898 401152 516134
rect 406847 516218 407083 516454
rect 406847 515898 407083 516134
rect 427916 516218 428152 516454
rect 427916 515898 428152 516134
rect 433847 516218 434083 516454
rect 433847 515898 434083 516134
rect 454916 516218 455152 516454
rect 454916 515898 455152 516134
rect 460847 516218 461083 516454
rect 460847 515898 461083 516134
rect 481916 516218 482152 516454
rect 481916 515898 482152 516134
rect 487847 516218 488083 516454
rect 487847 515898 488083 516134
rect 508916 516218 509152 516454
rect 508916 515898 509152 516134
rect 514847 516218 515083 516454
rect 514847 515898 515083 516134
rect 535916 516218 536152 516454
rect 535916 515898 536152 516134
rect 541847 516218 542083 516454
rect 541847 515898 542083 516134
rect 19952 507218 20188 507454
rect 19952 506898 20188 507134
rect 25882 507218 26118 507454
rect 25882 506898 26118 507134
rect 31813 507218 32049 507454
rect 31813 506898 32049 507134
rect 46952 507218 47188 507454
rect 46952 506898 47188 507134
rect 52882 507218 53118 507454
rect 52882 506898 53118 507134
rect 58813 507218 59049 507454
rect 58813 506898 59049 507134
rect 73952 507218 74188 507454
rect 73952 506898 74188 507134
rect 79882 507218 80118 507454
rect 79882 506898 80118 507134
rect 85813 507218 86049 507454
rect 85813 506898 86049 507134
rect 100952 507218 101188 507454
rect 100952 506898 101188 507134
rect 106882 507218 107118 507454
rect 106882 506898 107118 507134
rect 112813 507218 113049 507454
rect 112813 506898 113049 507134
rect 127952 507218 128188 507454
rect 127952 506898 128188 507134
rect 133882 507218 134118 507454
rect 133882 506898 134118 507134
rect 139813 507218 140049 507454
rect 139813 506898 140049 507134
rect 154952 507218 155188 507454
rect 154952 506898 155188 507134
rect 160882 507218 161118 507454
rect 160882 506898 161118 507134
rect 166813 507218 167049 507454
rect 166813 506898 167049 507134
rect 181952 507218 182188 507454
rect 181952 506898 182188 507134
rect 187882 507218 188118 507454
rect 187882 506898 188118 507134
rect 193813 507218 194049 507454
rect 193813 506898 194049 507134
rect 208952 507218 209188 507454
rect 208952 506898 209188 507134
rect 214882 507218 215118 507454
rect 214882 506898 215118 507134
rect 220813 507218 221049 507454
rect 220813 506898 221049 507134
rect 235952 507218 236188 507454
rect 235952 506898 236188 507134
rect 241882 507218 242118 507454
rect 241882 506898 242118 507134
rect 247813 507218 248049 507454
rect 247813 506898 248049 507134
rect 262952 507218 263188 507454
rect 262952 506898 263188 507134
rect 268882 507218 269118 507454
rect 268882 506898 269118 507134
rect 274813 507218 275049 507454
rect 274813 506898 275049 507134
rect 289952 507218 290188 507454
rect 289952 506898 290188 507134
rect 295882 507218 296118 507454
rect 295882 506898 296118 507134
rect 301813 507218 302049 507454
rect 301813 506898 302049 507134
rect 316952 507218 317188 507454
rect 316952 506898 317188 507134
rect 322882 507218 323118 507454
rect 322882 506898 323118 507134
rect 328813 507218 329049 507454
rect 328813 506898 329049 507134
rect 343952 507218 344188 507454
rect 343952 506898 344188 507134
rect 349882 507218 350118 507454
rect 349882 506898 350118 507134
rect 355813 507218 356049 507454
rect 355813 506898 356049 507134
rect 370952 507218 371188 507454
rect 370952 506898 371188 507134
rect 376882 507218 377118 507454
rect 376882 506898 377118 507134
rect 382813 507218 383049 507454
rect 382813 506898 383049 507134
rect 397952 507218 398188 507454
rect 397952 506898 398188 507134
rect 403882 507218 404118 507454
rect 403882 506898 404118 507134
rect 409813 507218 410049 507454
rect 409813 506898 410049 507134
rect 424952 507218 425188 507454
rect 424952 506898 425188 507134
rect 430882 507218 431118 507454
rect 430882 506898 431118 507134
rect 436813 507218 437049 507454
rect 436813 506898 437049 507134
rect 451952 507218 452188 507454
rect 451952 506898 452188 507134
rect 457882 507218 458118 507454
rect 457882 506898 458118 507134
rect 463813 507218 464049 507454
rect 463813 506898 464049 507134
rect 478952 507218 479188 507454
rect 478952 506898 479188 507134
rect 484882 507218 485118 507454
rect 484882 506898 485118 507134
rect 490813 507218 491049 507454
rect 490813 506898 491049 507134
rect 505952 507218 506188 507454
rect 505952 506898 506188 507134
rect 511882 507218 512118 507454
rect 511882 506898 512118 507134
rect 517813 507218 518049 507454
rect 517813 506898 518049 507134
rect 532952 507218 533188 507454
rect 532952 506898 533188 507134
rect 538882 507218 539118 507454
rect 538882 506898 539118 507134
rect 544813 507218 545049 507454
rect 544813 506898 545049 507134
rect 559826 507218 560062 507454
rect 560146 507218 560382 507454
rect 559826 506898 560062 507134
rect 560146 506898 560382 507134
rect 10826 498218 11062 498454
rect 11146 498218 11382 498454
rect 10826 497898 11062 498134
rect 11146 497898 11382 498134
rect 19826 499158 20062 499394
rect 20146 499158 20382 499394
rect 19826 498838 20062 499074
rect 20146 498838 20382 499074
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 37826 499158 38062 499394
rect 38146 499158 38382 499394
rect 37826 498838 38062 499074
rect 38146 498838 38382 499074
rect 46826 498218 47062 498454
rect 47146 498218 47382 498454
rect 46826 497898 47062 498134
rect 47146 497898 47382 498134
rect 55826 499158 56062 499394
rect 56146 499158 56382 499394
rect 55826 498838 56062 499074
rect 56146 498838 56382 499074
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 73826 499158 74062 499394
rect 74146 499158 74382 499394
rect 73826 498838 74062 499074
rect 74146 498838 74382 499074
rect 82826 498218 83062 498454
rect 83146 498218 83382 498454
rect 82826 497898 83062 498134
rect 83146 497898 83382 498134
rect 91826 499158 92062 499394
rect 92146 499158 92382 499394
rect 91826 498838 92062 499074
rect 92146 498838 92382 499074
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 109826 499158 110062 499394
rect 110146 499158 110382 499394
rect 109826 498838 110062 499074
rect 110146 498838 110382 499074
rect 118826 498218 119062 498454
rect 119146 498218 119382 498454
rect 118826 497898 119062 498134
rect 119146 497898 119382 498134
rect 127826 499158 128062 499394
rect 128146 499158 128382 499394
rect 127826 498838 128062 499074
rect 128146 498838 128382 499074
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 145826 499158 146062 499394
rect 146146 499158 146382 499394
rect 145826 498838 146062 499074
rect 146146 498838 146382 499074
rect 154826 498218 155062 498454
rect 155146 498218 155382 498454
rect 154826 497898 155062 498134
rect 155146 497898 155382 498134
rect 163826 499158 164062 499394
rect 164146 499158 164382 499394
rect 163826 498838 164062 499074
rect 164146 498838 164382 499074
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 181826 499158 182062 499394
rect 182146 499158 182382 499394
rect 181826 498838 182062 499074
rect 182146 498838 182382 499074
rect 190826 498218 191062 498454
rect 191146 498218 191382 498454
rect 190826 497898 191062 498134
rect 191146 497898 191382 498134
rect 199826 499158 200062 499394
rect 200146 499158 200382 499394
rect 199826 498838 200062 499074
rect 200146 498838 200382 499074
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 217826 499158 218062 499394
rect 218146 499158 218382 499394
rect 217826 498838 218062 499074
rect 218146 498838 218382 499074
rect 226826 498218 227062 498454
rect 227146 498218 227382 498454
rect 226826 497898 227062 498134
rect 227146 497898 227382 498134
rect 235826 499158 236062 499394
rect 236146 499158 236382 499394
rect 235826 498838 236062 499074
rect 236146 498838 236382 499074
rect 244826 498218 245062 498454
rect 245146 498218 245382 498454
rect 244826 497898 245062 498134
rect 245146 497898 245382 498134
rect 253826 499158 254062 499394
rect 254146 499158 254382 499394
rect 253826 498838 254062 499074
rect 254146 498838 254382 499074
rect 262826 498218 263062 498454
rect 263146 498218 263382 498454
rect 262826 497898 263062 498134
rect 263146 497898 263382 498134
rect 271826 499158 272062 499394
rect 272146 499158 272382 499394
rect 271826 498838 272062 499074
rect 272146 498838 272382 499074
rect 280826 498218 281062 498454
rect 281146 498218 281382 498454
rect 280826 497898 281062 498134
rect 281146 497898 281382 498134
rect 289826 499158 290062 499394
rect 290146 499158 290382 499394
rect 289826 498838 290062 499074
rect 290146 498838 290382 499074
rect 298826 498218 299062 498454
rect 299146 498218 299382 498454
rect 298826 497898 299062 498134
rect 299146 497898 299382 498134
rect 307826 499158 308062 499394
rect 308146 499158 308382 499394
rect 307826 498838 308062 499074
rect 308146 498838 308382 499074
rect 316826 498218 317062 498454
rect 317146 498218 317382 498454
rect 316826 497898 317062 498134
rect 317146 497898 317382 498134
rect 325826 499158 326062 499394
rect 326146 499158 326382 499394
rect 325826 498838 326062 499074
rect 326146 498838 326382 499074
rect 334826 498218 335062 498454
rect 335146 498218 335382 498454
rect 334826 497898 335062 498134
rect 335146 497898 335382 498134
rect 343826 499158 344062 499394
rect 344146 499158 344382 499394
rect 343826 498838 344062 499074
rect 344146 498838 344382 499074
rect 352826 498218 353062 498454
rect 353146 498218 353382 498454
rect 352826 497898 353062 498134
rect 353146 497898 353382 498134
rect 361826 499158 362062 499394
rect 362146 499158 362382 499394
rect 361826 498838 362062 499074
rect 362146 498838 362382 499074
rect 370826 498218 371062 498454
rect 371146 498218 371382 498454
rect 370826 497898 371062 498134
rect 371146 497898 371382 498134
rect 379826 499158 380062 499394
rect 380146 499158 380382 499394
rect 379826 498838 380062 499074
rect 380146 498838 380382 499074
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 397826 499158 398062 499394
rect 398146 499158 398382 499394
rect 397826 498838 398062 499074
rect 398146 498838 398382 499074
rect 406826 498218 407062 498454
rect 407146 498218 407382 498454
rect 406826 497898 407062 498134
rect 407146 497898 407382 498134
rect 415826 499158 416062 499394
rect 416146 499158 416382 499394
rect 415826 498838 416062 499074
rect 416146 498838 416382 499074
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 433826 499158 434062 499394
rect 434146 499158 434382 499394
rect 433826 498838 434062 499074
rect 434146 498838 434382 499074
rect 442826 498218 443062 498454
rect 443146 498218 443382 498454
rect 442826 497898 443062 498134
rect 443146 497898 443382 498134
rect 451826 499158 452062 499394
rect 452146 499158 452382 499394
rect 451826 498838 452062 499074
rect 452146 498838 452382 499074
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 469826 499158 470062 499394
rect 470146 499158 470382 499394
rect 469826 498838 470062 499074
rect 470146 498838 470382 499074
rect 478826 498218 479062 498454
rect 479146 498218 479382 498454
rect 478826 497898 479062 498134
rect 479146 497898 479382 498134
rect 487826 499158 488062 499394
rect 488146 499158 488382 499394
rect 487826 498838 488062 499074
rect 488146 498838 488382 499074
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 505826 499158 506062 499394
rect 506146 499158 506382 499394
rect 505826 498838 506062 499074
rect 506146 498838 506382 499074
rect 514826 498218 515062 498454
rect 515146 498218 515382 498454
rect 514826 497898 515062 498134
rect 515146 497898 515382 498134
rect 523826 499158 524062 499394
rect 524146 499158 524382 499394
rect 523826 498838 524062 499074
rect 524146 498838 524382 499074
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 541826 499158 542062 499394
rect 542146 499158 542382 499394
rect 541826 498838 542062 499074
rect 542146 498838 542382 499074
rect 550826 498218 551062 498454
rect 551146 498218 551382 498454
rect 550826 497898 551062 498134
rect 551146 497898 551382 498134
rect 19952 489218 20188 489454
rect 19952 488898 20188 489134
rect 25882 489218 26118 489454
rect 25882 488898 26118 489134
rect 31813 489218 32049 489454
rect 31813 488898 32049 489134
rect 46952 489218 47188 489454
rect 46952 488898 47188 489134
rect 52882 489218 53118 489454
rect 52882 488898 53118 489134
rect 58813 489218 59049 489454
rect 58813 488898 59049 489134
rect 73952 489218 74188 489454
rect 73952 488898 74188 489134
rect 79882 489218 80118 489454
rect 79882 488898 80118 489134
rect 85813 489218 86049 489454
rect 85813 488898 86049 489134
rect 100952 489218 101188 489454
rect 100952 488898 101188 489134
rect 106882 489218 107118 489454
rect 106882 488898 107118 489134
rect 112813 489218 113049 489454
rect 112813 488898 113049 489134
rect 127952 489218 128188 489454
rect 127952 488898 128188 489134
rect 133882 489218 134118 489454
rect 133882 488898 134118 489134
rect 139813 489218 140049 489454
rect 139813 488898 140049 489134
rect 154952 489218 155188 489454
rect 154952 488898 155188 489134
rect 160882 489218 161118 489454
rect 160882 488898 161118 489134
rect 166813 489218 167049 489454
rect 166813 488898 167049 489134
rect 181952 489218 182188 489454
rect 181952 488898 182188 489134
rect 187882 489218 188118 489454
rect 187882 488898 188118 489134
rect 193813 489218 194049 489454
rect 193813 488898 194049 489134
rect 208952 489218 209188 489454
rect 208952 488898 209188 489134
rect 214882 489218 215118 489454
rect 214882 488898 215118 489134
rect 220813 489218 221049 489454
rect 220813 488898 221049 489134
rect 235952 489218 236188 489454
rect 235952 488898 236188 489134
rect 241882 489218 242118 489454
rect 241882 488898 242118 489134
rect 247813 489218 248049 489454
rect 247813 488898 248049 489134
rect 262952 489218 263188 489454
rect 262952 488898 263188 489134
rect 268882 489218 269118 489454
rect 268882 488898 269118 489134
rect 274813 489218 275049 489454
rect 274813 488898 275049 489134
rect 289952 489218 290188 489454
rect 289952 488898 290188 489134
rect 295882 489218 296118 489454
rect 295882 488898 296118 489134
rect 301813 489218 302049 489454
rect 301813 488898 302049 489134
rect 316952 489218 317188 489454
rect 316952 488898 317188 489134
rect 322882 489218 323118 489454
rect 322882 488898 323118 489134
rect 328813 489218 329049 489454
rect 328813 488898 329049 489134
rect 343952 489218 344188 489454
rect 343952 488898 344188 489134
rect 349882 489218 350118 489454
rect 349882 488898 350118 489134
rect 355813 489218 356049 489454
rect 355813 488898 356049 489134
rect 370952 489218 371188 489454
rect 370952 488898 371188 489134
rect 376882 489218 377118 489454
rect 376882 488898 377118 489134
rect 382813 489218 383049 489454
rect 382813 488898 383049 489134
rect 397952 489218 398188 489454
rect 397952 488898 398188 489134
rect 403882 489218 404118 489454
rect 403882 488898 404118 489134
rect 409813 489218 410049 489454
rect 409813 488898 410049 489134
rect 424952 489218 425188 489454
rect 424952 488898 425188 489134
rect 430882 489218 431118 489454
rect 430882 488898 431118 489134
rect 436813 489218 437049 489454
rect 436813 488898 437049 489134
rect 451952 489218 452188 489454
rect 451952 488898 452188 489134
rect 457882 489218 458118 489454
rect 457882 488898 458118 489134
rect 463813 489218 464049 489454
rect 463813 488898 464049 489134
rect 478952 489218 479188 489454
rect 478952 488898 479188 489134
rect 484882 489218 485118 489454
rect 484882 488898 485118 489134
rect 490813 489218 491049 489454
rect 490813 488898 491049 489134
rect 505952 489218 506188 489454
rect 505952 488898 506188 489134
rect 511882 489218 512118 489454
rect 511882 488898 512118 489134
rect 517813 489218 518049 489454
rect 517813 488898 518049 489134
rect 532952 489218 533188 489454
rect 532952 488898 533188 489134
rect 538882 489218 539118 489454
rect 538882 488898 539118 489134
rect 544813 489218 545049 489454
rect 544813 488898 545049 489134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 22916 480218 23152 480454
rect 22916 479898 23152 480134
rect 28847 480218 29083 480454
rect 28847 479898 29083 480134
rect 49916 480218 50152 480454
rect 49916 479898 50152 480134
rect 55847 480218 56083 480454
rect 55847 479898 56083 480134
rect 76916 480218 77152 480454
rect 76916 479898 77152 480134
rect 82847 480218 83083 480454
rect 82847 479898 83083 480134
rect 103916 480218 104152 480454
rect 103916 479898 104152 480134
rect 109847 480218 110083 480454
rect 109847 479898 110083 480134
rect 130916 480218 131152 480454
rect 130916 479898 131152 480134
rect 136847 480218 137083 480454
rect 136847 479898 137083 480134
rect 157916 480218 158152 480454
rect 157916 479898 158152 480134
rect 163847 480218 164083 480454
rect 163847 479898 164083 480134
rect 184916 480218 185152 480454
rect 184916 479898 185152 480134
rect 190847 480218 191083 480454
rect 190847 479898 191083 480134
rect 211916 480218 212152 480454
rect 211916 479898 212152 480134
rect 217847 480218 218083 480454
rect 217847 479898 218083 480134
rect 238916 480218 239152 480454
rect 238916 479898 239152 480134
rect 244847 480218 245083 480454
rect 244847 479898 245083 480134
rect 265916 480218 266152 480454
rect 265916 479898 266152 480134
rect 271847 480218 272083 480454
rect 271847 479898 272083 480134
rect 292916 480218 293152 480454
rect 292916 479898 293152 480134
rect 298847 480218 299083 480454
rect 298847 479898 299083 480134
rect 319916 480218 320152 480454
rect 319916 479898 320152 480134
rect 325847 480218 326083 480454
rect 325847 479898 326083 480134
rect 346916 480218 347152 480454
rect 346916 479898 347152 480134
rect 352847 480218 353083 480454
rect 352847 479898 353083 480134
rect 373916 480218 374152 480454
rect 373916 479898 374152 480134
rect 379847 480218 380083 480454
rect 379847 479898 380083 480134
rect 400916 480218 401152 480454
rect 400916 479898 401152 480134
rect 406847 480218 407083 480454
rect 406847 479898 407083 480134
rect 427916 480218 428152 480454
rect 427916 479898 428152 480134
rect 433847 480218 434083 480454
rect 433847 479898 434083 480134
rect 454916 480218 455152 480454
rect 454916 479898 455152 480134
rect 460847 480218 461083 480454
rect 460847 479898 461083 480134
rect 481916 480218 482152 480454
rect 481916 479898 482152 480134
rect 487847 480218 488083 480454
rect 487847 479898 488083 480134
rect 508916 480218 509152 480454
rect 508916 479898 509152 480134
rect 514847 480218 515083 480454
rect 514847 479898 515083 480134
rect 535916 480218 536152 480454
rect 535916 479898 536152 480134
rect 541847 480218 542083 480454
rect 541847 479898 542083 480134
rect 19826 471218 20062 471454
rect 20146 471218 20382 471454
rect 19826 470898 20062 471134
rect 20146 470898 20382 471134
rect 28826 472158 29062 472394
rect 29146 472158 29382 472394
rect 28826 471838 29062 472074
rect 29146 471838 29382 472074
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 46826 472158 47062 472394
rect 47146 472158 47382 472394
rect 46826 471838 47062 472074
rect 47146 471838 47382 472074
rect 55826 471218 56062 471454
rect 56146 471218 56382 471454
rect 55826 470898 56062 471134
rect 56146 470898 56382 471134
rect 64826 472158 65062 472394
rect 65146 472158 65382 472394
rect 64826 471838 65062 472074
rect 65146 471838 65382 472074
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 82826 472158 83062 472394
rect 83146 472158 83382 472394
rect 82826 471838 83062 472074
rect 83146 471838 83382 472074
rect 91826 471218 92062 471454
rect 92146 471218 92382 471454
rect 91826 470898 92062 471134
rect 92146 470898 92382 471134
rect 100826 472158 101062 472394
rect 101146 472158 101382 472394
rect 100826 471838 101062 472074
rect 101146 471838 101382 472074
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 118826 472158 119062 472394
rect 119146 472158 119382 472394
rect 118826 471838 119062 472074
rect 119146 471838 119382 472074
rect 127826 471218 128062 471454
rect 128146 471218 128382 471454
rect 127826 470898 128062 471134
rect 128146 470898 128382 471134
rect 136826 472158 137062 472394
rect 137146 472158 137382 472394
rect 136826 471838 137062 472074
rect 137146 471838 137382 472074
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 154826 472158 155062 472394
rect 155146 472158 155382 472394
rect 154826 471838 155062 472074
rect 155146 471838 155382 472074
rect 163826 471218 164062 471454
rect 164146 471218 164382 471454
rect 163826 470898 164062 471134
rect 164146 470898 164382 471134
rect 172826 472158 173062 472394
rect 173146 472158 173382 472394
rect 172826 471838 173062 472074
rect 173146 471838 173382 472074
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 190826 472158 191062 472394
rect 191146 472158 191382 472394
rect 190826 471838 191062 472074
rect 191146 471838 191382 472074
rect 199826 471218 200062 471454
rect 200146 471218 200382 471454
rect 199826 470898 200062 471134
rect 200146 470898 200382 471134
rect 208826 472158 209062 472394
rect 209146 472158 209382 472394
rect 208826 471838 209062 472074
rect 209146 471838 209382 472074
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 226826 472158 227062 472394
rect 227146 472158 227382 472394
rect 226826 471838 227062 472074
rect 227146 471838 227382 472074
rect 235826 471218 236062 471454
rect 236146 471218 236382 471454
rect 235826 470898 236062 471134
rect 236146 470898 236382 471134
rect 244826 472158 245062 472394
rect 245146 472158 245382 472394
rect 244826 471838 245062 472074
rect 245146 471838 245382 472074
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 262826 472158 263062 472394
rect 263146 472158 263382 472394
rect 262826 471838 263062 472074
rect 263146 471838 263382 472074
rect 271826 471218 272062 471454
rect 272146 471218 272382 471454
rect 271826 470898 272062 471134
rect 272146 470898 272382 471134
rect 280826 472158 281062 472394
rect 281146 472158 281382 472394
rect 280826 471838 281062 472074
rect 281146 471838 281382 472074
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 298826 472158 299062 472394
rect 299146 472158 299382 472394
rect 298826 471838 299062 472074
rect 299146 471838 299382 472074
rect 307826 471218 308062 471454
rect 308146 471218 308382 471454
rect 307826 470898 308062 471134
rect 308146 470898 308382 471134
rect 316826 472158 317062 472394
rect 317146 472158 317382 472394
rect 316826 471838 317062 472074
rect 317146 471838 317382 472074
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 334826 472158 335062 472394
rect 335146 472158 335382 472394
rect 334826 471838 335062 472074
rect 335146 471838 335382 472074
rect 343826 471218 344062 471454
rect 344146 471218 344382 471454
rect 343826 470898 344062 471134
rect 344146 470898 344382 471134
rect 352826 472158 353062 472394
rect 353146 472158 353382 472394
rect 352826 471838 353062 472074
rect 353146 471838 353382 472074
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 370826 472158 371062 472394
rect 371146 472158 371382 472394
rect 370826 471838 371062 472074
rect 371146 471838 371382 472074
rect 379826 471218 380062 471454
rect 380146 471218 380382 471454
rect 379826 470898 380062 471134
rect 380146 470898 380382 471134
rect 388826 472158 389062 472394
rect 389146 472158 389382 472394
rect 388826 471838 389062 472074
rect 389146 471838 389382 472074
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 406826 472158 407062 472394
rect 407146 472158 407382 472394
rect 406826 471838 407062 472074
rect 407146 471838 407382 472074
rect 415826 471218 416062 471454
rect 416146 471218 416382 471454
rect 415826 470898 416062 471134
rect 416146 470898 416382 471134
rect 424826 472158 425062 472394
rect 425146 472158 425382 472394
rect 424826 471838 425062 472074
rect 425146 471838 425382 472074
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 442826 472158 443062 472394
rect 443146 472158 443382 472394
rect 442826 471838 443062 472074
rect 443146 471838 443382 472074
rect 451826 471218 452062 471454
rect 452146 471218 452382 471454
rect 451826 470898 452062 471134
rect 452146 470898 452382 471134
rect 460826 472158 461062 472394
rect 461146 472158 461382 472394
rect 460826 471838 461062 472074
rect 461146 471838 461382 472074
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 478826 472158 479062 472394
rect 479146 472158 479382 472394
rect 478826 471838 479062 472074
rect 479146 471838 479382 472074
rect 487826 471218 488062 471454
rect 488146 471218 488382 471454
rect 487826 470898 488062 471134
rect 488146 470898 488382 471134
rect 496826 472158 497062 472394
rect 497146 472158 497382 472394
rect 496826 471838 497062 472074
rect 497146 471838 497382 472074
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 514826 472158 515062 472394
rect 515146 472158 515382 472394
rect 514826 471838 515062 472074
rect 515146 471838 515382 472074
rect 523826 471218 524062 471454
rect 524146 471218 524382 471454
rect 523826 470898 524062 471134
rect 524146 470898 524382 471134
rect 532826 472158 533062 472394
rect 533146 472158 533382 472394
rect 532826 471838 533062 472074
rect 533146 471838 533382 472074
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 550826 472158 551062 472394
rect 551146 472158 551382 472394
rect 550826 471838 551062 472074
rect 551146 471838 551382 472074
rect 559826 471218 560062 471454
rect 560146 471218 560382 471454
rect 559826 470898 560062 471134
rect 560146 470898 560382 471134
rect 10826 462218 11062 462454
rect 11146 462218 11382 462454
rect 10826 461898 11062 462134
rect 11146 461898 11382 462134
rect 22916 462218 23152 462454
rect 22916 461898 23152 462134
rect 28847 462218 29083 462454
rect 28847 461898 29083 462134
rect 49916 462218 50152 462454
rect 49916 461898 50152 462134
rect 55847 462218 56083 462454
rect 55847 461898 56083 462134
rect 76916 462218 77152 462454
rect 76916 461898 77152 462134
rect 82847 462218 83083 462454
rect 82847 461898 83083 462134
rect 103916 462218 104152 462454
rect 103916 461898 104152 462134
rect 109847 462218 110083 462454
rect 109847 461898 110083 462134
rect 130916 462218 131152 462454
rect 130916 461898 131152 462134
rect 136847 462218 137083 462454
rect 136847 461898 137083 462134
rect 157916 462218 158152 462454
rect 157916 461898 158152 462134
rect 163847 462218 164083 462454
rect 163847 461898 164083 462134
rect 184916 462218 185152 462454
rect 184916 461898 185152 462134
rect 190847 462218 191083 462454
rect 190847 461898 191083 462134
rect 211916 462218 212152 462454
rect 211916 461898 212152 462134
rect 217847 462218 218083 462454
rect 217847 461898 218083 462134
rect 238916 462218 239152 462454
rect 238916 461898 239152 462134
rect 244847 462218 245083 462454
rect 244847 461898 245083 462134
rect 265916 462218 266152 462454
rect 265916 461898 266152 462134
rect 271847 462218 272083 462454
rect 271847 461898 272083 462134
rect 292916 462218 293152 462454
rect 292916 461898 293152 462134
rect 298847 462218 299083 462454
rect 298847 461898 299083 462134
rect 319916 462218 320152 462454
rect 319916 461898 320152 462134
rect 325847 462218 326083 462454
rect 325847 461898 326083 462134
rect 346916 462218 347152 462454
rect 346916 461898 347152 462134
rect 352847 462218 353083 462454
rect 352847 461898 353083 462134
rect 373916 462218 374152 462454
rect 373916 461898 374152 462134
rect 379847 462218 380083 462454
rect 379847 461898 380083 462134
rect 400916 462218 401152 462454
rect 400916 461898 401152 462134
rect 406847 462218 407083 462454
rect 406847 461898 407083 462134
rect 427916 462218 428152 462454
rect 427916 461898 428152 462134
rect 433847 462218 434083 462454
rect 433847 461898 434083 462134
rect 454916 462218 455152 462454
rect 454916 461898 455152 462134
rect 460847 462218 461083 462454
rect 460847 461898 461083 462134
rect 481916 462218 482152 462454
rect 481916 461898 482152 462134
rect 487847 462218 488083 462454
rect 487847 461898 488083 462134
rect 508916 462218 509152 462454
rect 508916 461898 509152 462134
rect 514847 462218 515083 462454
rect 514847 461898 515083 462134
rect 535916 462218 536152 462454
rect 535916 461898 536152 462134
rect 541847 462218 542083 462454
rect 541847 461898 542083 462134
rect 19952 453218 20188 453454
rect 19952 452898 20188 453134
rect 25882 453218 26118 453454
rect 25882 452898 26118 453134
rect 31813 453218 32049 453454
rect 31813 452898 32049 453134
rect 46952 453218 47188 453454
rect 46952 452898 47188 453134
rect 52882 453218 53118 453454
rect 52882 452898 53118 453134
rect 58813 453218 59049 453454
rect 58813 452898 59049 453134
rect 73952 453218 74188 453454
rect 73952 452898 74188 453134
rect 79882 453218 80118 453454
rect 79882 452898 80118 453134
rect 85813 453218 86049 453454
rect 85813 452898 86049 453134
rect 100952 453218 101188 453454
rect 100952 452898 101188 453134
rect 106882 453218 107118 453454
rect 106882 452898 107118 453134
rect 112813 453218 113049 453454
rect 112813 452898 113049 453134
rect 127952 453218 128188 453454
rect 127952 452898 128188 453134
rect 133882 453218 134118 453454
rect 133882 452898 134118 453134
rect 139813 453218 140049 453454
rect 139813 452898 140049 453134
rect 154952 453218 155188 453454
rect 154952 452898 155188 453134
rect 160882 453218 161118 453454
rect 160882 452898 161118 453134
rect 166813 453218 167049 453454
rect 166813 452898 167049 453134
rect 181952 453218 182188 453454
rect 181952 452898 182188 453134
rect 187882 453218 188118 453454
rect 187882 452898 188118 453134
rect 193813 453218 194049 453454
rect 193813 452898 194049 453134
rect 208952 453218 209188 453454
rect 208952 452898 209188 453134
rect 214882 453218 215118 453454
rect 214882 452898 215118 453134
rect 220813 453218 221049 453454
rect 220813 452898 221049 453134
rect 235952 453218 236188 453454
rect 235952 452898 236188 453134
rect 241882 453218 242118 453454
rect 241882 452898 242118 453134
rect 247813 453218 248049 453454
rect 247813 452898 248049 453134
rect 262952 453218 263188 453454
rect 262952 452898 263188 453134
rect 268882 453218 269118 453454
rect 268882 452898 269118 453134
rect 274813 453218 275049 453454
rect 274813 452898 275049 453134
rect 289952 453218 290188 453454
rect 289952 452898 290188 453134
rect 295882 453218 296118 453454
rect 295882 452898 296118 453134
rect 301813 453218 302049 453454
rect 301813 452898 302049 453134
rect 316952 453218 317188 453454
rect 316952 452898 317188 453134
rect 322882 453218 323118 453454
rect 322882 452898 323118 453134
rect 328813 453218 329049 453454
rect 328813 452898 329049 453134
rect 343952 453218 344188 453454
rect 343952 452898 344188 453134
rect 349882 453218 350118 453454
rect 349882 452898 350118 453134
rect 355813 453218 356049 453454
rect 355813 452898 356049 453134
rect 370952 453218 371188 453454
rect 370952 452898 371188 453134
rect 376882 453218 377118 453454
rect 376882 452898 377118 453134
rect 382813 453218 383049 453454
rect 382813 452898 383049 453134
rect 397952 453218 398188 453454
rect 397952 452898 398188 453134
rect 403882 453218 404118 453454
rect 403882 452898 404118 453134
rect 409813 453218 410049 453454
rect 409813 452898 410049 453134
rect 424952 453218 425188 453454
rect 424952 452898 425188 453134
rect 430882 453218 431118 453454
rect 430882 452898 431118 453134
rect 436813 453218 437049 453454
rect 436813 452898 437049 453134
rect 451952 453218 452188 453454
rect 451952 452898 452188 453134
rect 457882 453218 458118 453454
rect 457882 452898 458118 453134
rect 463813 453218 464049 453454
rect 463813 452898 464049 453134
rect 478952 453218 479188 453454
rect 478952 452898 479188 453134
rect 484882 453218 485118 453454
rect 484882 452898 485118 453134
rect 490813 453218 491049 453454
rect 490813 452898 491049 453134
rect 505952 453218 506188 453454
rect 505952 452898 506188 453134
rect 511882 453218 512118 453454
rect 511882 452898 512118 453134
rect 517813 453218 518049 453454
rect 517813 452898 518049 453134
rect 532952 453218 533188 453454
rect 532952 452898 533188 453134
rect 538882 453218 539118 453454
rect 538882 452898 539118 453134
rect 544813 453218 545049 453454
rect 544813 452898 545049 453134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 19826 445158 20062 445394
rect 20146 445158 20382 445394
rect 19826 444838 20062 445074
rect 20146 444838 20382 445074
rect 28826 444218 29062 444454
rect 29146 444218 29382 444454
rect 28826 443898 29062 444134
rect 29146 443898 29382 444134
rect 37826 445158 38062 445394
rect 38146 445158 38382 445394
rect 37826 444838 38062 445074
rect 38146 444838 38382 445074
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 55826 445158 56062 445394
rect 56146 445158 56382 445394
rect 55826 444838 56062 445074
rect 56146 444838 56382 445074
rect 64826 444218 65062 444454
rect 65146 444218 65382 444454
rect 64826 443898 65062 444134
rect 65146 443898 65382 444134
rect 73826 445158 74062 445394
rect 74146 445158 74382 445394
rect 73826 444838 74062 445074
rect 74146 444838 74382 445074
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 91826 445158 92062 445394
rect 92146 445158 92382 445394
rect 91826 444838 92062 445074
rect 92146 444838 92382 445074
rect 100826 444218 101062 444454
rect 101146 444218 101382 444454
rect 100826 443898 101062 444134
rect 101146 443898 101382 444134
rect 109826 445158 110062 445394
rect 110146 445158 110382 445394
rect 109826 444838 110062 445074
rect 110146 444838 110382 445074
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 127826 445158 128062 445394
rect 128146 445158 128382 445394
rect 127826 444838 128062 445074
rect 128146 444838 128382 445074
rect 136826 444218 137062 444454
rect 137146 444218 137382 444454
rect 136826 443898 137062 444134
rect 137146 443898 137382 444134
rect 145826 445158 146062 445394
rect 146146 445158 146382 445394
rect 145826 444838 146062 445074
rect 146146 444838 146382 445074
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 163826 445158 164062 445394
rect 164146 445158 164382 445394
rect 163826 444838 164062 445074
rect 164146 444838 164382 445074
rect 172826 444218 173062 444454
rect 173146 444218 173382 444454
rect 172826 443898 173062 444134
rect 173146 443898 173382 444134
rect 181826 445158 182062 445394
rect 182146 445158 182382 445394
rect 181826 444838 182062 445074
rect 182146 444838 182382 445074
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 199826 445158 200062 445394
rect 200146 445158 200382 445394
rect 199826 444838 200062 445074
rect 200146 444838 200382 445074
rect 208826 444218 209062 444454
rect 209146 444218 209382 444454
rect 208826 443898 209062 444134
rect 209146 443898 209382 444134
rect 217826 445158 218062 445394
rect 218146 445158 218382 445394
rect 217826 444838 218062 445074
rect 218146 444838 218382 445074
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 235826 445158 236062 445394
rect 236146 445158 236382 445394
rect 235826 444838 236062 445074
rect 236146 444838 236382 445074
rect 244826 444218 245062 444454
rect 245146 444218 245382 444454
rect 244826 443898 245062 444134
rect 245146 443898 245382 444134
rect 253826 445158 254062 445394
rect 254146 445158 254382 445394
rect 253826 444838 254062 445074
rect 254146 444838 254382 445074
rect 262826 444218 263062 444454
rect 263146 444218 263382 444454
rect 262826 443898 263062 444134
rect 263146 443898 263382 444134
rect 271826 445158 272062 445394
rect 272146 445158 272382 445394
rect 271826 444838 272062 445074
rect 272146 444838 272382 445074
rect 280826 444218 281062 444454
rect 281146 444218 281382 444454
rect 280826 443898 281062 444134
rect 281146 443898 281382 444134
rect 289826 445158 290062 445394
rect 290146 445158 290382 445394
rect 289826 444838 290062 445074
rect 290146 444838 290382 445074
rect 298826 444218 299062 444454
rect 299146 444218 299382 444454
rect 298826 443898 299062 444134
rect 299146 443898 299382 444134
rect 307826 445158 308062 445394
rect 308146 445158 308382 445394
rect 307826 444838 308062 445074
rect 308146 444838 308382 445074
rect 316826 444218 317062 444454
rect 317146 444218 317382 444454
rect 316826 443898 317062 444134
rect 317146 443898 317382 444134
rect 325826 445158 326062 445394
rect 326146 445158 326382 445394
rect 325826 444838 326062 445074
rect 326146 444838 326382 445074
rect 334826 444218 335062 444454
rect 335146 444218 335382 444454
rect 334826 443898 335062 444134
rect 335146 443898 335382 444134
rect 343826 445158 344062 445394
rect 344146 445158 344382 445394
rect 343826 444838 344062 445074
rect 344146 444838 344382 445074
rect 352826 444218 353062 444454
rect 353146 444218 353382 444454
rect 352826 443898 353062 444134
rect 353146 443898 353382 444134
rect 361826 445158 362062 445394
rect 362146 445158 362382 445394
rect 361826 444838 362062 445074
rect 362146 444838 362382 445074
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 379826 445158 380062 445394
rect 380146 445158 380382 445394
rect 379826 444838 380062 445074
rect 380146 444838 380382 445074
rect 388826 444218 389062 444454
rect 389146 444218 389382 444454
rect 388826 443898 389062 444134
rect 389146 443898 389382 444134
rect 397826 445158 398062 445394
rect 398146 445158 398382 445394
rect 397826 444838 398062 445074
rect 398146 444838 398382 445074
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 415826 445158 416062 445394
rect 416146 445158 416382 445394
rect 415826 444838 416062 445074
rect 416146 444838 416382 445074
rect 424826 444218 425062 444454
rect 425146 444218 425382 444454
rect 424826 443898 425062 444134
rect 425146 443898 425382 444134
rect 433826 445158 434062 445394
rect 434146 445158 434382 445394
rect 433826 444838 434062 445074
rect 434146 444838 434382 445074
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 451826 445158 452062 445394
rect 452146 445158 452382 445394
rect 451826 444838 452062 445074
rect 452146 444838 452382 445074
rect 460826 444218 461062 444454
rect 461146 444218 461382 444454
rect 460826 443898 461062 444134
rect 461146 443898 461382 444134
rect 469826 445158 470062 445394
rect 470146 445158 470382 445394
rect 469826 444838 470062 445074
rect 470146 444838 470382 445074
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 487826 445158 488062 445394
rect 488146 445158 488382 445394
rect 487826 444838 488062 445074
rect 488146 444838 488382 445074
rect 496826 444218 497062 444454
rect 497146 444218 497382 444454
rect 496826 443898 497062 444134
rect 497146 443898 497382 444134
rect 505826 445158 506062 445394
rect 506146 445158 506382 445394
rect 505826 444838 506062 445074
rect 506146 444838 506382 445074
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 523826 445158 524062 445394
rect 524146 445158 524382 445394
rect 523826 444838 524062 445074
rect 524146 444838 524382 445074
rect 532826 444218 533062 444454
rect 533146 444218 533382 444454
rect 532826 443898 533062 444134
rect 533146 443898 533382 444134
rect 541826 445158 542062 445394
rect 542146 445158 542382 445394
rect 541826 444838 542062 445074
rect 542146 444838 542382 445074
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 19952 435218 20188 435454
rect 19952 434898 20188 435134
rect 25882 435218 26118 435454
rect 25882 434898 26118 435134
rect 31813 435218 32049 435454
rect 31813 434898 32049 435134
rect 46952 435218 47188 435454
rect 46952 434898 47188 435134
rect 52882 435218 53118 435454
rect 52882 434898 53118 435134
rect 58813 435218 59049 435454
rect 58813 434898 59049 435134
rect 73952 435218 74188 435454
rect 73952 434898 74188 435134
rect 79882 435218 80118 435454
rect 79882 434898 80118 435134
rect 85813 435218 86049 435454
rect 85813 434898 86049 435134
rect 100952 435218 101188 435454
rect 100952 434898 101188 435134
rect 106882 435218 107118 435454
rect 106882 434898 107118 435134
rect 112813 435218 113049 435454
rect 112813 434898 113049 435134
rect 127952 435218 128188 435454
rect 127952 434898 128188 435134
rect 133882 435218 134118 435454
rect 133882 434898 134118 435134
rect 139813 435218 140049 435454
rect 139813 434898 140049 435134
rect 154952 435218 155188 435454
rect 154952 434898 155188 435134
rect 160882 435218 161118 435454
rect 160882 434898 161118 435134
rect 166813 435218 167049 435454
rect 166813 434898 167049 435134
rect 181952 435218 182188 435454
rect 181952 434898 182188 435134
rect 187882 435218 188118 435454
rect 187882 434898 188118 435134
rect 193813 435218 194049 435454
rect 193813 434898 194049 435134
rect 208952 435218 209188 435454
rect 208952 434898 209188 435134
rect 214882 435218 215118 435454
rect 214882 434898 215118 435134
rect 220813 435218 221049 435454
rect 220813 434898 221049 435134
rect 235952 435218 236188 435454
rect 235952 434898 236188 435134
rect 241882 435218 242118 435454
rect 241882 434898 242118 435134
rect 247813 435218 248049 435454
rect 247813 434898 248049 435134
rect 262952 435218 263188 435454
rect 262952 434898 263188 435134
rect 268882 435218 269118 435454
rect 268882 434898 269118 435134
rect 274813 435218 275049 435454
rect 274813 434898 275049 435134
rect 289952 435218 290188 435454
rect 289952 434898 290188 435134
rect 295882 435218 296118 435454
rect 295882 434898 296118 435134
rect 301813 435218 302049 435454
rect 301813 434898 302049 435134
rect 316952 435218 317188 435454
rect 316952 434898 317188 435134
rect 322882 435218 323118 435454
rect 322882 434898 323118 435134
rect 328813 435218 329049 435454
rect 328813 434898 329049 435134
rect 343952 435218 344188 435454
rect 343952 434898 344188 435134
rect 349882 435218 350118 435454
rect 349882 434898 350118 435134
rect 355813 435218 356049 435454
rect 355813 434898 356049 435134
rect 370952 435218 371188 435454
rect 370952 434898 371188 435134
rect 376882 435218 377118 435454
rect 376882 434898 377118 435134
rect 382813 435218 383049 435454
rect 382813 434898 383049 435134
rect 397952 435218 398188 435454
rect 397952 434898 398188 435134
rect 403882 435218 404118 435454
rect 403882 434898 404118 435134
rect 409813 435218 410049 435454
rect 409813 434898 410049 435134
rect 424952 435218 425188 435454
rect 424952 434898 425188 435134
rect 430882 435218 431118 435454
rect 430882 434898 431118 435134
rect 436813 435218 437049 435454
rect 436813 434898 437049 435134
rect 451952 435218 452188 435454
rect 451952 434898 452188 435134
rect 457882 435218 458118 435454
rect 457882 434898 458118 435134
rect 463813 435218 464049 435454
rect 463813 434898 464049 435134
rect 478952 435218 479188 435454
rect 478952 434898 479188 435134
rect 484882 435218 485118 435454
rect 484882 434898 485118 435134
rect 490813 435218 491049 435454
rect 490813 434898 491049 435134
rect 505952 435218 506188 435454
rect 505952 434898 506188 435134
rect 511882 435218 512118 435454
rect 511882 434898 512118 435134
rect 517813 435218 518049 435454
rect 517813 434898 518049 435134
rect 532952 435218 533188 435454
rect 532952 434898 533188 435134
rect 538882 435218 539118 435454
rect 538882 434898 539118 435134
rect 544813 435218 545049 435454
rect 544813 434898 545049 435134
rect 559826 435218 560062 435454
rect 560146 435218 560382 435454
rect 559826 434898 560062 435134
rect 560146 434898 560382 435134
rect 10826 426218 11062 426454
rect 11146 426218 11382 426454
rect 10826 425898 11062 426134
rect 11146 425898 11382 426134
rect 22916 426218 23152 426454
rect 22916 425898 23152 426134
rect 28847 426218 29083 426454
rect 28847 425898 29083 426134
rect 49916 426218 50152 426454
rect 49916 425898 50152 426134
rect 55847 426218 56083 426454
rect 55847 425898 56083 426134
rect 76916 426218 77152 426454
rect 76916 425898 77152 426134
rect 82847 426218 83083 426454
rect 82847 425898 83083 426134
rect 103916 426218 104152 426454
rect 103916 425898 104152 426134
rect 109847 426218 110083 426454
rect 109847 425898 110083 426134
rect 130916 426218 131152 426454
rect 130916 425898 131152 426134
rect 136847 426218 137083 426454
rect 136847 425898 137083 426134
rect 157916 426218 158152 426454
rect 157916 425898 158152 426134
rect 163847 426218 164083 426454
rect 163847 425898 164083 426134
rect 184916 426218 185152 426454
rect 184916 425898 185152 426134
rect 190847 426218 191083 426454
rect 190847 425898 191083 426134
rect 211916 426218 212152 426454
rect 211916 425898 212152 426134
rect 217847 426218 218083 426454
rect 217847 425898 218083 426134
rect 238916 426218 239152 426454
rect 238916 425898 239152 426134
rect 244847 426218 245083 426454
rect 244847 425898 245083 426134
rect 265916 426218 266152 426454
rect 265916 425898 266152 426134
rect 271847 426218 272083 426454
rect 271847 425898 272083 426134
rect 292916 426218 293152 426454
rect 292916 425898 293152 426134
rect 298847 426218 299083 426454
rect 298847 425898 299083 426134
rect 319916 426218 320152 426454
rect 319916 425898 320152 426134
rect 325847 426218 326083 426454
rect 325847 425898 326083 426134
rect 346916 426218 347152 426454
rect 346916 425898 347152 426134
rect 352847 426218 353083 426454
rect 352847 425898 353083 426134
rect 373916 426218 374152 426454
rect 373916 425898 374152 426134
rect 379847 426218 380083 426454
rect 379847 425898 380083 426134
rect 400916 426218 401152 426454
rect 400916 425898 401152 426134
rect 406847 426218 407083 426454
rect 406847 425898 407083 426134
rect 427916 426218 428152 426454
rect 427916 425898 428152 426134
rect 433847 426218 434083 426454
rect 433847 425898 434083 426134
rect 454916 426218 455152 426454
rect 454916 425898 455152 426134
rect 460847 426218 461083 426454
rect 460847 425898 461083 426134
rect 481916 426218 482152 426454
rect 481916 425898 482152 426134
rect 487847 426218 488083 426454
rect 487847 425898 488083 426134
rect 508916 426218 509152 426454
rect 508916 425898 509152 426134
rect 514847 426218 515083 426454
rect 514847 425898 515083 426134
rect 535916 426218 536152 426454
rect 535916 425898 536152 426134
rect 541847 426218 542083 426454
rect 541847 425898 542083 426134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 28826 418158 29062 418394
rect 29146 418158 29382 418394
rect 28826 417838 29062 418074
rect 29146 417838 29382 418074
rect 37826 417218 38062 417454
rect 38146 417218 38382 417454
rect 37826 416898 38062 417134
rect 38146 416898 38382 417134
rect 46826 418158 47062 418394
rect 47146 418158 47382 418394
rect 46826 417838 47062 418074
rect 47146 417838 47382 418074
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 64826 418158 65062 418394
rect 65146 418158 65382 418394
rect 64826 417838 65062 418074
rect 65146 417838 65382 418074
rect 73826 417218 74062 417454
rect 74146 417218 74382 417454
rect 73826 416898 74062 417134
rect 74146 416898 74382 417134
rect 82826 418158 83062 418394
rect 83146 418158 83382 418394
rect 82826 417838 83062 418074
rect 83146 417838 83382 418074
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 100826 418158 101062 418394
rect 101146 418158 101382 418394
rect 100826 417838 101062 418074
rect 101146 417838 101382 418074
rect 109826 417218 110062 417454
rect 110146 417218 110382 417454
rect 109826 416898 110062 417134
rect 110146 416898 110382 417134
rect 118826 418158 119062 418394
rect 119146 418158 119382 418394
rect 118826 417838 119062 418074
rect 119146 417838 119382 418074
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 136826 418158 137062 418394
rect 137146 418158 137382 418394
rect 136826 417838 137062 418074
rect 137146 417838 137382 418074
rect 145826 417218 146062 417454
rect 146146 417218 146382 417454
rect 145826 416898 146062 417134
rect 146146 416898 146382 417134
rect 154826 418158 155062 418394
rect 155146 418158 155382 418394
rect 154826 417838 155062 418074
rect 155146 417838 155382 418074
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 172826 418158 173062 418394
rect 173146 418158 173382 418394
rect 172826 417838 173062 418074
rect 173146 417838 173382 418074
rect 181826 417218 182062 417454
rect 182146 417218 182382 417454
rect 181826 416898 182062 417134
rect 182146 416898 182382 417134
rect 190826 418158 191062 418394
rect 191146 418158 191382 418394
rect 190826 417838 191062 418074
rect 191146 417838 191382 418074
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 208826 418158 209062 418394
rect 209146 418158 209382 418394
rect 208826 417838 209062 418074
rect 209146 417838 209382 418074
rect 217826 417218 218062 417454
rect 218146 417218 218382 417454
rect 217826 416898 218062 417134
rect 218146 416898 218382 417134
rect 226826 418158 227062 418394
rect 227146 418158 227382 418394
rect 226826 417838 227062 418074
rect 227146 417838 227382 418074
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 244826 418158 245062 418394
rect 245146 418158 245382 418394
rect 244826 417838 245062 418074
rect 245146 417838 245382 418074
rect 253826 417218 254062 417454
rect 254146 417218 254382 417454
rect 253826 416898 254062 417134
rect 254146 416898 254382 417134
rect 262826 418158 263062 418394
rect 263146 418158 263382 418394
rect 262826 417838 263062 418074
rect 263146 417838 263382 418074
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 280826 418158 281062 418394
rect 281146 418158 281382 418394
rect 280826 417838 281062 418074
rect 281146 417838 281382 418074
rect 289826 417218 290062 417454
rect 290146 417218 290382 417454
rect 289826 416898 290062 417134
rect 290146 416898 290382 417134
rect 298826 418158 299062 418394
rect 299146 418158 299382 418394
rect 298826 417838 299062 418074
rect 299146 417838 299382 418074
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 316826 418158 317062 418394
rect 317146 418158 317382 418394
rect 316826 417838 317062 418074
rect 317146 417838 317382 418074
rect 325826 417218 326062 417454
rect 326146 417218 326382 417454
rect 325826 416898 326062 417134
rect 326146 416898 326382 417134
rect 334826 418158 335062 418394
rect 335146 418158 335382 418394
rect 334826 417838 335062 418074
rect 335146 417838 335382 418074
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 352826 418158 353062 418394
rect 353146 418158 353382 418394
rect 352826 417838 353062 418074
rect 353146 417838 353382 418074
rect 361826 417218 362062 417454
rect 362146 417218 362382 417454
rect 361826 416898 362062 417134
rect 362146 416898 362382 417134
rect 370826 418158 371062 418394
rect 371146 418158 371382 418394
rect 370826 417838 371062 418074
rect 371146 417838 371382 418074
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 388826 418158 389062 418394
rect 389146 418158 389382 418394
rect 388826 417838 389062 418074
rect 389146 417838 389382 418074
rect 397826 417218 398062 417454
rect 398146 417218 398382 417454
rect 397826 416898 398062 417134
rect 398146 416898 398382 417134
rect 406826 418158 407062 418394
rect 407146 418158 407382 418394
rect 406826 417838 407062 418074
rect 407146 417838 407382 418074
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 424826 418158 425062 418394
rect 425146 418158 425382 418394
rect 424826 417838 425062 418074
rect 425146 417838 425382 418074
rect 433826 417218 434062 417454
rect 434146 417218 434382 417454
rect 433826 416898 434062 417134
rect 434146 416898 434382 417134
rect 442826 418158 443062 418394
rect 443146 418158 443382 418394
rect 442826 417838 443062 418074
rect 443146 417838 443382 418074
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 460826 418158 461062 418394
rect 461146 418158 461382 418394
rect 460826 417838 461062 418074
rect 461146 417838 461382 418074
rect 469826 417218 470062 417454
rect 470146 417218 470382 417454
rect 469826 416898 470062 417134
rect 470146 416898 470382 417134
rect 478826 418158 479062 418394
rect 479146 418158 479382 418394
rect 478826 417838 479062 418074
rect 479146 417838 479382 418074
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 496826 418158 497062 418394
rect 497146 418158 497382 418394
rect 496826 417838 497062 418074
rect 497146 417838 497382 418074
rect 505826 417218 506062 417454
rect 506146 417218 506382 417454
rect 505826 416898 506062 417134
rect 506146 416898 506382 417134
rect 514826 418158 515062 418394
rect 515146 418158 515382 418394
rect 514826 417838 515062 418074
rect 515146 417838 515382 418074
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 532826 418158 533062 418394
rect 533146 418158 533382 418394
rect 532826 417838 533062 418074
rect 533146 417838 533382 418074
rect 541826 417218 542062 417454
rect 542146 417218 542382 417454
rect 541826 416898 542062 417134
rect 542146 416898 542382 417134
rect 550826 418158 551062 418394
rect 551146 418158 551382 418394
rect 550826 417838 551062 418074
rect 551146 417838 551382 418074
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 22916 408218 23152 408454
rect 22916 407898 23152 408134
rect 28847 408218 29083 408454
rect 28847 407898 29083 408134
rect 49916 408218 50152 408454
rect 49916 407898 50152 408134
rect 55847 408218 56083 408454
rect 55847 407898 56083 408134
rect 76916 408218 77152 408454
rect 76916 407898 77152 408134
rect 82847 408218 83083 408454
rect 82847 407898 83083 408134
rect 103916 408218 104152 408454
rect 103916 407898 104152 408134
rect 109847 408218 110083 408454
rect 109847 407898 110083 408134
rect 130916 408218 131152 408454
rect 130916 407898 131152 408134
rect 136847 408218 137083 408454
rect 136847 407898 137083 408134
rect 157916 408218 158152 408454
rect 157916 407898 158152 408134
rect 163847 408218 164083 408454
rect 163847 407898 164083 408134
rect 184916 408218 185152 408454
rect 184916 407898 185152 408134
rect 190847 408218 191083 408454
rect 190847 407898 191083 408134
rect 211916 408218 212152 408454
rect 211916 407898 212152 408134
rect 217847 408218 218083 408454
rect 217847 407898 218083 408134
rect 238916 408218 239152 408454
rect 238916 407898 239152 408134
rect 244847 408218 245083 408454
rect 244847 407898 245083 408134
rect 265916 408218 266152 408454
rect 265916 407898 266152 408134
rect 271847 408218 272083 408454
rect 271847 407898 272083 408134
rect 292916 408218 293152 408454
rect 292916 407898 293152 408134
rect 298847 408218 299083 408454
rect 298847 407898 299083 408134
rect 319916 408218 320152 408454
rect 319916 407898 320152 408134
rect 325847 408218 326083 408454
rect 325847 407898 326083 408134
rect 346916 408218 347152 408454
rect 346916 407898 347152 408134
rect 352847 408218 353083 408454
rect 352847 407898 353083 408134
rect 373916 408218 374152 408454
rect 373916 407898 374152 408134
rect 379847 408218 380083 408454
rect 379847 407898 380083 408134
rect 400916 408218 401152 408454
rect 400916 407898 401152 408134
rect 406847 408218 407083 408454
rect 406847 407898 407083 408134
rect 427916 408218 428152 408454
rect 427916 407898 428152 408134
rect 433847 408218 434083 408454
rect 433847 407898 434083 408134
rect 454916 408218 455152 408454
rect 454916 407898 455152 408134
rect 460847 408218 461083 408454
rect 460847 407898 461083 408134
rect 481916 408218 482152 408454
rect 481916 407898 482152 408134
rect 487847 408218 488083 408454
rect 487847 407898 488083 408134
rect 508916 408218 509152 408454
rect 508916 407898 509152 408134
rect 514847 408218 515083 408454
rect 514847 407898 515083 408134
rect 535916 408218 536152 408454
rect 535916 407898 536152 408134
rect 541847 408218 542083 408454
rect 541847 407898 542083 408134
rect 19952 399218 20188 399454
rect 19952 398898 20188 399134
rect 25882 399218 26118 399454
rect 25882 398898 26118 399134
rect 31813 399218 32049 399454
rect 31813 398898 32049 399134
rect 46952 399218 47188 399454
rect 46952 398898 47188 399134
rect 52882 399218 53118 399454
rect 52882 398898 53118 399134
rect 58813 399218 59049 399454
rect 58813 398898 59049 399134
rect 73952 399218 74188 399454
rect 73952 398898 74188 399134
rect 79882 399218 80118 399454
rect 79882 398898 80118 399134
rect 85813 399218 86049 399454
rect 85813 398898 86049 399134
rect 100952 399218 101188 399454
rect 100952 398898 101188 399134
rect 106882 399218 107118 399454
rect 106882 398898 107118 399134
rect 112813 399218 113049 399454
rect 112813 398898 113049 399134
rect 127952 399218 128188 399454
rect 127952 398898 128188 399134
rect 133882 399218 134118 399454
rect 133882 398898 134118 399134
rect 139813 399218 140049 399454
rect 139813 398898 140049 399134
rect 154952 399218 155188 399454
rect 154952 398898 155188 399134
rect 160882 399218 161118 399454
rect 160882 398898 161118 399134
rect 166813 399218 167049 399454
rect 166813 398898 167049 399134
rect 181952 399218 182188 399454
rect 181952 398898 182188 399134
rect 187882 399218 188118 399454
rect 187882 398898 188118 399134
rect 193813 399218 194049 399454
rect 193813 398898 194049 399134
rect 208952 399218 209188 399454
rect 208952 398898 209188 399134
rect 214882 399218 215118 399454
rect 214882 398898 215118 399134
rect 220813 399218 221049 399454
rect 220813 398898 221049 399134
rect 235952 399218 236188 399454
rect 235952 398898 236188 399134
rect 241882 399218 242118 399454
rect 241882 398898 242118 399134
rect 247813 399218 248049 399454
rect 247813 398898 248049 399134
rect 262952 399218 263188 399454
rect 262952 398898 263188 399134
rect 268882 399218 269118 399454
rect 268882 398898 269118 399134
rect 274813 399218 275049 399454
rect 274813 398898 275049 399134
rect 289952 399218 290188 399454
rect 289952 398898 290188 399134
rect 295882 399218 296118 399454
rect 295882 398898 296118 399134
rect 301813 399218 302049 399454
rect 301813 398898 302049 399134
rect 316952 399218 317188 399454
rect 316952 398898 317188 399134
rect 322882 399218 323118 399454
rect 322882 398898 323118 399134
rect 328813 399218 329049 399454
rect 328813 398898 329049 399134
rect 343952 399218 344188 399454
rect 343952 398898 344188 399134
rect 349882 399218 350118 399454
rect 349882 398898 350118 399134
rect 355813 399218 356049 399454
rect 355813 398898 356049 399134
rect 370952 399218 371188 399454
rect 370952 398898 371188 399134
rect 376882 399218 377118 399454
rect 376882 398898 377118 399134
rect 382813 399218 383049 399454
rect 382813 398898 383049 399134
rect 397952 399218 398188 399454
rect 397952 398898 398188 399134
rect 403882 399218 404118 399454
rect 403882 398898 404118 399134
rect 409813 399218 410049 399454
rect 409813 398898 410049 399134
rect 424952 399218 425188 399454
rect 424952 398898 425188 399134
rect 430882 399218 431118 399454
rect 430882 398898 431118 399134
rect 436813 399218 437049 399454
rect 436813 398898 437049 399134
rect 451952 399218 452188 399454
rect 451952 398898 452188 399134
rect 457882 399218 458118 399454
rect 457882 398898 458118 399134
rect 463813 399218 464049 399454
rect 463813 398898 464049 399134
rect 478952 399218 479188 399454
rect 478952 398898 479188 399134
rect 484882 399218 485118 399454
rect 484882 398898 485118 399134
rect 490813 399218 491049 399454
rect 490813 398898 491049 399134
rect 505952 399218 506188 399454
rect 505952 398898 506188 399134
rect 511882 399218 512118 399454
rect 511882 398898 512118 399134
rect 517813 399218 518049 399454
rect 517813 398898 518049 399134
rect 532952 399218 533188 399454
rect 532952 398898 533188 399134
rect 538882 399218 539118 399454
rect 538882 398898 539118 399134
rect 544813 399218 545049 399454
rect 544813 398898 545049 399134
rect 559826 399218 560062 399454
rect 560146 399218 560382 399454
rect 559826 398898 560062 399134
rect 560146 398898 560382 399134
rect 10826 390218 11062 390454
rect 11146 390218 11382 390454
rect 10826 389898 11062 390134
rect 11146 389898 11382 390134
rect 19826 391158 20062 391394
rect 20146 391158 20382 391394
rect 19826 390838 20062 391074
rect 20146 390838 20382 391074
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 37826 391158 38062 391394
rect 38146 391158 38382 391394
rect 37826 390838 38062 391074
rect 38146 390838 38382 391074
rect 46826 390218 47062 390454
rect 47146 390218 47382 390454
rect 46826 389898 47062 390134
rect 47146 389898 47382 390134
rect 55826 391158 56062 391394
rect 56146 391158 56382 391394
rect 55826 390838 56062 391074
rect 56146 390838 56382 391074
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 73826 391158 74062 391394
rect 74146 391158 74382 391394
rect 73826 390838 74062 391074
rect 74146 390838 74382 391074
rect 82826 390218 83062 390454
rect 83146 390218 83382 390454
rect 82826 389898 83062 390134
rect 83146 389898 83382 390134
rect 91826 391158 92062 391394
rect 92146 391158 92382 391394
rect 91826 390838 92062 391074
rect 92146 390838 92382 391074
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 109826 391158 110062 391394
rect 110146 391158 110382 391394
rect 109826 390838 110062 391074
rect 110146 390838 110382 391074
rect 118826 390218 119062 390454
rect 119146 390218 119382 390454
rect 118826 389898 119062 390134
rect 119146 389898 119382 390134
rect 127826 391158 128062 391394
rect 128146 391158 128382 391394
rect 127826 390838 128062 391074
rect 128146 390838 128382 391074
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 145826 391158 146062 391394
rect 146146 391158 146382 391394
rect 145826 390838 146062 391074
rect 146146 390838 146382 391074
rect 154826 390218 155062 390454
rect 155146 390218 155382 390454
rect 154826 389898 155062 390134
rect 155146 389898 155382 390134
rect 163826 391158 164062 391394
rect 164146 391158 164382 391394
rect 163826 390838 164062 391074
rect 164146 390838 164382 391074
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 181826 391158 182062 391394
rect 182146 391158 182382 391394
rect 181826 390838 182062 391074
rect 182146 390838 182382 391074
rect 190826 390218 191062 390454
rect 191146 390218 191382 390454
rect 190826 389898 191062 390134
rect 191146 389898 191382 390134
rect 199826 391158 200062 391394
rect 200146 391158 200382 391394
rect 199826 390838 200062 391074
rect 200146 390838 200382 391074
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 217826 391158 218062 391394
rect 218146 391158 218382 391394
rect 217826 390838 218062 391074
rect 218146 390838 218382 391074
rect 226826 390218 227062 390454
rect 227146 390218 227382 390454
rect 226826 389898 227062 390134
rect 227146 389898 227382 390134
rect 235826 391158 236062 391394
rect 236146 391158 236382 391394
rect 235826 390838 236062 391074
rect 236146 390838 236382 391074
rect 244826 390218 245062 390454
rect 245146 390218 245382 390454
rect 244826 389898 245062 390134
rect 245146 389898 245382 390134
rect 253826 391158 254062 391394
rect 254146 391158 254382 391394
rect 253826 390838 254062 391074
rect 254146 390838 254382 391074
rect 262826 390218 263062 390454
rect 263146 390218 263382 390454
rect 262826 389898 263062 390134
rect 263146 389898 263382 390134
rect 271826 391158 272062 391394
rect 272146 391158 272382 391394
rect 271826 390838 272062 391074
rect 272146 390838 272382 391074
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 289826 391158 290062 391394
rect 290146 391158 290382 391394
rect 289826 390838 290062 391074
rect 290146 390838 290382 391074
rect 298826 390218 299062 390454
rect 299146 390218 299382 390454
rect 298826 389898 299062 390134
rect 299146 389898 299382 390134
rect 307826 391158 308062 391394
rect 308146 391158 308382 391394
rect 307826 390838 308062 391074
rect 308146 390838 308382 391074
rect 316826 390218 317062 390454
rect 317146 390218 317382 390454
rect 316826 389898 317062 390134
rect 317146 389898 317382 390134
rect 325826 391158 326062 391394
rect 326146 391158 326382 391394
rect 325826 390838 326062 391074
rect 326146 390838 326382 391074
rect 334826 390218 335062 390454
rect 335146 390218 335382 390454
rect 334826 389898 335062 390134
rect 335146 389898 335382 390134
rect 343826 391158 344062 391394
rect 344146 391158 344382 391394
rect 343826 390838 344062 391074
rect 344146 390838 344382 391074
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 361826 391158 362062 391394
rect 362146 391158 362382 391394
rect 361826 390838 362062 391074
rect 362146 390838 362382 391074
rect 370826 390218 371062 390454
rect 371146 390218 371382 390454
rect 370826 389898 371062 390134
rect 371146 389898 371382 390134
rect 379826 391158 380062 391394
rect 380146 391158 380382 391394
rect 379826 390838 380062 391074
rect 380146 390838 380382 391074
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 397826 391158 398062 391394
rect 398146 391158 398382 391394
rect 397826 390838 398062 391074
rect 398146 390838 398382 391074
rect 406826 390218 407062 390454
rect 407146 390218 407382 390454
rect 406826 389898 407062 390134
rect 407146 389898 407382 390134
rect 415826 391158 416062 391394
rect 416146 391158 416382 391394
rect 415826 390838 416062 391074
rect 416146 390838 416382 391074
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 433826 391158 434062 391394
rect 434146 391158 434382 391394
rect 433826 390838 434062 391074
rect 434146 390838 434382 391074
rect 442826 390218 443062 390454
rect 443146 390218 443382 390454
rect 442826 389898 443062 390134
rect 443146 389898 443382 390134
rect 451826 391158 452062 391394
rect 452146 391158 452382 391394
rect 451826 390838 452062 391074
rect 452146 390838 452382 391074
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 469826 391158 470062 391394
rect 470146 391158 470382 391394
rect 469826 390838 470062 391074
rect 470146 390838 470382 391074
rect 478826 390218 479062 390454
rect 479146 390218 479382 390454
rect 478826 389898 479062 390134
rect 479146 389898 479382 390134
rect 487826 391158 488062 391394
rect 488146 391158 488382 391394
rect 487826 390838 488062 391074
rect 488146 390838 488382 391074
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 505826 391158 506062 391394
rect 506146 391158 506382 391394
rect 505826 390838 506062 391074
rect 506146 390838 506382 391074
rect 514826 390218 515062 390454
rect 515146 390218 515382 390454
rect 514826 389898 515062 390134
rect 515146 389898 515382 390134
rect 523826 391158 524062 391394
rect 524146 391158 524382 391394
rect 523826 390838 524062 391074
rect 524146 390838 524382 391074
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 541826 391158 542062 391394
rect 542146 391158 542382 391394
rect 541826 390838 542062 391074
rect 542146 390838 542382 391074
rect 550826 390218 551062 390454
rect 551146 390218 551382 390454
rect 550826 389898 551062 390134
rect 551146 389898 551382 390134
rect 19952 381218 20188 381454
rect 19952 380898 20188 381134
rect 25882 381218 26118 381454
rect 25882 380898 26118 381134
rect 31813 381218 32049 381454
rect 31813 380898 32049 381134
rect 46952 381218 47188 381454
rect 46952 380898 47188 381134
rect 52882 381218 53118 381454
rect 52882 380898 53118 381134
rect 58813 381218 59049 381454
rect 58813 380898 59049 381134
rect 73952 381218 74188 381454
rect 73952 380898 74188 381134
rect 79882 381218 80118 381454
rect 79882 380898 80118 381134
rect 85813 381218 86049 381454
rect 85813 380898 86049 381134
rect 100952 381218 101188 381454
rect 100952 380898 101188 381134
rect 106882 381218 107118 381454
rect 106882 380898 107118 381134
rect 112813 381218 113049 381454
rect 112813 380898 113049 381134
rect 127952 381218 128188 381454
rect 127952 380898 128188 381134
rect 133882 381218 134118 381454
rect 133882 380898 134118 381134
rect 139813 381218 140049 381454
rect 139813 380898 140049 381134
rect 154952 381218 155188 381454
rect 154952 380898 155188 381134
rect 160882 381218 161118 381454
rect 160882 380898 161118 381134
rect 166813 381218 167049 381454
rect 166813 380898 167049 381134
rect 181952 381218 182188 381454
rect 181952 380898 182188 381134
rect 187882 381218 188118 381454
rect 187882 380898 188118 381134
rect 193813 381218 194049 381454
rect 193813 380898 194049 381134
rect 208952 381218 209188 381454
rect 208952 380898 209188 381134
rect 214882 381218 215118 381454
rect 214882 380898 215118 381134
rect 220813 381218 221049 381454
rect 220813 380898 221049 381134
rect 235952 381218 236188 381454
rect 235952 380898 236188 381134
rect 241882 381218 242118 381454
rect 241882 380898 242118 381134
rect 247813 381218 248049 381454
rect 247813 380898 248049 381134
rect 262952 381218 263188 381454
rect 262952 380898 263188 381134
rect 268882 381218 269118 381454
rect 268882 380898 269118 381134
rect 274813 381218 275049 381454
rect 274813 380898 275049 381134
rect 289952 381218 290188 381454
rect 289952 380898 290188 381134
rect 295882 381218 296118 381454
rect 295882 380898 296118 381134
rect 301813 381218 302049 381454
rect 301813 380898 302049 381134
rect 316952 381218 317188 381454
rect 316952 380898 317188 381134
rect 322882 381218 323118 381454
rect 322882 380898 323118 381134
rect 328813 381218 329049 381454
rect 328813 380898 329049 381134
rect 343952 381218 344188 381454
rect 343952 380898 344188 381134
rect 349882 381218 350118 381454
rect 349882 380898 350118 381134
rect 355813 381218 356049 381454
rect 355813 380898 356049 381134
rect 370952 381218 371188 381454
rect 370952 380898 371188 381134
rect 376882 381218 377118 381454
rect 376882 380898 377118 381134
rect 382813 381218 383049 381454
rect 382813 380898 383049 381134
rect 397952 381218 398188 381454
rect 397952 380898 398188 381134
rect 403882 381218 404118 381454
rect 403882 380898 404118 381134
rect 409813 381218 410049 381454
rect 409813 380898 410049 381134
rect 424952 381218 425188 381454
rect 424952 380898 425188 381134
rect 430882 381218 431118 381454
rect 430882 380898 431118 381134
rect 436813 381218 437049 381454
rect 436813 380898 437049 381134
rect 451952 381218 452188 381454
rect 451952 380898 452188 381134
rect 457882 381218 458118 381454
rect 457882 380898 458118 381134
rect 463813 381218 464049 381454
rect 463813 380898 464049 381134
rect 478952 381218 479188 381454
rect 478952 380898 479188 381134
rect 484882 381218 485118 381454
rect 484882 380898 485118 381134
rect 490813 381218 491049 381454
rect 490813 380898 491049 381134
rect 505952 381218 506188 381454
rect 505952 380898 506188 381134
rect 511882 381218 512118 381454
rect 511882 380898 512118 381134
rect 517813 381218 518049 381454
rect 517813 380898 518049 381134
rect 532952 381218 533188 381454
rect 532952 380898 533188 381134
rect 538882 381218 539118 381454
rect 538882 380898 539118 381134
rect 544813 381218 545049 381454
rect 544813 380898 545049 381134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 22916 372218 23152 372454
rect 22916 371898 23152 372134
rect 28847 372218 29083 372454
rect 28847 371898 29083 372134
rect 49916 372218 50152 372454
rect 49916 371898 50152 372134
rect 55847 372218 56083 372454
rect 55847 371898 56083 372134
rect 76916 372218 77152 372454
rect 76916 371898 77152 372134
rect 82847 372218 83083 372454
rect 82847 371898 83083 372134
rect 103916 372218 104152 372454
rect 103916 371898 104152 372134
rect 109847 372218 110083 372454
rect 109847 371898 110083 372134
rect 130916 372218 131152 372454
rect 130916 371898 131152 372134
rect 136847 372218 137083 372454
rect 136847 371898 137083 372134
rect 157916 372218 158152 372454
rect 157916 371898 158152 372134
rect 163847 372218 164083 372454
rect 163847 371898 164083 372134
rect 184916 372218 185152 372454
rect 184916 371898 185152 372134
rect 190847 372218 191083 372454
rect 190847 371898 191083 372134
rect 211916 372218 212152 372454
rect 211916 371898 212152 372134
rect 217847 372218 218083 372454
rect 217847 371898 218083 372134
rect 238916 372218 239152 372454
rect 238916 371898 239152 372134
rect 244847 372218 245083 372454
rect 244847 371898 245083 372134
rect 265916 372218 266152 372454
rect 265916 371898 266152 372134
rect 271847 372218 272083 372454
rect 271847 371898 272083 372134
rect 292916 372218 293152 372454
rect 292916 371898 293152 372134
rect 298847 372218 299083 372454
rect 298847 371898 299083 372134
rect 319916 372218 320152 372454
rect 319916 371898 320152 372134
rect 325847 372218 326083 372454
rect 325847 371898 326083 372134
rect 346916 372218 347152 372454
rect 346916 371898 347152 372134
rect 352847 372218 353083 372454
rect 352847 371898 353083 372134
rect 373916 372218 374152 372454
rect 373916 371898 374152 372134
rect 379847 372218 380083 372454
rect 379847 371898 380083 372134
rect 400916 372218 401152 372454
rect 400916 371898 401152 372134
rect 406847 372218 407083 372454
rect 406847 371898 407083 372134
rect 427916 372218 428152 372454
rect 427916 371898 428152 372134
rect 433847 372218 434083 372454
rect 433847 371898 434083 372134
rect 454916 372218 455152 372454
rect 454916 371898 455152 372134
rect 460847 372218 461083 372454
rect 460847 371898 461083 372134
rect 481916 372218 482152 372454
rect 481916 371898 482152 372134
rect 487847 372218 488083 372454
rect 487847 371898 488083 372134
rect 508916 372218 509152 372454
rect 508916 371898 509152 372134
rect 514847 372218 515083 372454
rect 514847 371898 515083 372134
rect 535916 372218 536152 372454
rect 535916 371898 536152 372134
rect 541847 372218 542083 372454
rect 541847 371898 542083 372134
rect 19826 363218 20062 363454
rect 20146 363218 20382 363454
rect 19826 362898 20062 363134
rect 20146 362898 20382 363134
rect 28826 364158 29062 364394
rect 29146 364158 29382 364394
rect 28826 363838 29062 364074
rect 29146 363838 29382 364074
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 46826 364158 47062 364394
rect 47146 364158 47382 364394
rect 46826 363838 47062 364074
rect 47146 363838 47382 364074
rect 55826 363218 56062 363454
rect 56146 363218 56382 363454
rect 55826 362898 56062 363134
rect 56146 362898 56382 363134
rect 64826 364158 65062 364394
rect 65146 364158 65382 364394
rect 64826 363838 65062 364074
rect 65146 363838 65382 364074
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 82826 364158 83062 364394
rect 83146 364158 83382 364394
rect 82826 363838 83062 364074
rect 83146 363838 83382 364074
rect 91826 363218 92062 363454
rect 92146 363218 92382 363454
rect 91826 362898 92062 363134
rect 92146 362898 92382 363134
rect 100826 364158 101062 364394
rect 101146 364158 101382 364394
rect 100826 363838 101062 364074
rect 101146 363838 101382 364074
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 118826 364158 119062 364394
rect 119146 364158 119382 364394
rect 118826 363838 119062 364074
rect 119146 363838 119382 364074
rect 127826 363218 128062 363454
rect 128146 363218 128382 363454
rect 127826 362898 128062 363134
rect 128146 362898 128382 363134
rect 136826 364158 137062 364394
rect 137146 364158 137382 364394
rect 136826 363838 137062 364074
rect 137146 363838 137382 364074
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 154826 364158 155062 364394
rect 155146 364158 155382 364394
rect 154826 363838 155062 364074
rect 155146 363838 155382 364074
rect 163826 363218 164062 363454
rect 164146 363218 164382 363454
rect 163826 362898 164062 363134
rect 164146 362898 164382 363134
rect 172826 364158 173062 364394
rect 173146 364158 173382 364394
rect 172826 363838 173062 364074
rect 173146 363838 173382 364074
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 190826 364158 191062 364394
rect 191146 364158 191382 364394
rect 190826 363838 191062 364074
rect 191146 363838 191382 364074
rect 199826 363218 200062 363454
rect 200146 363218 200382 363454
rect 199826 362898 200062 363134
rect 200146 362898 200382 363134
rect 208826 364158 209062 364394
rect 209146 364158 209382 364394
rect 208826 363838 209062 364074
rect 209146 363838 209382 364074
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 226826 364158 227062 364394
rect 227146 364158 227382 364394
rect 226826 363838 227062 364074
rect 227146 363838 227382 364074
rect 235826 363218 236062 363454
rect 236146 363218 236382 363454
rect 235826 362898 236062 363134
rect 236146 362898 236382 363134
rect 244826 364158 245062 364394
rect 245146 364158 245382 364394
rect 244826 363838 245062 364074
rect 245146 363838 245382 364074
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 262826 364158 263062 364394
rect 263146 364158 263382 364394
rect 262826 363838 263062 364074
rect 263146 363838 263382 364074
rect 271826 363218 272062 363454
rect 272146 363218 272382 363454
rect 271826 362898 272062 363134
rect 272146 362898 272382 363134
rect 280826 364158 281062 364394
rect 281146 364158 281382 364394
rect 280826 363838 281062 364074
rect 281146 363838 281382 364074
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 298826 364158 299062 364394
rect 299146 364158 299382 364394
rect 298826 363838 299062 364074
rect 299146 363838 299382 364074
rect 307826 363218 308062 363454
rect 308146 363218 308382 363454
rect 307826 362898 308062 363134
rect 308146 362898 308382 363134
rect 316826 364158 317062 364394
rect 317146 364158 317382 364394
rect 316826 363838 317062 364074
rect 317146 363838 317382 364074
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 334826 364158 335062 364394
rect 335146 364158 335382 364394
rect 334826 363838 335062 364074
rect 335146 363838 335382 364074
rect 343826 363218 344062 363454
rect 344146 363218 344382 363454
rect 343826 362898 344062 363134
rect 344146 362898 344382 363134
rect 352826 364158 353062 364394
rect 353146 364158 353382 364394
rect 352826 363838 353062 364074
rect 353146 363838 353382 364074
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 370826 364158 371062 364394
rect 371146 364158 371382 364394
rect 370826 363838 371062 364074
rect 371146 363838 371382 364074
rect 379826 363218 380062 363454
rect 380146 363218 380382 363454
rect 379826 362898 380062 363134
rect 380146 362898 380382 363134
rect 388826 364158 389062 364394
rect 389146 364158 389382 364394
rect 388826 363838 389062 364074
rect 389146 363838 389382 364074
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 406826 364158 407062 364394
rect 407146 364158 407382 364394
rect 406826 363838 407062 364074
rect 407146 363838 407382 364074
rect 415826 363218 416062 363454
rect 416146 363218 416382 363454
rect 415826 362898 416062 363134
rect 416146 362898 416382 363134
rect 424826 364158 425062 364394
rect 425146 364158 425382 364394
rect 424826 363838 425062 364074
rect 425146 363838 425382 364074
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 442826 364158 443062 364394
rect 443146 364158 443382 364394
rect 442826 363838 443062 364074
rect 443146 363838 443382 364074
rect 451826 363218 452062 363454
rect 452146 363218 452382 363454
rect 451826 362898 452062 363134
rect 452146 362898 452382 363134
rect 460826 364158 461062 364394
rect 461146 364158 461382 364394
rect 460826 363838 461062 364074
rect 461146 363838 461382 364074
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 478826 364158 479062 364394
rect 479146 364158 479382 364394
rect 478826 363838 479062 364074
rect 479146 363838 479382 364074
rect 487826 363218 488062 363454
rect 488146 363218 488382 363454
rect 487826 362898 488062 363134
rect 488146 362898 488382 363134
rect 496826 364158 497062 364394
rect 497146 364158 497382 364394
rect 496826 363838 497062 364074
rect 497146 363838 497382 364074
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 514826 364158 515062 364394
rect 515146 364158 515382 364394
rect 514826 363838 515062 364074
rect 515146 363838 515382 364074
rect 523826 363218 524062 363454
rect 524146 363218 524382 363454
rect 523826 362898 524062 363134
rect 524146 362898 524382 363134
rect 532826 364158 533062 364394
rect 533146 364158 533382 364394
rect 532826 363838 533062 364074
rect 533146 363838 533382 364074
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 550826 364158 551062 364394
rect 551146 364158 551382 364394
rect 550826 363838 551062 364074
rect 551146 363838 551382 364074
rect 559826 363218 560062 363454
rect 560146 363218 560382 363454
rect 559826 362898 560062 363134
rect 560146 362898 560382 363134
rect 10826 354218 11062 354454
rect 11146 354218 11382 354454
rect 10826 353898 11062 354134
rect 11146 353898 11382 354134
rect 22916 354218 23152 354454
rect 22916 353898 23152 354134
rect 28847 354218 29083 354454
rect 28847 353898 29083 354134
rect 49916 354218 50152 354454
rect 49916 353898 50152 354134
rect 55847 354218 56083 354454
rect 55847 353898 56083 354134
rect 76916 354218 77152 354454
rect 76916 353898 77152 354134
rect 82847 354218 83083 354454
rect 82847 353898 83083 354134
rect 103916 354218 104152 354454
rect 103916 353898 104152 354134
rect 109847 354218 110083 354454
rect 109847 353898 110083 354134
rect 130916 354218 131152 354454
rect 130916 353898 131152 354134
rect 136847 354218 137083 354454
rect 136847 353898 137083 354134
rect 157916 354218 158152 354454
rect 157916 353898 158152 354134
rect 163847 354218 164083 354454
rect 163847 353898 164083 354134
rect 184916 354218 185152 354454
rect 184916 353898 185152 354134
rect 190847 354218 191083 354454
rect 190847 353898 191083 354134
rect 211916 354218 212152 354454
rect 211916 353898 212152 354134
rect 217847 354218 218083 354454
rect 217847 353898 218083 354134
rect 238916 354218 239152 354454
rect 238916 353898 239152 354134
rect 244847 354218 245083 354454
rect 244847 353898 245083 354134
rect 265916 354218 266152 354454
rect 265916 353898 266152 354134
rect 271847 354218 272083 354454
rect 271847 353898 272083 354134
rect 292916 354218 293152 354454
rect 292916 353898 293152 354134
rect 298847 354218 299083 354454
rect 298847 353898 299083 354134
rect 319916 354218 320152 354454
rect 319916 353898 320152 354134
rect 325847 354218 326083 354454
rect 325847 353898 326083 354134
rect 346916 354218 347152 354454
rect 346916 353898 347152 354134
rect 352847 354218 353083 354454
rect 352847 353898 353083 354134
rect 373916 354218 374152 354454
rect 373916 353898 374152 354134
rect 379847 354218 380083 354454
rect 379847 353898 380083 354134
rect 400916 354218 401152 354454
rect 400916 353898 401152 354134
rect 406847 354218 407083 354454
rect 406847 353898 407083 354134
rect 427916 354218 428152 354454
rect 427916 353898 428152 354134
rect 433847 354218 434083 354454
rect 433847 353898 434083 354134
rect 454916 354218 455152 354454
rect 454916 353898 455152 354134
rect 460847 354218 461083 354454
rect 460847 353898 461083 354134
rect 481916 354218 482152 354454
rect 481916 353898 482152 354134
rect 487847 354218 488083 354454
rect 487847 353898 488083 354134
rect 508916 354218 509152 354454
rect 508916 353898 509152 354134
rect 514847 354218 515083 354454
rect 514847 353898 515083 354134
rect 535916 354218 536152 354454
rect 535916 353898 536152 354134
rect 541847 354218 542083 354454
rect 541847 353898 542083 354134
rect 19952 345218 20188 345454
rect 19952 344898 20188 345134
rect 25882 345218 26118 345454
rect 25882 344898 26118 345134
rect 31813 345218 32049 345454
rect 31813 344898 32049 345134
rect 46952 345218 47188 345454
rect 46952 344898 47188 345134
rect 52882 345218 53118 345454
rect 52882 344898 53118 345134
rect 58813 345218 59049 345454
rect 58813 344898 59049 345134
rect 73952 345218 74188 345454
rect 73952 344898 74188 345134
rect 79882 345218 80118 345454
rect 79882 344898 80118 345134
rect 85813 345218 86049 345454
rect 85813 344898 86049 345134
rect 100952 345218 101188 345454
rect 100952 344898 101188 345134
rect 106882 345218 107118 345454
rect 106882 344898 107118 345134
rect 112813 345218 113049 345454
rect 112813 344898 113049 345134
rect 127952 345218 128188 345454
rect 127952 344898 128188 345134
rect 133882 345218 134118 345454
rect 133882 344898 134118 345134
rect 139813 345218 140049 345454
rect 139813 344898 140049 345134
rect 154952 345218 155188 345454
rect 154952 344898 155188 345134
rect 160882 345218 161118 345454
rect 160882 344898 161118 345134
rect 166813 345218 167049 345454
rect 166813 344898 167049 345134
rect 181952 345218 182188 345454
rect 181952 344898 182188 345134
rect 187882 345218 188118 345454
rect 187882 344898 188118 345134
rect 193813 345218 194049 345454
rect 193813 344898 194049 345134
rect 208952 345218 209188 345454
rect 208952 344898 209188 345134
rect 214882 345218 215118 345454
rect 214882 344898 215118 345134
rect 220813 345218 221049 345454
rect 220813 344898 221049 345134
rect 235952 345218 236188 345454
rect 235952 344898 236188 345134
rect 241882 345218 242118 345454
rect 241882 344898 242118 345134
rect 247813 345218 248049 345454
rect 247813 344898 248049 345134
rect 262952 345218 263188 345454
rect 262952 344898 263188 345134
rect 268882 345218 269118 345454
rect 268882 344898 269118 345134
rect 274813 345218 275049 345454
rect 274813 344898 275049 345134
rect 289952 345218 290188 345454
rect 289952 344898 290188 345134
rect 295882 345218 296118 345454
rect 295882 344898 296118 345134
rect 301813 345218 302049 345454
rect 301813 344898 302049 345134
rect 316952 345218 317188 345454
rect 316952 344898 317188 345134
rect 322882 345218 323118 345454
rect 322882 344898 323118 345134
rect 328813 345218 329049 345454
rect 328813 344898 329049 345134
rect 343952 345218 344188 345454
rect 343952 344898 344188 345134
rect 349882 345218 350118 345454
rect 349882 344898 350118 345134
rect 355813 345218 356049 345454
rect 355813 344898 356049 345134
rect 370952 345218 371188 345454
rect 370952 344898 371188 345134
rect 376882 345218 377118 345454
rect 376882 344898 377118 345134
rect 382813 345218 383049 345454
rect 382813 344898 383049 345134
rect 397952 345218 398188 345454
rect 397952 344898 398188 345134
rect 403882 345218 404118 345454
rect 403882 344898 404118 345134
rect 409813 345218 410049 345454
rect 409813 344898 410049 345134
rect 424952 345218 425188 345454
rect 424952 344898 425188 345134
rect 430882 345218 431118 345454
rect 430882 344898 431118 345134
rect 436813 345218 437049 345454
rect 436813 344898 437049 345134
rect 451952 345218 452188 345454
rect 451952 344898 452188 345134
rect 457882 345218 458118 345454
rect 457882 344898 458118 345134
rect 463813 345218 464049 345454
rect 463813 344898 464049 345134
rect 478952 345218 479188 345454
rect 478952 344898 479188 345134
rect 484882 345218 485118 345454
rect 484882 344898 485118 345134
rect 490813 345218 491049 345454
rect 490813 344898 491049 345134
rect 505952 345218 506188 345454
rect 505952 344898 506188 345134
rect 511882 345218 512118 345454
rect 511882 344898 512118 345134
rect 517813 345218 518049 345454
rect 517813 344898 518049 345134
rect 532952 345218 533188 345454
rect 532952 344898 533188 345134
rect 538882 345218 539118 345454
rect 538882 344898 539118 345134
rect 544813 345218 545049 345454
rect 544813 344898 545049 345134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 19826 337158 20062 337394
rect 20146 337158 20382 337394
rect 19826 336838 20062 337074
rect 20146 336838 20382 337074
rect 28826 336218 29062 336454
rect 29146 336218 29382 336454
rect 28826 335898 29062 336134
rect 29146 335898 29382 336134
rect 37826 337158 38062 337394
rect 38146 337158 38382 337394
rect 37826 336838 38062 337074
rect 38146 336838 38382 337074
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 55826 337158 56062 337394
rect 56146 337158 56382 337394
rect 55826 336838 56062 337074
rect 56146 336838 56382 337074
rect 64826 336218 65062 336454
rect 65146 336218 65382 336454
rect 64826 335898 65062 336134
rect 65146 335898 65382 336134
rect 73826 337158 74062 337394
rect 74146 337158 74382 337394
rect 73826 336838 74062 337074
rect 74146 336838 74382 337074
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 91826 337158 92062 337394
rect 92146 337158 92382 337394
rect 91826 336838 92062 337074
rect 92146 336838 92382 337074
rect 100826 336218 101062 336454
rect 101146 336218 101382 336454
rect 100826 335898 101062 336134
rect 101146 335898 101382 336134
rect 109826 337158 110062 337394
rect 110146 337158 110382 337394
rect 109826 336838 110062 337074
rect 110146 336838 110382 337074
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 127826 337158 128062 337394
rect 128146 337158 128382 337394
rect 127826 336838 128062 337074
rect 128146 336838 128382 337074
rect 136826 336218 137062 336454
rect 137146 336218 137382 336454
rect 136826 335898 137062 336134
rect 137146 335898 137382 336134
rect 145826 337158 146062 337394
rect 146146 337158 146382 337394
rect 145826 336838 146062 337074
rect 146146 336838 146382 337074
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 163826 337158 164062 337394
rect 164146 337158 164382 337394
rect 163826 336838 164062 337074
rect 164146 336838 164382 337074
rect 172826 336218 173062 336454
rect 173146 336218 173382 336454
rect 172826 335898 173062 336134
rect 173146 335898 173382 336134
rect 181826 337158 182062 337394
rect 182146 337158 182382 337394
rect 181826 336838 182062 337074
rect 182146 336838 182382 337074
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 199826 337158 200062 337394
rect 200146 337158 200382 337394
rect 199826 336838 200062 337074
rect 200146 336838 200382 337074
rect 208826 336218 209062 336454
rect 209146 336218 209382 336454
rect 208826 335898 209062 336134
rect 209146 335898 209382 336134
rect 217826 337158 218062 337394
rect 218146 337158 218382 337394
rect 217826 336838 218062 337074
rect 218146 336838 218382 337074
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 235826 337158 236062 337394
rect 236146 337158 236382 337394
rect 235826 336838 236062 337074
rect 236146 336838 236382 337074
rect 244826 336218 245062 336454
rect 245146 336218 245382 336454
rect 244826 335898 245062 336134
rect 245146 335898 245382 336134
rect 253826 337158 254062 337394
rect 254146 337158 254382 337394
rect 253826 336838 254062 337074
rect 254146 336838 254382 337074
rect 262826 336218 263062 336454
rect 263146 336218 263382 336454
rect 262826 335898 263062 336134
rect 263146 335898 263382 336134
rect 271826 337158 272062 337394
rect 272146 337158 272382 337394
rect 271826 336838 272062 337074
rect 272146 336838 272382 337074
rect 280826 336218 281062 336454
rect 281146 336218 281382 336454
rect 280826 335898 281062 336134
rect 281146 335898 281382 336134
rect 289826 337158 290062 337394
rect 290146 337158 290382 337394
rect 289826 336838 290062 337074
rect 290146 336838 290382 337074
rect 298826 336218 299062 336454
rect 299146 336218 299382 336454
rect 298826 335898 299062 336134
rect 299146 335898 299382 336134
rect 307826 337158 308062 337394
rect 308146 337158 308382 337394
rect 307826 336838 308062 337074
rect 308146 336838 308382 337074
rect 316826 336218 317062 336454
rect 317146 336218 317382 336454
rect 316826 335898 317062 336134
rect 317146 335898 317382 336134
rect 325826 337158 326062 337394
rect 326146 337158 326382 337394
rect 325826 336838 326062 337074
rect 326146 336838 326382 337074
rect 334826 336218 335062 336454
rect 335146 336218 335382 336454
rect 334826 335898 335062 336134
rect 335146 335898 335382 336134
rect 343826 337158 344062 337394
rect 344146 337158 344382 337394
rect 343826 336838 344062 337074
rect 344146 336838 344382 337074
rect 352826 336218 353062 336454
rect 353146 336218 353382 336454
rect 352826 335898 353062 336134
rect 353146 335898 353382 336134
rect 361826 337158 362062 337394
rect 362146 337158 362382 337394
rect 361826 336838 362062 337074
rect 362146 336838 362382 337074
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 379826 337158 380062 337394
rect 380146 337158 380382 337394
rect 379826 336838 380062 337074
rect 380146 336838 380382 337074
rect 388826 336218 389062 336454
rect 389146 336218 389382 336454
rect 388826 335898 389062 336134
rect 389146 335898 389382 336134
rect 397826 337158 398062 337394
rect 398146 337158 398382 337394
rect 397826 336838 398062 337074
rect 398146 336838 398382 337074
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 415826 337158 416062 337394
rect 416146 337158 416382 337394
rect 415826 336838 416062 337074
rect 416146 336838 416382 337074
rect 424826 336218 425062 336454
rect 425146 336218 425382 336454
rect 424826 335898 425062 336134
rect 425146 335898 425382 336134
rect 433826 337158 434062 337394
rect 434146 337158 434382 337394
rect 433826 336838 434062 337074
rect 434146 336838 434382 337074
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 451826 337158 452062 337394
rect 452146 337158 452382 337394
rect 451826 336838 452062 337074
rect 452146 336838 452382 337074
rect 460826 336218 461062 336454
rect 461146 336218 461382 336454
rect 460826 335898 461062 336134
rect 461146 335898 461382 336134
rect 469826 337158 470062 337394
rect 470146 337158 470382 337394
rect 469826 336838 470062 337074
rect 470146 336838 470382 337074
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 487826 337158 488062 337394
rect 488146 337158 488382 337394
rect 487826 336838 488062 337074
rect 488146 336838 488382 337074
rect 496826 336218 497062 336454
rect 497146 336218 497382 336454
rect 496826 335898 497062 336134
rect 497146 335898 497382 336134
rect 505826 337158 506062 337394
rect 506146 337158 506382 337394
rect 505826 336838 506062 337074
rect 506146 336838 506382 337074
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 523826 337158 524062 337394
rect 524146 337158 524382 337394
rect 523826 336838 524062 337074
rect 524146 336838 524382 337074
rect 532826 336218 533062 336454
rect 533146 336218 533382 336454
rect 532826 335898 533062 336134
rect 533146 335898 533382 336134
rect 541826 337158 542062 337394
rect 542146 337158 542382 337394
rect 541826 336838 542062 337074
rect 542146 336838 542382 337074
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 19952 327218 20188 327454
rect 19952 326898 20188 327134
rect 25882 327218 26118 327454
rect 25882 326898 26118 327134
rect 31813 327218 32049 327454
rect 31813 326898 32049 327134
rect 46952 327218 47188 327454
rect 46952 326898 47188 327134
rect 52882 327218 53118 327454
rect 52882 326898 53118 327134
rect 58813 327218 59049 327454
rect 58813 326898 59049 327134
rect 73952 327218 74188 327454
rect 73952 326898 74188 327134
rect 79882 327218 80118 327454
rect 79882 326898 80118 327134
rect 85813 327218 86049 327454
rect 85813 326898 86049 327134
rect 100952 327218 101188 327454
rect 100952 326898 101188 327134
rect 106882 327218 107118 327454
rect 106882 326898 107118 327134
rect 112813 327218 113049 327454
rect 112813 326898 113049 327134
rect 127952 327218 128188 327454
rect 127952 326898 128188 327134
rect 133882 327218 134118 327454
rect 133882 326898 134118 327134
rect 139813 327218 140049 327454
rect 139813 326898 140049 327134
rect 154952 327218 155188 327454
rect 154952 326898 155188 327134
rect 160882 327218 161118 327454
rect 160882 326898 161118 327134
rect 166813 327218 167049 327454
rect 166813 326898 167049 327134
rect 181952 327218 182188 327454
rect 181952 326898 182188 327134
rect 187882 327218 188118 327454
rect 187882 326898 188118 327134
rect 193813 327218 194049 327454
rect 193813 326898 194049 327134
rect 208952 327218 209188 327454
rect 208952 326898 209188 327134
rect 214882 327218 215118 327454
rect 214882 326898 215118 327134
rect 220813 327218 221049 327454
rect 220813 326898 221049 327134
rect 235952 327218 236188 327454
rect 235952 326898 236188 327134
rect 241882 327218 242118 327454
rect 241882 326898 242118 327134
rect 247813 327218 248049 327454
rect 247813 326898 248049 327134
rect 262952 327218 263188 327454
rect 262952 326898 263188 327134
rect 268882 327218 269118 327454
rect 268882 326898 269118 327134
rect 274813 327218 275049 327454
rect 274813 326898 275049 327134
rect 289952 327218 290188 327454
rect 289952 326898 290188 327134
rect 295882 327218 296118 327454
rect 295882 326898 296118 327134
rect 301813 327218 302049 327454
rect 301813 326898 302049 327134
rect 316952 327218 317188 327454
rect 316952 326898 317188 327134
rect 322882 327218 323118 327454
rect 322882 326898 323118 327134
rect 328813 327218 329049 327454
rect 328813 326898 329049 327134
rect 343952 327218 344188 327454
rect 343952 326898 344188 327134
rect 349882 327218 350118 327454
rect 349882 326898 350118 327134
rect 355813 327218 356049 327454
rect 355813 326898 356049 327134
rect 370952 327218 371188 327454
rect 370952 326898 371188 327134
rect 376882 327218 377118 327454
rect 376882 326898 377118 327134
rect 382813 327218 383049 327454
rect 382813 326898 383049 327134
rect 397952 327218 398188 327454
rect 397952 326898 398188 327134
rect 403882 327218 404118 327454
rect 403882 326898 404118 327134
rect 409813 327218 410049 327454
rect 409813 326898 410049 327134
rect 424952 327218 425188 327454
rect 424952 326898 425188 327134
rect 430882 327218 431118 327454
rect 430882 326898 431118 327134
rect 436813 327218 437049 327454
rect 436813 326898 437049 327134
rect 451952 327218 452188 327454
rect 451952 326898 452188 327134
rect 457882 327218 458118 327454
rect 457882 326898 458118 327134
rect 463813 327218 464049 327454
rect 463813 326898 464049 327134
rect 478952 327218 479188 327454
rect 478952 326898 479188 327134
rect 484882 327218 485118 327454
rect 484882 326898 485118 327134
rect 490813 327218 491049 327454
rect 490813 326898 491049 327134
rect 505952 327218 506188 327454
rect 505952 326898 506188 327134
rect 511882 327218 512118 327454
rect 511882 326898 512118 327134
rect 517813 327218 518049 327454
rect 517813 326898 518049 327134
rect 532952 327218 533188 327454
rect 532952 326898 533188 327134
rect 538882 327218 539118 327454
rect 538882 326898 539118 327134
rect 544813 327218 545049 327454
rect 544813 326898 545049 327134
rect 559826 327218 560062 327454
rect 560146 327218 560382 327454
rect 559826 326898 560062 327134
rect 560146 326898 560382 327134
rect 10826 318218 11062 318454
rect 11146 318218 11382 318454
rect 10826 317898 11062 318134
rect 11146 317898 11382 318134
rect 22916 318218 23152 318454
rect 22916 317898 23152 318134
rect 28847 318218 29083 318454
rect 28847 317898 29083 318134
rect 49916 318218 50152 318454
rect 49916 317898 50152 318134
rect 55847 318218 56083 318454
rect 55847 317898 56083 318134
rect 76916 318218 77152 318454
rect 76916 317898 77152 318134
rect 82847 318218 83083 318454
rect 82847 317898 83083 318134
rect 103916 318218 104152 318454
rect 103916 317898 104152 318134
rect 109847 318218 110083 318454
rect 109847 317898 110083 318134
rect 130916 318218 131152 318454
rect 130916 317898 131152 318134
rect 136847 318218 137083 318454
rect 136847 317898 137083 318134
rect 157916 318218 158152 318454
rect 157916 317898 158152 318134
rect 163847 318218 164083 318454
rect 163847 317898 164083 318134
rect 184916 318218 185152 318454
rect 184916 317898 185152 318134
rect 190847 318218 191083 318454
rect 190847 317898 191083 318134
rect 211916 318218 212152 318454
rect 211916 317898 212152 318134
rect 217847 318218 218083 318454
rect 217847 317898 218083 318134
rect 238916 318218 239152 318454
rect 238916 317898 239152 318134
rect 244847 318218 245083 318454
rect 244847 317898 245083 318134
rect 265916 318218 266152 318454
rect 265916 317898 266152 318134
rect 271847 318218 272083 318454
rect 271847 317898 272083 318134
rect 292916 318218 293152 318454
rect 292916 317898 293152 318134
rect 298847 318218 299083 318454
rect 298847 317898 299083 318134
rect 319916 318218 320152 318454
rect 319916 317898 320152 318134
rect 325847 318218 326083 318454
rect 325847 317898 326083 318134
rect 346916 318218 347152 318454
rect 346916 317898 347152 318134
rect 352847 318218 353083 318454
rect 352847 317898 353083 318134
rect 373916 318218 374152 318454
rect 373916 317898 374152 318134
rect 379847 318218 380083 318454
rect 379847 317898 380083 318134
rect 400916 318218 401152 318454
rect 400916 317898 401152 318134
rect 406847 318218 407083 318454
rect 406847 317898 407083 318134
rect 427916 318218 428152 318454
rect 427916 317898 428152 318134
rect 433847 318218 434083 318454
rect 433847 317898 434083 318134
rect 454916 318218 455152 318454
rect 454916 317898 455152 318134
rect 460847 318218 461083 318454
rect 460847 317898 461083 318134
rect 481916 318218 482152 318454
rect 481916 317898 482152 318134
rect 487847 318218 488083 318454
rect 487847 317898 488083 318134
rect 508916 318218 509152 318454
rect 508916 317898 509152 318134
rect 514847 318218 515083 318454
rect 514847 317898 515083 318134
rect 535916 318218 536152 318454
rect 535916 317898 536152 318134
rect 541847 318218 542083 318454
rect 541847 317898 542083 318134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 28826 310158 29062 310394
rect 29146 310158 29382 310394
rect 28826 309838 29062 310074
rect 29146 309838 29382 310074
rect 37826 309218 38062 309454
rect 38146 309218 38382 309454
rect 37826 308898 38062 309134
rect 38146 308898 38382 309134
rect 46826 310158 47062 310394
rect 47146 310158 47382 310394
rect 46826 309838 47062 310074
rect 47146 309838 47382 310074
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 64826 310158 65062 310394
rect 65146 310158 65382 310394
rect 64826 309838 65062 310074
rect 65146 309838 65382 310074
rect 73826 309218 74062 309454
rect 74146 309218 74382 309454
rect 73826 308898 74062 309134
rect 74146 308898 74382 309134
rect 82826 310158 83062 310394
rect 83146 310158 83382 310394
rect 82826 309838 83062 310074
rect 83146 309838 83382 310074
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 100826 310158 101062 310394
rect 101146 310158 101382 310394
rect 100826 309838 101062 310074
rect 101146 309838 101382 310074
rect 109826 309218 110062 309454
rect 110146 309218 110382 309454
rect 109826 308898 110062 309134
rect 110146 308898 110382 309134
rect 118826 310158 119062 310394
rect 119146 310158 119382 310394
rect 118826 309838 119062 310074
rect 119146 309838 119382 310074
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 136826 310158 137062 310394
rect 137146 310158 137382 310394
rect 136826 309838 137062 310074
rect 137146 309838 137382 310074
rect 145826 309218 146062 309454
rect 146146 309218 146382 309454
rect 145826 308898 146062 309134
rect 146146 308898 146382 309134
rect 154826 310158 155062 310394
rect 155146 310158 155382 310394
rect 154826 309838 155062 310074
rect 155146 309838 155382 310074
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 172826 310158 173062 310394
rect 173146 310158 173382 310394
rect 172826 309838 173062 310074
rect 173146 309838 173382 310074
rect 181826 309218 182062 309454
rect 182146 309218 182382 309454
rect 181826 308898 182062 309134
rect 182146 308898 182382 309134
rect 190826 310158 191062 310394
rect 191146 310158 191382 310394
rect 190826 309838 191062 310074
rect 191146 309838 191382 310074
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 208826 310158 209062 310394
rect 209146 310158 209382 310394
rect 208826 309838 209062 310074
rect 209146 309838 209382 310074
rect 217826 309218 218062 309454
rect 218146 309218 218382 309454
rect 217826 308898 218062 309134
rect 218146 308898 218382 309134
rect 226826 310158 227062 310394
rect 227146 310158 227382 310394
rect 226826 309838 227062 310074
rect 227146 309838 227382 310074
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 244826 310158 245062 310394
rect 245146 310158 245382 310394
rect 244826 309838 245062 310074
rect 245146 309838 245382 310074
rect 253826 309218 254062 309454
rect 254146 309218 254382 309454
rect 253826 308898 254062 309134
rect 254146 308898 254382 309134
rect 262826 310158 263062 310394
rect 263146 310158 263382 310394
rect 262826 309838 263062 310074
rect 263146 309838 263382 310074
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 280826 310158 281062 310394
rect 281146 310158 281382 310394
rect 280826 309838 281062 310074
rect 281146 309838 281382 310074
rect 289826 309218 290062 309454
rect 290146 309218 290382 309454
rect 289826 308898 290062 309134
rect 290146 308898 290382 309134
rect 298826 310158 299062 310394
rect 299146 310158 299382 310394
rect 298826 309838 299062 310074
rect 299146 309838 299382 310074
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 316826 310158 317062 310394
rect 317146 310158 317382 310394
rect 316826 309838 317062 310074
rect 317146 309838 317382 310074
rect 325826 309218 326062 309454
rect 326146 309218 326382 309454
rect 325826 308898 326062 309134
rect 326146 308898 326382 309134
rect 334826 310158 335062 310394
rect 335146 310158 335382 310394
rect 334826 309838 335062 310074
rect 335146 309838 335382 310074
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 352826 310158 353062 310394
rect 353146 310158 353382 310394
rect 352826 309838 353062 310074
rect 353146 309838 353382 310074
rect 361826 309218 362062 309454
rect 362146 309218 362382 309454
rect 361826 308898 362062 309134
rect 362146 308898 362382 309134
rect 370826 310158 371062 310394
rect 371146 310158 371382 310394
rect 370826 309838 371062 310074
rect 371146 309838 371382 310074
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 388826 310158 389062 310394
rect 389146 310158 389382 310394
rect 388826 309838 389062 310074
rect 389146 309838 389382 310074
rect 397826 309218 398062 309454
rect 398146 309218 398382 309454
rect 397826 308898 398062 309134
rect 398146 308898 398382 309134
rect 406826 310158 407062 310394
rect 407146 310158 407382 310394
rect 406826 309838 407062 310074
rect 407146 309838 407382 310074
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 424826 310158 425062 310394
rect 425146 310158 425382 310394
rect 424826 309838 425062 310074
rect 425146 309838 425382 310074
rect 433826 309218 434062 309454
rect 434146 309218 434382 309454
rect 433826 308898 434062 309134
rect 434146 308898 434382 309134
rect 442826 310158 443062 310394
rect 443146 310158 443382 310394
rect 442826 309838 443062 310074
rect 443146 309838 443382 310074
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 460826 310158 461062 310394
rect 461146 310158 461382 310394
rect 460826 309838 461062 310074
rect 461146 309838 461382 310074
rect 469826 309218 470062 309454
rect 470146 309218 470382 309454
rect 469826 308898 470062 309134
rect 470146 308898 470382 309134
rect 478826 310158 479062 310394
rect 479146 310158 479382 310394
rect 478826 309838 479062 310074
rect 479146 309838 479382 310074
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 496826 310158 497062 310394
rect 497146 310158 497382 310394
rect 496826 309838 497062 310074
rect 497146 309838 497382 310074
rect 505826 309218 506062 309454
rect 506146 309218 506382 309454
rect 505826 308898 506062 309134
rect 506146 308898 506382 309134
rect 514826 310158 515062 310394
rect 515146 310158 515382 310394
rect 514826 309838 515062 310074
rect 515146 309838 515382 310074
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 532826 310158 533062 310394
rect 533146 310158 533382 310394
rect 532826 309838 533062 310074
rect 533146 309838 533382 310074
rect 541826 309218 542062 309454
rect 542146 309218 542382 309454
rect 541826 308898 542062 309134
rect 542146 308898 542382 309134
rect 550826 310158 551062 310394
rect 551146 310158 551382 310394
rect 550826 309838 551062 310074
rect 551146 309838 551382 310074
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 22916 300218 23152 300454
rect 22916 299898 23152 300134
rect 28847 300218 29083 300454
rect 28847 299898 29083 300134
rect 49916 300218 50152 300454
rect 49916 299898 50152 300134
rect 55847 300218 56083 300454
rect 55847 299898 56083 300134
rect 76916 300218 77152 300454
rect 76916 299898 77152 300134
rect 82847 300218 83083 300454
rect 82847 299898 83083 300134
rect 103916 300218 104152 300454
rect 103916 299898 104152 300134
rect 109847 300218 110083 300454
rect 109847 299898 110083 300134
rect 130916 300218 131152 300454
rect 130916 299898 131152 300134
rect 136847 300218 137083 300454
rect 136847 299898 137083 300134
rect 157916 300218 158152 300454
rect 157916 299898 158152 300134
rect 163847 300218 164083 300454
rect 163847 299898 164083 300134
rect 184916 300218 185152 300454
rect 184916 299898 185152 300134
rect 190847 300218 191083 300454
rect 190847 299898 191083 300134
rect 211916 300218 212152 300454
rect 211916 299898 212152 300134
rect 217847 300218 218083 300454
rect 217847 299898 218083 300134
rect 238916 300218 239152 300454
rect 238916 299898 239152 300134
rect 244847 300218 245083 300454
rect 244847 299898 245083 300134
rect 265916 300218 266152 300454
rect 265916 299898 266152 300134
rect 271847 300218 272083 300454
rect 271847 299898 272083 300134
rect 292916 300218 293152 300454
rect 292916 299898 293152 300134
rect 298847 300218 299083 300454
rect 298847 299898 299083 300134
rect 319916 300218 320152 300454
rect 319916 299898 320152 300134
rect 325847 300218 326083 300454
rect 325847 299898 326083 300134
rect 346916 300218 347152 300454
rect 346916 299898 347152 300134
rect 352847 300218 353083 300454
rect 352847 299898 353083 300134
rect 373916 300218 374152 300454
rect 373916 299898 374152 300134
rect 379847 300218 380083 300454
rect 379847 299898 380083 300134
rect 400916 300218 401152 300454
rect 400916 299898 401152 300134
rect 406847 300218 407083 300454
rect 406847 299898 407083 300134
rect 427916 300218 428152 300454
rect 427916 299898 428152 300134
rect 433847 300218 434083 300454
rect 433847 299898 434083 300134
rect 454916 300218 455152 300454
rect 454916 299898 455152 300134
rect 460847 300218 461083 300454
rect 460847 299898 461083 300134
rect 481916 300218 482152 300454
rect 481916 299898 482152 300134
rect 487847 300218 488083 300454
rect 487847 299898 488083 300134
rect 508916 300218 509152 300454
rect 508916 299898 509152 300134
rect 514847 300218 515083 300454
rect 514847 299898 515083 300134
rect 535916 300218 536152 300454
rect 535916 299898 536152 300134
rect 541847 300218 542083 300454
rect 541847 299898 542083 300134
rect 19952 291218 20188 291454
rect 19952 290898 20188 291134
rect 25882 291218 26118 291454
rect 25882 290898 26118 291134
rect 31813 291218 32049 291454
rect 31813 290898 32049 291134
rect 46952 291218 47188 291454
rect 46952 290898 47188 291134
rect 52882 291218 53118 291454
rect 52882 290898 53118 291134
rect 58813 291218 59049 291454
rect 58813 290898 59049 291134
rect 73952 291218 74188 291454
rect 73952 290898 74188 291134
rect 79882 291218 80118 291454
rect 79882 290898 80118 291134
rect 85813 291218 86049 291454
rect 85813 290898 86049 291134
rect 100952 291218 101188 291454
rect 100952 290898 101188 291134
rect 106882 291218 107118 291454
rect 106882 290898 107118 291134
rect 112813 291218 113049 291454
rect 112813 290898 113049 291134
rect 127952 291218 128188 291454
rect 127952 290898 128188 291134
rect 133882 291218 134118 291454
rect 133882 290898 134118 291134
rect 139813 291218 140049 291454
rect 139813 290898 140049 291134
rect 154952 291218 155188 291454
rect 154952 290898 155188 291134
rect 160882 291218 161118 291454
rect 160882 290898 161118 291134
rect 166813 291218 167049 291454
rect 166813 290898 167049 291134
rect 181952 291218 182188 291454
rect 181952 290898 182188 291134
rect 187882 291218 188118 291454
rect 187882 290898 188118 291134
rect 193813 291218 194049 291454
rect 193813 290898 194049 291134
rect 208952 291218 209188 291454
rect 208952 290898 209188 291134
rect 214882 291218 215118 291454
rect 214882 290898 215118 291134
rect 220813 291218 221049 291454
rect 220813 290898 221049 291134
rect 235952 291218 236188 291454
rect 235952 290898 236188 291134
rect 241882 291218 242118 291454
rect 241882 290898 242118 291134
rect 247813 291218 248049 291454
rect 247813 290898 248049 291134
rect 262952 291218 263188 291454
rect 262952 290898 263188 291134
rect 268882 291218 269118 291454
rect 268882 290898 269118 291134
rect 274813 291218 275049 291454
rect 274813 290898 275049 291134
rect 289952 291218 290188 291454
rect 289952 290898 290188 291134
rect 295882 291218 296118 291454
rect 295882 290898 296118 291134
rect 301813 291218 302049 291454
rect 301813 290898 302049 291134
rect 316952 291218 317188 291454
rect 316952 290898 317188 291134
rect 322882 291218 323118 291454
rect 322882 290898 323118 291134
rect 328813 291218 329049 291454
rect 328813 290898 329049 291134
rect 343952 291218 344188 291454
rect 343952 290898 344188 291134
rect 349882 291218 350118 291454
rect 349882 290898 350118 291134
rect 355813 291218 356049 291454
rect 355813 290898 356049 291134
rect 370952 291218 371188 291454
rect 370952 290898 371188 291134
rect 376882 291218 377118 291454
rect 376882 290898 377118 291134
rect 382813 291218 383049 291454
rect 382813 290898 383049 291134
rect 397952 291218 398188 291454
rect 397952 290898 398188 291134
rect 403882 291218 404118 291454
rect 403882 290898 404118 291134
rect 409813 291218 410049 291454
rect 409813 290898 410049 291134
rect 424952 291218 425188 291454
rect 424952 290898 425188 291134
rect 430882 291218 431118 291454
rect 430882 290898 431118 291134
rect 436813 291218 437049 291454
rect 436813 290898 437049 291134
rect 451952 291218 452188 291454
rect 451952 290898 452188 291134
rect 457882 291218 458118 291454
rect 457882 290898 458118 291134
rect 463813 291218 464049 291454
rect 463813 290898 464049 291134
rect 478952 291218 479188 291454
rect 478952 290898 479188 291134
rect 484882 291218 485118 291454
rect 484882 290898 485118 291134
rect 490813 291218 491049 291454
rect 490813 290898 491049 291134
rect 505952 291218 506188 291454
rect 505952 290898 506188 291134
rect 511882 291218 512118 291454
rect 511882 290898 512118 291134
rect 517813 291218 518049 291454
rect 517813 290898 518049 291134
rect 532952 291218 533188 291454
rect 532952 290898 533188 291134
rect 538882 291218 539118 291454
rect 538882 290898 539118 291134
rect 544813 291218 545049 291454
rect 544813 290898 545049 291134
rect 559826 291218 560062 291454
rect 560146 291218 560382 291454
rect 559826 290898 560062 291134
rect 560146 290898 560382 291134
rect 10826 282218 11062 282454
rect 11146 282218 11382 282454
rect 10826 281898 11062 282134
rect 11146 281898 11382 282134
rect 19826 283158 20062 283394
rect 20146 283158 20382 283394
rect 19826 282838 20062 283074
rect 20146 282838 20382 283074
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 37826 283158 38062 283394
rect 38146 283158 38382 283394
rect 37826 282838 38062 283074
rect 38146 282838 38382 283074
rect 46826 282218 47062 282454
rect 47146 282218 47382 282454
rect 46826 281898 47062 282134
rect 47146 281898 47382 282134
rect 55826 283158 56062 283394
rect 56146 283158 56382 283394
rect 55826 282838 56062 283074
rect 56146 282838 56382 283074
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 73826 283158 74062 283394
rect 74146 283158 74382 283394
rect 73826 282838 74062 283074
rect 74146 282838 74382 283074
rect 82826 282218 83062 282454
rect 83146 282218 83382 282454
rect 82826 281898 83062 282134
rect 83146 281898 83382 282134
rect 91826 283158 92062 283394
rect 92146 283158 92382 283394
rect 91826 282838 92062 283074
rect 92146 282838 92382 283074
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 109826 283158 110062 283394
rect 110146 283158 110382 283394
rect 109826 282838 110062 283074
rect 110146 282838 110382 283074
rect 118826 282218 119062 282454
rect 119146 282218 119382 282454
rect 118826 281898 119062 282134
rect 119146 281898 119382 282134
rect 127826 283158 128062 283394
rect 128146 283158 128382 283394
rect 127826 282838 128062 283074
rect 128146 282838 128382 283074
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 145826 283158 146062 283394
rect 146146 283158 146382 283394
rect 145826 282838 146062 283074
rect 146146 282838 146382 283074
rect 154826 282218 155062 282454
rect 155146 282218 155382 282454
rect 154826 281898 155062 282134
rect 155146 281898 155382 282134
rect 163826 283158 164062 283394
rect 164146 283158 164382 283394
rect 163826 282838 164062 283074
rect 164146 282838 164382 283074
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 181826 283158 182062 283394
rect 182146 283158 182382 283394
rect 181826 282838 182062 283074
rect 182146 282838 182382 283074
rect 190826 282218 191062 282454
rect 191146 282218 191382 282454
rect 190826 281898 191062 282134
rect 191146 281898 191382 282134
rect 199826 283158 200062 283394
rect 200146 283158 200382 283394
rect 199826 282838 200062 283074
rect 200146 282838 200382 283074
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 217826 283158 218062 283394
rect 218146 283158 218382 283394
rect 217826 282838 218062 283074
rect 218146 282838 218382 283074
rect 226826 282218 227062 282454
rect 227146 282218 227382 282454
rect 226826 281898 227062 282134
rect 227146 281898 227382 282134
rect 235826 283158 236062 283394
rect 236146 283158 236382 283394
rect 235826 282838 236062 283074
rect 236146 282838 236382 283074
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 253826 283158 254062 283394
rect 254146 283158 254382 283394
rect 253826 282838 254062 283074
rect 254146 282838 254382 283074
rect 262826 282218 263062 282454
rect 263146 282218 263382 282454
rect 262826 281898 263062 282134
rect 263146 281898 263382 282134
rect 271826 283158 272062 283394
rect 272146 283158 272382 283394
rect 271826 282838 272062 283074
rect 272146 282838 272382 283074
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 289826 283158 290062 283394
rect 290146 283158 290382 283394
rect 289826 282838 290062 283074
rect 290146 282838 290382 283074
rect 298826 282218 299062 282454
rect 299146 282218 299382 282454
rect 298826 281898 299062 282134
rect 299146 281898 299382 282134
rect 307826 283158 308062 283394
rect 308146 283158 308382 283394
rect 307826 282838 308062 283074
rect 308146 282838 308382 283074
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 325826 283158 326062 283394
rect 326146 283158 326382 283394
rect 325826 282838 326062 283074
rect 326146 282838 326382 283074
rect 334826 282218 335062 282454
rect 335146 282218 335382 282454
rect 334826 281898 335062 282134
rect 335146 281898 335382 282134
rect 343826 283158 344062 283394
rect 344146 283158 344382 283394
rect 343826 282838 344062 283074
rect 344146 282838 344382 283074
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 361826 283158 362062 283394
rect 362146 283158 362382 283394
rect 361826 282838 362062 283074
rect 362146 282838 362382 283074
rect 370826 282218 371062 282454
rect 371146 282218 371382 282454
rect 370826 281898 371062 282134
rect 371146 281898 371382 282134
rect 379826 283158 380062 283394
rect 380146 283158 380382 283394
rect 379826 282838 380062 283074
rect 380146 282838 380382 283074
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 397826 283158 398062 283394
rect 398146 283158 398382 283394
rect 397826 282838 398062 283074
rect 398146 282838 398382 283074
rect 406826 282218 407062 282454
rect 407146 282218 407382 282454
rect 406826 281898 407062 282134
rect 407146 281898 407382 282134
rect 415826 283158 416062 283394
rect 416146 283158 416382 283394
rect 415826 282838 416062 283074
rect 416146 282838 416382 283074
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 433826 283158 434062 283394
rect 434146 283158 434382 283394
rect 433826 282838 434062 283074
rect 434146 282838 434382 283074
rect 442826 282218 443062 282454
rect 443146 282218 443382 282454
rect 442826 281898 443062 282134
rect 443146 281898 443382 282134
rect 451826 283158 452062 283394
rect 452146 283158 452382 283394
rect 451826 282838 452062 283074
rect 452146 282838 452382 283074
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 469826 283158 470062 283394
rect 470146 283158 470382 283394
rect 469826 282838 470062 283074
rect 470146 282838 470382 283074
rect 478826 282218 479062 282454
rect 479146 282218 479382 282454
rect 478826 281898 479062 282134
rect 479146 281898 479382 282134
rect 487826 283158 488062 283394
rect 488146 283158 488382 283394
rect 487826 282838 488062 283074
rect 488146 282838 488382 283074
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 505826 283158 506062 283394
rect 506146 283158 506382 283394
rect 505826 282838 506062 283074
rect 506146 282838 506382 283074
rect 514826 282218 515062 282454
rect 515146 282218 515382 282454
rect 514826 281898 515062 282134
rect 515146 281898 515382 282134
rect 523826 283158 524062 283394
rect 524146 283158 524382 283394
rect 523826 282838 524062 283074
rect 524146 282838 524382 283074
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 541826 283158 542062 283394
rect 542146 283158 542382 283394
rect 541826 282838 542062 283074
rect 542146 282838 542382 283074
rect 550826 282218 551062 282454
rect 551146 282218 551382 282454
rect 550826 281898 551062 282134
rect 551146 281898 551382 282134
rect 19952 273218 20188 273454
rect 19952 272898 20188 273134
rect 25882 273218 26118 273454
rect 25882 272898 26118 273134
rect 31813 273218 32049 273454
rect 31813 272898 32049 273134
rect 46952 273218 47188 273454
rect 46952 272898 47188 273134
rect 52882 273218 53118 273454
rect 52882 272898 53118 273134
rect 58813 273218 59049 273454
rect 58813 272898 59049 273134
rect 73952 273218 74188 273454
rect 73952 272898 74188 273134
rect 79882 273218 80118 273454
rect 79882 272898 80118 273134
rect 85813 273218 86049 273454
rect 85813 272898 86049 273134
rect 100952 273218 101188 273454
rect 100952 272898 101188 273134
rect 106882 273218 107118 273454
rect 106882 272898 107118 273134
rect 112813 273218 113049 273454
rect 112813 272898 113049 273134
rect 127952 273218 128188 273454
rect 127952 272898 128188 273134
rect 133882 273218 134118 273454
rect 133882 272898 134118 273134
rect 139813 273218 140049 273454
rect 139813 272898 140049 273134
rect 154952 273218 155188 273454
rect 154952 272898 155188 273134
rect 160882 273218 161118 273454
rect 160882 272898 161118 273134
rect 166813 273218 167049 273454
rect 166813 272898 167049 273134
rect 181952 273218 182188 273454
rect 181952 272898 182188 273134
rect 187882 273218 188118 273454
rect 187882 272898 188118 273134
rect 193813 273218 194049 273454
rect 193813 272898 194049 273134
rect 208952 273218 209188 273454
rect 208952 272898 209188 273134
rect 214882 273218 215118 273454
rect 214882 272898 215118 273134
rect 220813 273218 221049 273454
rect 220813 272898 221049 273134
rect 235952 273218 236188 273454
rect 235952 272898 236188 273134
rect 241882 273218 242118 273454
rect 241882 272898 242118 273134
rect 247813 273218 248049 273454
rect 247813 272898 248049 273134
rect 262952 273218 263188 273454
rect 262952 272898 263188 273134
rect 268882 273218 269118 273454
rect 268882 272898 269118 273134
rect 274813 273218 275049 273454
rect 274813 272898 275049 273134
rect 289952 273218 290188 273454
rect 289952 272898 290188 273134
rect 295882 273218 296118 273454
rect 295882 272898 296118 273134
rect 301813 273218 302049 273454
rect 301813 272898 302049 273134
rect 316952 273218 317188 273454
rect 316952 272898 317188 273134
rect 322882 273218 323118 273454
rect 322882 272898 323118 273134
rect 328813 273218 329049 273454
rect 328813 272898 329049 273134
rect 343952 273218 344188 273454
rect 343952 272898 344188 273134
rect 349882 273218 350118 273454
rect 349882 272898 350118 273134
rect 355813 273218 356049 273454
rect 355813 272898 356049 273134
rect 370952 273218 371188 273454
rect 370952 272898 371188 273134
rect 376882 273218 377118 273454
rect 376882 272898 377118 273134
rect 382813 273218 383049 273454
rect 382813 272898 383049 273134
rect 397952 273218 398188 273454
rect 397952 272898 398188 273134
rect 403882 273218 404118 273454
rect 403882 272898 404118 273134
rect 409813 273218 410049 273454
rect 409813 272898 410049 273134
rect 424952 273218 425188 273454
rect 424952 272898 425188 273134
rect 430882 273218 431118 273454
rect 430882 272898 431118 273134
rect 436813 273218 437049 273454
rect 436813 272898 437049 273134
rect 451952 273218 452188 273454
rect 451952 272898 452188 273134
rect 457882 273218 458118 273454
rect 457882 272898 458118 273134
rect 463813 273218 464049 273454
rect 463813 272898 464049 273134
rect 478952 273218 479188 273454
rect 478952 272898 479188 273134
rect 484882 273218 485118 273454
rect 484882 272898 485118 273134
rect 490813 273218 491049 273454
rect 490813 272898 491049 273134
rect 505952 273218 506188 273454
rect 505952 272898 506188 273134
rect 511882 273218 512118 273454
rect 511882 272898 512118 273134
rect 517813 273218 518049 273454
rect 517813 272898 518049 273134
rect 532952 273218 533188 273454
rect 532952 272898 533188 273134
rect 538882 273218 539118 273454
rect 538882 272898 539118 273134
rect 544813 273218 545049 273454
rect 544813 272898 545049 273134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 22916 264218 23152 264454
rect 22916 263898 23152 264134
rect 28847 264218 29083 264454
rect 28847 263898 29083 264134
rect 49916 264218 50152 264454
rect 49916 263898 50152 264134
rect 55847 264218 56083 264454
rect 55847 263898 56083 264134
rect 76916 264218 77152 264454
rect 76916 263898 77152 264134
rect 82847 264218 83083 264454
rect 82847 263898 83083 264134
rect 103916 264218 104152 264454
rect 103916 263898 104152 264134
rect 109847 264218 110083 264454
rect 109847 263898 110083 264134
rect 130916 264218 131152 264454
rect 130916 263898 131152 264134
rect 136847 264218 137083 264454
rect 136847 263898 137083 264134
rect 157916 264218 158152 264454
rect 157916 263898 158152 264134
rect 163847 264218 164083 264454
rect 163847 263898 164083 264134
rect 184916 264218 185152 264454
rect 184916 263898 185152 264134
rect 190847 264218 191083 264454
rect 190847 263898 191083 264134
rect 211916 264218 212152 264454
rect 211916 263898 212152 264134
rect 217847 264218 218083 264454
rect 217847 263898 218083 264134
rect 238916 264218 239152 264454
rect 238916 263898 239152 264134
rect 244847 264218 245083 264454
rect 244847 263898 245083 264134
rect 265916 264218 266152 264454
rect 265916 263898 266152 264134
rect 271847 264218 272083 264454
rect 271847 263898 272083 264134
rect 292916 264218 293152 264454
rect 292916 263898 293152 264134
rect 298847 264218 299083 264454
rect 298847 263898 299083 264134
rect 319916 264218 320152 264454
rect 319916 263898 320152 264134
rect 325847 264218 326083 264454
rect 325847 263898 326083 264134
rect 346916 264218 347152 264454
rect 346916 263898 347152 264134
rect 352847 264218 353083 264454
rect 352847 263898 353083 264134
rect 373916 264218 374152 264454
rect 373916 263898 374152 264134
rect 379847 264218 380083 264454
rect 379847 263898 380083 264134
rect 400916 264218 401152 264454
rect 400916 263898 401152 264134
rect 406847 264218 407083 264454
rect 406847 263898 407083 264134
rect 427916 264218 428152 264454
rect 427916 263898 428152 264134
rect 433847 264218 434083 264454
rect 433847 263898 434083 264134
rect 454916 264218 455152 264454
rect 454916 263898 455152 264134
rect 460847 264218 461083 264454
rect 460847 263898 461083 264134
rect 481916 264218 482152 264454
rect 481916 263898 482152 264134
rect 487847 264218 488083 264454
rect 487847 263898 488083 264134
rect 508916 264218 509152 264454
rect 508916 263898 509152 264134
rect 514847 264218 515083 264454
rect 514847 263898 515083 264134
rect 535916 264218 536152 264454
rect 535916 263898 536152 264134
rect 541847 264218 542083 264454
rect 541847 263898 542083 264134
rect 19826 255218 20062 255454
rect 20146 255218 20382 255454
rect 19826 254898 20062 255134
rect 20146 254898 20382 255134
rect 28826 256158 29062 256394
rect 29146 256158 29382 256394
rect 28826 255838 29062 256074
rect 29146 255838 29382 256074
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 46826 256158 47062 256394
rect 47146 256158 47382 256394
rect 46826 255838 47062 256074
rect 47146 255838 47382 256074
rect 55826 255218 56062 255454
rect 56146 255218 56382 255454
rect 55826 254898 56062 255134
rect 56146 254898 56382 255134
rect 64826 256158 65062 256394
rect 65146 256158 65382 256394
rect 64826 255838 65062 256074
rect 65146 255838 65382 256074
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 82826 256158 83062 256394
rect 83146 256158 83382 256394
rect 82826 255838 83062 256074
rect 83146 255838 83382 256074
rect 91826 255218 92062 255454
rect 92146 255218 92382 255454
rect 91826 254898 92062 255134
rect 92146 254898 92382 255134
rect 100826 256158 101062 256394
rect 101146 256158 101382 256394
rect 100826 255838 101062 256074
rect 101146 255838 101382 256074
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 118826 256158 119062 256394
rect 119146 256158 119382 256394
rect 118826 255838 119062 256074
rect 119146 255838 119382 256074
rect 127826 255218 128062 255454
rect 128146 255218 128382 255454
rect 127826 254898 128062 255134
rect 128146 254898 128382 255134
rect 136826 256158 137062 256394
rect 137146 256158 137382 256394
rect 136826 255838 137062 256074
rect 137146 255838 137382 256074
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 154826 256158 155062 256394
rect 155146 256158 155382 256394
rect 154826 255838 155062 256074
rect 155146 255838 155382 256074
rect 163826 255218 164062 255454
rect 164146 255218 164382 255454
rect 163826 254898 164062 255134
rect 164146 254898 164382 255134
rect 172826 256158 173062 256394
rect 173146 256158 173382 256394
rect 172826 255838 173062 256074
rect 173146 255838 173382 256074
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 190826 256158 191062 256394
rect 191146 256158 191382 256394
rect 190826 255838 191062 256074
rect 191146 255838 191382 256074
rect 199826 255218 200062 255454
rect 200146 255218 200382 255454
rect 199826 254898 200062 255134
rect 200146 254898 200382 255134
rect 208826 256158 209062 256394
rect 209146 256158 209382 256394
rect 208826 255838 209062 256074
rect 209146 255838 209382 256074
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 226826 256158 227062 256394
rect 227146 256158 227382 256394
rect 226826 255838 227062 256074
rect 227146 255838 227382 256074
rect 235826 255218 236062 255454
rect 236146 255218 236382 255454
rect 235826 254898 236062 255134
rect 236146 254898 236382 255134
rect 244826 256158 245062 256394
rect 245146 256158 245382 256394
rect 244826 255838 245062 256074
rect 245146 255838 245382 256074
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 262826 256158 263062 256394
rect 263146 256158 263382 256394
rect 262826 255838 263062 256074
rect 263146 255838 263382 256074
rect 271826 255218 272062 255454
rect 272146 255218 272382 255454
rect 271826 254898 272062 255134
rect 272146 254898 272382 255134
rect 280826 256158 281062 256394
rect 281146 256158 281382 256394
rect 280826 255838 281062 256074
rect 281146 255838 281382 256074
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 298826 256158 299062 256394
rect 299146 256158 299382 256394
rect 298826 255838 299062 256074
rect 299146 255838 299382 256074
rect 307826 255218 308062 255454
rect 308146 255218 308382 255454
rect 307826 254898 308062 255134
rect 308146 254898 308382 255134
rect 316826 256158 317062 256394
rect 317146 256158 317382 256394
rect 316826 255838 317062 256074
rect 317146 255838 317382 256074
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 334826 256158 335062 256394
rect 335146 256158 335382 256394
rect 334826 255838 335062 256074
rect 335146 255838 335382 256074
rect 343826 255218 344062 255454
rect 344146 255218 344382 255454
rect 343826 254898 344062 255134
rect 344146 254898 344382 255134
rect 352826 256158 353062 256394
rect 353146 256158 353382 256394
rect 352826 255838 353062 256074
rect 353146 255838 353382 256074
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 370826 256158 371062 256394
rect 371146 256158 371382 256394
rect 370826 255838 371062 256074
rect 371146 255838 371382 256074
rect 379826 255218 380062 255454
rect 380146 255218 380382 255454
rect 379826 254898 380062 255134
rect 380146 254898 380382 255134
rect 388826 256158 389062 256394
rect 389146 256158 389382 256394
rect 388826 255838 389062 256074
rect 389146 255838 389382 256074
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 406826 256158 407062 256394
rect 407146 256158 407382 256394
rect 406826 255838 407062 256074
rect 407146 255838 407382 256074
rect 415826 255218 416062 255454
rect 416146 255218 416382 255454
rect 415826 254898 416062 255134
rect 416146 254898 416382 255134
rect 424826 256158 425062 256394
rect 425146 256158 425382 256394
rect 424826 255838 425062 256074
rect 425146 255838 425382 256074
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 442826 256158 443062 256394
rect 443146 256158 443382 256394
rect 442826 255838 443062 256074
rect 443146 255838 443382 256074
rect 451826 255218 452062 255454
rect 452146 255218 452382 255454
rect 451826 254898 452062 255134
rect 452146 254898 452382 255134
rect 460826 256158 461062 256394
rect 461146 256158 461382 256394
rect 460826 255838 461062 256074
rect 461146 255838 461382 256074
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 478826 256158 479062 256394
rect 479146 256158 479382 256394
rect 478826 255838 479062 256074
rect 479146 255838 479382 256074
rect 487826 255218 488062 255454
rect 488146 255218 488382 255454
rect 487826 254898 488062 255134
rect 488146 254898 488382 255134
rect 496826 256158 497062 256394
rect 497146 256158 497382 256394
rect 496826 255838 497062 256074
rect 497146 255838 497382 256074
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 514826 256158 515062 256394
rect 515146 256158 515382 256394
rect 514826 255838 515062 256074
rect 515146 255838 515382 256074
rect 523826 255218 524062 255454
rect 524146 255218 524382 255454
rect 523826 254898 524062 255134
rect 524146 254898 524382 255134
rect 532826 256158 533062 256394
rect 533146 256158 533382 256394
rect 532826 255838 533062 256074
rect 533146 255838 533382 256074
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 550826 256158 551062 256394
rect 551146 256158 551382 256394
rect 550826 255838 551062 256074
rect 551146 255838 551382 256074
rect 559826 255218 560062 255454
rect 560146 255218 560382 255454
rect 559826 254898 560062 255134
rect 560146 254898 560382 255134
rect 10826 246218 11062 246454
rect 11146 246218 11382 246454
rect 10826 245898 11062 246134
rect 11146 245898 11382 246134
rect 22916 246218 23152 246454
rect 22916 245898 23152 246134
rect 28847 246218 29083 246454
rect 28847 245898 29083 246134
rect 49916 246218 50152 246454
rect 49916 245898 50152 246134
rect 55847 246218 56083 246454
rect 55847 245898 56083 246134
rect 76916 246218 77152 246454
rect 76916 245898 77152 246134
rect 82847 246218 83083 246454
rect 82847 245898 83083 246134
rect 103916 246218 104152 246454
rect 103916 245898 104152 246134
rect 109847 246218 110083 246454
rect 109847 245898 110083 246134
rect 130916 246218 131152 246454
rect 130916 245898 131152 246134
rect 136847 246218 137083 246454
rect 136847 245898 137083 246134
rect 157916 246218 158152 246454
rect 157916 245898 158152 246134
rect 163847 246218 164083 246454
rect 163847 245898 164083 246134
rect 184916 246218 185152 246454
rect 184916 245898 185152 246134
rect 190847 246218 191083 246454
rect 190847 245898 191083 246134
rect 211916 246218 212152 246454
rect 211916 245898 212152 246134
rect 217847 246218 218083 246454
rect 217847 245898 218083 246134
rect 238916 246218 239152 246454
rect 238916 245898 239152 246134
rect 244847 246218 245083 246454
rect 244847 245898 245083 246134
rect 265916 246218 266152 246454
rect 265916 245898 266152 246134
rect 271847 246218 272083 246454
rect 271847 245898 272083 246134
rect 292916 246218 293152 246454
rect 292916 245898 293152 246134
rect 298847 246218 299083 246454
rect 298847 245898 299083 246134
rect 319916 246218 320152 246454
rect 319916 245898 320152 246134
rect 325847 246218 326083 246454
rect 325847 245898 326083 246134
rect 346916 246218 347152 246454
rect 346916 245898 347152 246134
rect 352847 246218 353083 246454
rect 352847 245898 353083 246134
rect 373916 246218 374152 246454
rect 373916 245898 374152 246134
rect 379847 246218 380083 246454
rect 379847 245898 380083 246134
rect 400916 246218 401152 246454
rect 400916 245898 401152 246134
rect 406847 246218 407083 246454
rect 406847 245898 407083 246134
rect 427916 246218 428152 246454
rect 427916 245898 428152 246134
rect 433847 246218 434083 246454
rect 433847 245898 434083 246134
rect 454916 246218 455152 246454
rect 454916 245898 455152 246134
rect 460847 246218 461083 246454
rect 460847 245898 461083 246134
rect 481916 246218 482152 246454
rect 481916 245898 482152 246134
rect 487847 246218 488083 246454
rect 487847 245898 488083 246134
rect 508916 246218 509152 246454
rect 508916 245898 509152 246134
rect 514847 246218 515083 246454
rect 514847 245898 515083 246134
rect 535916 246218 536152 246454
rect 535916 245898 536152 246134
rect 541847 246218 542083 246454
rect 541847 245898 542083 246134
rect 19952 237218 20188 237454
rect 19952 236898 20188 237134
rect 25882 237218 26118 237454
rect 25882 236898 26118 237134
rect 31813 237218 32049 237454
rect 31813 236898 32049 237134
rect 46952 237218 47188 237454
rect 46952 236898 47188 237134
rect 52882 237218 53118 237454
rect 52882 236898 53118 237134
rect 58813 237218 59049 237454
rect 58813 236898 59049 237134
rect 73952 237218 74188 237454
rect 73952 236898 74188 237134
rect 79882 237218 80118 237454
rect 79882 236898 80118 237134
rect 85813 237218 86049 237454
rect 85813 236898 86049 237134
rect 100952 237218 101188 237454
rect 100952 236898 101188 237134
rect 106882 237218 107118 237454
rect 106882 236898 107118 237134
rect 112813 237218 113049 237454
rect 112813 236898 113049 237134
rect 127952 237218 128188 237454
rect 127952 236898 128188 237134
rect 133882 237218 134118 237454
rect 133882 236898 134118 237134
rect 139813 237218 140049 237454
rect 139813 236898 140049 237134
rect 154952 237218 155188 237454
rect 154952 236898 155188 237134
rect 160882 237218 161118 237454
rect 160882 236898 161118 237134
rect 166813 237218 167049 237454
rect 166813 236898 167049 237134
rect 181952 237218 182188 237454
rect 181952 236898 182188 237134
rect 187882 237218 188118 237454
rect 187882 236898 188118 237134
rect 193813 237218 194049 237454
rect 193813 236898 194049 237134
rect 208952 237218 209188 237454
rect 208952 236898 209188 237134
rect 214882 237218 215118 237454
rect 214882 236898 215118 237134
rect 220813 237218 221049 237454
rect 220813 236898 221049 237134
rect 235952 237218 236188 237454
rect 235952 236898 236188 237134
rect 241882 237218 242118 237454
rect 241882 236898 242118 237134
rect 247813 237218 248049 237454
rect 247813 236898 248049 237134
rect 262952 237218 263188 237454
rect 262952 236898 263188 237134
rect 268882 237218 269118 237454
rect 268882 236898 269118 237134
rect 274813 237218 275049 237454
rect 274813 236898 275049 237134
rect 289952 237218 290188 237454
rect 289952 236898 290188 237134
rect 295882 237218 296118 237454
rect 295882 236898 296118 237134
rect 301813 237218 302049 237454
rect 301813 236898 302049 237134
rect 316952 237218 317188 237454
rect 316952 236898 317188 237134
rect 322882 237218 323118 237454
rect 322882 236898 323118 237134
rect 328813 237218 329049 237454
rect 328813 236898 329049 237134
rect 343952 237218 344188 237454
rect 343952 236898 344188 237134
rect 349882 237218 350118 237454
rect 349882 236898 350118 237134
rect 355813 237218 356049 237454
rect 355813 236898 356049 237134
rect 370952 237218 371188 237454
rect 370952 236898 371188 237134
rect 376882 237218 377118 237454
rect 376882 236898 377118 237134
rect 382813 237218 383049 237454
rect 382813 236898 383049 237134
rect 397952 237218 398188 237454
rect 397952 236898 398188 237134
rect 403882 237218 404118 237454
rect 403882 236898 404118 237134
rect 409813 237218 410049 237454
rect 409813 236898 410049 237134
rect 424952 237218 425188 237454
rect 424952 236898 425188 237134
rect 430882 237218 431118 237454
rect 430882 236898 431118 237134
rect 436813 237218 437049 237454
rect 436813 236898 437049 237134
rect 451952 237218 452188 237454
rect 451952 236898 452188 237134
rect 457882 237218 458118 237454
rect 457882 236898 458118 237134
rect 463813 237218 464049 237454
rect 463813 236898 464049 237134
rect 478952 237218 479188 237454
rect 478952 236898 479188 237134
rect 484882 237218 485118 237454
rect 484882 236898 485118 237134
rect 490813 237218 491049 237454
rect 490813 236898 491049 237134
rect 505952 237218 506188 237454
rect 505952 236898 506188 237134
rect 511882 237218 512118 237454
rect 511882 236898 512118 237134
rect 517813 237218 518049 237454
rect 517813 236898 518049 237134
rect 532952 237218 533188 237454
rect 532952 236898 533188 237134
rect 538882 237218 539118 237454
rect 538882 236898 539118 237134
rect 544813 237218 545049 237454
rect 544813 236898 545049 237134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 19826 229158 20062 229394
rect 20146 229158 20382 229394
rect 19826 228838 20062 229074
rect 20146 228838 20382 229074
rect 28826 228218 29062 228454
rect 29146 228218 29382 228454
rect 28826 227898 29062 228134
rect 29146 227898 29382 228134
rect 37826 229158 38062 229394
rect 38146 229158 38382 229394
rect 37826 228838 38062 229074
rect 38146 228838 38382 229074
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 55826 229158 56062 229394
rect 56146 229158 56382 229394
rect 55826 228838 56062 229074
rect 56146 228838 56382 229074
rect 64826 228218 65062 228454
rect 65146 228218 65382 228454
rect 64826 227898 65062 228134
rect 65146 227898 65382 228134
rect 73826 229158 74062 229394
rect 74146 229158 74382 229394
rect 73826 228838 74062 229074
rect 74146 228838 74382 229074
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 91826 229158 92062 229394
rect 92146 229158 92382 229394
rect 91826 228838 92062 229074
rect 92146 228838 92382 229074
rect 100826 228218 101062 228454
rect 101146 228218 101382 228454
rect 100826 227898 101062 228134
rect 101146 227898 101382 228134
rect 109826 229158 110062 229394
rect 110146 229158 110382 229394
rect 109826 228838 110062 229074
rect 110146 228838 110382 229074
rect 118826 228218 119062 228454
rect 119146 228218 119382 228454
rect 118826 227898 119062 228134
rect 119146 227898 119382 228134
rect 127826 229158 128062 229394
rect 128146 229158 128382 229394
rect 127826 228838 128062 229074
rect 128146 228838 128382 229074
rect 136826 228218 137062 228454
rect 137146 228218 137382 228454
rect 136826 227898 137062 228134
rect 137146 227898 137382 228134
rect 145826 229158 146062 229394
rect 146146 229158 146382 229394
rect 145826 228838 146062 229074
rect 146146 228838 146382 229074
rect 154826 228218 155062 228454
rect 155146 228218 155382 228454
rect 154826 227898 155062 228134
rect 155146 227898 155382 228134
rect 163826 229158 164062 229394
rect 164146 229158 164382 229394
rect 163826 228838 164062 229074
rect 164146 228838 164382 229074
rect 172826 228218 173062 228454
rect 173146 228218 173382 228454
rect 172826 227898 173062 228134
rect 173146 227898 173382 228134
rect 181826 229158 182062 229394
rect 182146 229158 182382 229394
rect 181826 228838 182062 229074
rect 182146 228838 182382 229074
rect 190826 228218 191062 228454
rect 191146 228218 191382 228454
rect 190826 227898 191062 228134
rect 191146 227898 191382 228134
rect 199826 229158 200062 229394
rect 200146 229158 200382 229394
rect 199826 228838 200062 229074
rect 200146 228838 200382 229074
rect 208826 228218 209062 228454
rect 209146 228218 209382 228454
rect 208826 227898 209062 228134
rect 209146 227898 209382 228134
rect 217826 229158 218062 229394
rect 218146 229158 218382 229394
rect 217826 228838 218062 229074
rect 218146 228838 218382 229074
rect 226826 228218 227062 228454
rect 227146 228218 227382 228454
rect 226826 227898 227062 228134
rect 227146 227898 227382 228134
rect 235826 229158 236062 229394
rect 236146 229158 236382 229394
rect 235826 228838 236062 229074
rect 236146 228838 236382 229074
rect 244826 228218 245062 228454
rect 245146 228218 245382 228454
rect 244826 227898 245062 228134
rect 245146 227898 245382 228134
rect 253826 229158 254062 229394
rect 254146 229158 254382 229394
rect 253826 228838 254062 229074
rect 254146 228838 254382 229074
rect 262826 228218 263062 228454
rect 263146 228218 263382 228454
rect 262826 227898 263062 228134
rect 263146 227898 263382 228134
rect 271826 229158 272062 229394
rect 272146 229158 272382 229394
rect 271826 228838 272062 229074
rect 272146 228838 272382 229074
rect 280826 228218 281062 228454
rect 281146 228218 281382 228454
rect 280826 227898 281062 228134
rect 281146 227898 281382 228134
rect 289826 229158 290062 229394
rect 290146 229158 290382 229394
rect 289826 228838 290062 229074
rect 290146 228838 290382 229074
rect 298826 228218 299062 228454
rect 299146 228218 299382 228454
rect 298826 227898 299062 228134
rect 299146 227898 299382 228134
rect 307826 229158 308062 229394
rect 308146 229158 308382 229394
rect 307826 228838 308062 229074
rect 308146 228838 308382 229074
rect 316826 228218 317062 228454
rect 317146 228218 317382 228454
rect 316826 227898 317062 228134
rect 317146 227898 317382 228134
rect 325826 229158 326062 229394
rect 326146 229158 326382 229394
rect 325826 228838 326062 229074
rect 326146 228838 326382 229074
rect 334826 228218 335062 228454
rect 335146 228218 335382 228454
rect 334826 227898 335062 228134
rect 335146 227898 335382 228134
rect 343826 229158 344062 229394
rect 344146 229158 344382 229394
rect 343826 228838 344062 229074
rect 344146 228838 344382 229074
rect 352826 228218 353062 228454
rect 353146 228218 353382 228454
rect 352826 227898 353062 228134
rect 353146 227898 353382 228134
rect 361826 229158 362062 229394
rect 362146 229158 362382 229394
rect 361826 228838 362062 229074
rect 362146 228838 362382 229074
rect 370826 228218 371062 228454
rect 371146 228218 371382 228454
rect 370826 227898 371062 228134
rect 371146 227898 371382 228134
rect 379826 229158 380062 229394
rect 380146 229158 380382 229394
rect 379826 228838 380062 229074
rect 380146 228838 380382 229074
rect 388826 228218 389062 228454
rect 389146 228218 389382 228454
rect 388826 227898 389062 228134
rect 389146 227898 389382 228134
rect 397826 229158 398062 229394
rect 398146 229158 398382 229394
rect 397826 228838 398062 229074
rect 398146 228838 398382 229074
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 415826 229158 416062 229394
rect 416146 229158 416382 229394
rect 415826 228838 416062 229074
rect 416146 228838 416382 229074
rect 424826 228218 425062 228454
rect 425146 228218 425382 228454
rect 424826 227898 425062 228134
rect 425146 227898 425382 228134
rect 433826 229158 434062 229394
rect 434146 229158 434382 229394
rect 433826 228838 434062 229074
rect 434146 228838 434382 229074
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 451826 229158 452062 229394
rect 452146 229158 452382 229394
rect 451826 228838 452062 229074
rect 452146 228838 452382 229074
rect 460826 228218 461062 228454
rect 461146 228218 461382 228454
rect 460826 227898 461062 228134
rect 461146 227898 461382 228134
rect 469826 229158 470062 229394
rect 470146 229158 470382 229394
rect 469826 228838 470062 229074
rect 470146 228838 470382 229074
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 487826 229158 488062 229394
rect 488146 229158 488382 229394
rect 487826 228838 488062 229074
rect 488146 228838 488382 229074
rect 496826 228218 497062 228454
rect 497146 228218 497382 228454
rect 496826 227898 497062 228134
rect 497146 227898 497382 228134
rect 505826 229158 506062 229394
rect 506146 229158 506382 229394
rect 505826 228838 506062 229074
rect 506146 228838 506382 229074
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 523826 229158 524062 229394
rect 524146 229158 524382 229394
rect 523826 228838 524062 229074
rect 524146 228838 524382 229074
rect 532826 228218 533062 228454
rect 533146 228218 533382 228454
rect 532826 227898 533062 228134
rect 533146 227898 533382 228134
rect 541826 229158 542062 229394
rect 542146 229158 542382 229394
rect 541826 228838 542062 229074
rect 542146 228838 542382 229074
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 19952 219218 20188 219454
rect 19952 218898 20188 219134
rect 25882 219218 26118 219454
rect 25882 218898 26118 219134
rect 31813 219218 32049 219454
rect 31813 218898 32049 219134
rect 46952 219218 47188 219454
rect 46952 218898 47188 219134
rect 52882 219218 53118 219454
rect 52882 218898 53118 219134
rect 58813 219218 59049 219454
rect 58813 218898 59049 219134
rect 73952 219218 74188 219454
rect 73952 218898 74188 219134
rect 79882 219218 80118 219454
rect 79882 218898 80118 219134
rect 85813 219218 86049 219454
rect 85813 218898 86049 219134
rect 100952 219218 101188 219454
rect 100952 218898 101188 219134
rect 106882 219218 107118 219454
rect 106882 218898 107118 219134
rect 112813 219218 113049 219454
rect 112813 218898 113049 219134
rect 127952 219218 128188 219454
rect 127952 218898 128188 219134
rect 133882 219218 134118 219454
rect 133882 218898 134118 219134
rect 139813 219218 140049 219454
rect 139813 218898 140049 219134
rect 154952 219218 155188 219454
rect 154952 218898 155188 219134
rect 160882 219218 161118 219454
rect 160882 218898 161118 219134
rect 166813 219218 167049 219454
rect 166813 218898 167049 219134
rect 181952 219218 182188 219454
rect 181952 218898 182188 219134
rect 187882 219218 188118 219454
rect 187882 218898 188118 219134
rect 193813 219218 194049 219454
rect 193813 218898 194049 219134
rect 208952 219218 209188 219454
rect 208952 218898 209188 219134
rect 214882 219218 215118 219454
rect 214882 218898 215118 219134
rect 220813 219218 221049 219454
rect 220813 218898 221049 219134
rect 235952 219218 236188 219454
rect 235952 218898 236188 219134
rect 241882 219218 242118 219454
rect 241882 218898 242118 219134
rect 247813 219218 248049 219454
rect 247813 218898 248049 219134
rect 262952 219218 263188 219454
rect 262952 218898 263188 219134
rect 268882 219218 269118 219454
rect 268882 218898 269118 219134
rect 274813 219218 275049 219454
rect 274813 218898 275049 219134
rect 289952 219218 290188 219454
rect 289952 218898 290188 219134
rect 295882 219218 296118 219454
rect 295882 218898 296118 219134
rect 301813 219218 302049 219454
rect 301813 218898 302049 219134
rect 316952 219218 317188 219454
rect 316952 218898 317188 219134
rect 322882 219218 323118 219454
rect 322882 218898 323118 219134
rect 328813 219218 329049 219454
rect 328813 218898 329049 219134
rect 343952 219218 344188 219454
rect 343952 218898 344188 219134
rect 349882 219218 350118 219454
rect 349882 218898 350118 219134
rect 355813 219218 356049 219454
rect 355813 218898 356049 219134
rect 370952 219218 371188 219454
rect 370952 218898 371188 219134
rect 376882 219218 377118 219454
rect 376882 218898 377118 219134
rect 382813 219218 383049 219454
rect 382813 218898 383049 219134
rect 397952 219218 398188 219454
rect 397952 218898 398188 219134
rect 403882 219218 404118 219454
rect 403882 218898 404118 219134
rect 409813 219218 410049 219454
rect 409813 218898 410049 219134
rect 424952 219218 425188 219454
rect 424952 218898 425188 219134
rect 430882 219218 431118 219454
rect 430882 218898 431118 219134
rect 436813 219218 437049 219454
rect 436813 218898 437049 219134
rect 451952 219218 452188 219454
rect 451952 218898 452188 219134
rect 457882 219218 458118 219454
rect 457882 218898 458118 219134
rect 463813 219218 464049 219454
rect 463813 218898 464049 219134
rect 478952 219218 479188 219454
rect 478952 218898 479188 219134
rect 484882 219218 485118 219454
rect 484882 218898 485118 219134
rect 490813 219218 491049 219454
rect 490813 218898 491049 219134
rect 505952 219218 506188 219454
rect 505952 218898 506188 219134
rect 511882 219218 512118 219454
rect 511882 218898 512118 219134
rect 517813 219218 518049 219454
rect 517813 218898 518049 219134
rect 532952 219218 533188 219454
rect 532952 218898 533188 219134
rect 538882 219218 539118 219454
rect 538882 218898 539118 219134
rect 544813 219218 545049 219454
rect 544813 218898 545049 219134
rect 559826 219218 560062 219454
rect 560146 219218 560382 219454
rect 559826 218898 560062 219134
rect 560146 218898 560382 219134
rect 10826 210218 11062 210454
rect 11146 210218 11382 210454
rect 10826 209898 11062 210134
rect 11146 209898 11382 210134
rect 22916 210218 23152 210454
rect 22916 209898 23152 210134
rect 28847 210218 29083 210454
rect 28847 209898 29083 210134
rect 49916 210218 50152 210454
rect 49916 209898 50152 210134
rect 55847 210218 56083 210454
rect 55847 209898 56083 210134
rect 76916 210218 77152 210454
rect 76916 209898 77152 210134
rect 82847 210218 83083 210454
rect 82847 209898 83083 210134
rect 103916 210218 104152 210454
rect 103916 209898 104152 210134
rect 109847 210218 110083 210454
rect 109847 209898 110083 210134
rect 130916 210218 131152 210454
rect 130916 209898 131152 210134
rect 136847 210218 137083 210454
rect 136847 209898 137083 210134
rect 157916 210218 158152 210454
rect 157916 209898 158152 210134
rect 163847 210218 164083 210454
rect 163847 209898 164083 210134
rect 184916 210218 185152 210454
rect 184916 209898 185152 210134
rect 190847 210218 191083 210454
rect 190847 209898 191083 210134
rect 211916 210218 212152 210454
rect 211916 209898 212152 210134
rect 217847 210218 218083 210454
rect 217847 209898 218083 210134
rect 238916 210218 239152 210454
rect 238916 209898 239152 210134
rect 244847 210218 245083 210454
rect 244847 209898 245083 210134
rect 265916 210218 266152 210454
rect 265916 209898 266152 210134
rect 271847 210218 272083 210454
rect 271847 209898 272083 210134
rect 292916 210218 293152 210454
rect 292916 209898 293152 210134
rect 298847 210218 299083 210454
rect 298847 209898 299083 210134
rect 319916 210218 320152 210454
rect 319916 209898 320152 210134
rect 325847 210218 326083 210454
rect 325847 209898 326083 210134
rect 346916 210218 347152 210454
rect 346916 209898 347152 210134
rect 352847 210218 353083 210454
rect 352847 209898 353083 210134
rect 373916 210218 374152 210454
rect 373916 209898 374152 210134
rect 379847 210218 380083 210454
rect 379847 209898 380083 210134
rect 400916 210218 401152 210454
rect 400916 209898 401152 210134
rect 406847 210218 407083 210454
rect 406847 209898 407083 210134
rect 427916 210218 428152 210454
rect 427916 209898 428152 210134
rect 433847 210218 434083 210454
rect 433847 209898 434083 210134
rect 454916 210218 455152 210454
rect 454916 209898 455152 210134
rect 460847 210218 461083 210454
rect 460847 209898 461083 210134
rect 481916 210218 482152 210454
rect 481916 209898 482152 210134
rect 487847 210218 488083 210454
rect 487847 209898 488083 210134
rect 508916 210218 509152 210454
rect 508916 209898 509152 210134
rect 514847 210218 515083 210454
rect 514847 209898 515083 210134
rect 535916 210218 536152 210454
rect 535916 209898 536152 210134
rect 541847 210218 542083 210454
rect 541847 209898 542083 210134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 28826 202158 29062 202394
rect 29146 202158 29382 202394
rect 28826 201838 29062 202074
rect 29146 201838 29382 202074
rect 37826 201218 38062 201454
rect 38146 201218 38382 201454
rect 37826 200898 38062 201134
rect 38146 200898 38382 201134
rect 46826 202158 47062 202394
rect 47146 202158 47382 202394
rect 46826 201838 47062 202074
rect 47146 201838 47382 202074
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 64826 202158 65062 202394
rect 65146 202158 65382 202394
rect 64826 201838 65062 202074
rect 65146 201838 65382 202074
rect 73826 201218 74062 201454
rect 74146 201218 74382 201454
rect 73826 200898 74062 201134
rect 74146 200898 74382 201134
rect 82826 202158 83062 202394
rect 83146 202158 83382 202394
rect 82826 201838 83062 202074
rect 83146 201838 83382 202074
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 100826 202158 101062 202394
rect 101146 202158 101382 202394
rect 100826 201838 101062 202074
rect 101146 201838 101382 202074
rect 109826 201218 110062 201454
rect 110146 201218 110382 201454
rect 109826 200898 110062 201134
rect 110146 200898 110382 201134
rect 118826 202158 119062 202394
rect 119146 202158 119382 202394
rect 118826 201838 119062 202074
rect 119146 201838 119382 202074
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 136826 202158 137062 202394
rect 137146 202158 137382 202394
rect 136826 201838 137062 202074
rect 137146 201838 137382 202074
rect 145826 201218 146062 201454
rect 146146 201218 146382 201454
rect 145826 200898 146062 201134
rect 146146 200898 146382 201134
rect 154826 202158 155062 202394
rect 155146 202158 155382 202394
rect 154826 201838 155062 202074
rect 155146 201838 155382 202074
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 172826 202158 173062 202394
rect 173146 202158 173382 202394
rect 172826 201838 173062 202074
rect 173146 201838 173382 202074
rect 181826 201218 182062 201454
rect 182146 201218 182382 201454
rect 181826 200898 182062 201134
rect 182146 200898 182382 201134
rect 190826 202158 191062 202394
rect 191146 202158 191382 202394
rect 190826 201838 191062 202074
rect 191146 201838 191382 202074
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 208826 202158 209062 202394
rect 209146 202158 209382 202394
rect 208826 201838 209062 202074
rect 209146 201838 209382 202074
rect 217826 201218 218062 201454
rect 218146 201218 218382 201454
rect 217826 200898 218062 201134
rect 218146 200898 218382 201134
rect 226826 202158 227062 202394
rect 227146 202158 227382 202394
rect 226826 201838 227062 202074
rect 227146 201838 227382 202074
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 244826 202158 245062 202394
rect 245146 202158 245382 202394
rect 244826 201838 245062 202074
rect 245146 201838 245382 202074
rect 253826 201218 254062 201454
rect 254146 201218 254382 201454
rect 253826 200898 254062 201134
rect 254146 200898 254382 201134
rect 262826 202158 263062 202394
rect 263146 202158 263382 202394
rect 262826 201838 263062 202074
rect 263146 201838 263382 202074
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 280826 202158 281062 202394
rect 281146 202158 281382 202394
rect 280826 201838 281062 202074
rect 281146 201838 281382 202074
rect 289826 201218 290062 201454
rect 290146 201218 290382 201454
rect 289826 200898 290062 201134
rect 290146 200898 290382 201134
rect 298826 202158 299062 202394
rect 299146 202158 299382 202394
rect 298826 201838 299062 202074
rect 299146 201838 299382 202074
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 316826 202158 317062 202394
rect 317146 202158 317382 202394
rect 316826 201838 317062 202074
rect 317146 201838 317382 202074
rect 325826 201218 326062 201454
rect 326146 201218 326382 201454
rect 325826 200898 326062 201134
rect 326146 200898 326382 201134
rect 334826 202158 335062 202394
rect 335146 202158 335382 202394
rect 334826 201838 335062 202074
rect 335146 201838 335382 202074
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 352826 202158 353062 202394
rect 353146 202158 353382 202394
rect 352826 201838 353062 202074
rect 353146 201838 353382 202074
rect 361826 201218 362062 201454
rect 362146 201218 362382 201454
rect 361826 200898 362062 201134
rect 362146 200898 362382 201134
rect 370826 202158 371062 202394
rect 371146 202158 371382 202394
rect 370826 201838 371062 202074
rect 371146 201838 371382 202074
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 388826 202158 389062 202394
rect 389146 202158 389382 202394
rect 388826 201838 389062 202074
rect 389146 201838 389382 202074
rect 397826 201218 398062 201454
rect 398146 201218 398382 201454
rect 397826 200898 398062 201134
rect 398146 200898 398382 201134
rect 406826 202158 407062 202394
rect 407146 202158 407382 202394
rect 406826 201838 407062 202074
rect 407146 201838 407382 202074
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 424826 202158 425062 202394
rect 425146 202158 425382 202394
rect 424826 201838 425062 202074
rect 425146 201838 425382 202074
rect 433826 201218 434062 201454
rect 434146 201218 434382 201454
rect 433826 200898 434062 201134
rect 434146 200898 434382 201134
rect 442826 202158 443062 202394
rect 443146 202158 443382 202394
rect 442826 201838 443062 202074
rect 443146 201838 443382 202074
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 460826 202158 461062 202394
rect 461146 202158 461382 202394
rect 460826 201838 461062 202074
rect 461146 201838 461382 202074
rect 469826 201218 470062 201454
rect 470146 201218 470382 201454
rect 469826 200898 470062 201134
rect 470146 200898 470382 201134
rect 478826 202158 479062 202394
rect 479146 202158 479382 202394
rect 478826 201838 479062 202074
rect 479146 201838 479382 202074
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 496826 202158 497062 202394
rect 497146 202158 497382 202394
rect 496826 201838 497062 202074
rect 497146 201838 497382 202074
rect 505826 201218 506062 201454
rect 506146 201218 506382 201454
rect 505826 200898 506062 201134
rect 506146 200898 506382 201134
rect 514826 202158 515062 202394
rect 515146 202158 515382 202394
rect 514826 201838 515062 202074
rect 515146 201838 515382 202074
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 532826 202158 533062 202394
rect 533146 202158 533382 202394
rect 532826 201838 533062 202074
rect 533146 201838 533382 202074
rect 541826 201218 542062 201454
rect 542146 201218 542382 201454
rect 541826 200898 542062 201134
rect 542146 200898 542382 201134
rect 550826 202158 551062 202394
rect 551146 202158 551382 202394
rect 550826 201838 551062 202074
rect 551146 201838 551382 202074
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 22916 192218 23152 192454
rect 22916 191898 23152 192134
rect 28847 192218 29083 192454
rect 28847 191898 29083 192134
rect 49916 192218 50152 192454
rect 49916 191898 50152 192134
rect 55847 192218 56083 192454
rect 55847 191898 56083 192134
rect 76916 192218 77152 192454
rect 76916 191898 77152 192134
rect 82847 192218 83083 192454
rect 82847 191898 83083 192134
rect 103916 192218 104152 192454
rect 103916 191898 104152 192134
rect 109847 192218 110083 192454
rect 109847 191898 110083 192134
rect 130916 192218 131152 192454
rect 130916 191898 131152 192134
rect 136847 192218 137083 192454
rect 136847 191898 137083 192134
rect 157916 192218 158152 192454
rect 157916 191898 158152 192134
rect 163847 192218 164083 192454
rect 163847 191898 164083 192134
rect 184916 192218 185152 192454
rect 184916 191898 185152 192134
rect 190847 192218 191083 192454
rect 190847 191898 191083 192134
rect 211916 192218 212152 192454
rect 211916 191898 212152 192134
rect 217847 192218 218083 192454
rect 217847 191898 218083 192134
rect 238916 192218 239152 192454
rect 238916 191898 239152 192134
rect 244847 192218 245083 192454
rect 244847 191898 245083 192134
rect 265916 192218 266152 192454
rect 265916 191898 266152 192134
rect 271847 192218 272083 192454
rect 271847 191898 272083 192134
rect 292916 192218 293152 192454
rect 292916 191898 293152 192134
rect 298847 192218 299083 192454
rect 298847 191898 299083 192134
rect 319916 192218 320152 192454
rect 319916 191898 320152 192134
rect 325847 192218 326083 192454
rect 325847 191898 326083 192134
rect 346916 192218 347152 192454
rect 346916 191898 347152 192134
rect 352847 192218 353083 192454
rect 352847 191898 353083 192134
rect 373916 192218 374152 192454
rect 373916 191898 374152 192134
rect 379847 192218 380083 192454
rect 379847 191898 380083 192134
rect 400916 192218 401152 192454
rect 400916 191898 401152 192134
rect 406847 192218 407083 192454
rect 406847 191898 407083 192134
rect 427916 192218 428152 192454
rect 427916 191898 428152 192134
rect 433847 192218 434083 192454
rect 433847 191898 434083 192134
rect 454916 192218 455152 192454
rect 454916 191898 455152 192134
rect 460847 192218 461083 192454
rect 460847 191898 461083 192134
rect 481916 192218 482152 192454
rect 481916 191898 482152 192134
rect 487847 192218 488083 192454
rect 487847 191898 488083 192134
rect 508916 192218 509152 192454
rect 508916 191898 509152 192134
rect 514847 192218 515083 192454
rect 514847 191898 515083 192134
rect 535916 192218 536152 192454
rect 535916 191898 536152 192134
rect 541847 192218 542083 192454
rect 541847 191898 542083 192134
rect 19952 183218 20188 183454
rect 19952 182898 20188 183134
rect 25882 183218 26118 183454
rect 25882 182898 26118 183134
rect 31813 183218 32049 183454
rect 31813 182898 32049 183134
rect 46952 183218 47188 183454
rect 46952 182898 47188 183134
rect 52882 183218 53118 183454
rect 52882 182898 53118 183134
rect 58813 183218 59049 183454
rect 58813 182898 59049 183134
rect 73952 183218 74188 183454
rect 73952 182898 74188 183134
rect 79882 183218 80118 183454
rect 79882 182898 80118 183134
rect 85813 183218 86049 183454
rect 85813 182898 86049 183134
rect 100952 183218 101188 183454
rect 100952 182898 101188 183134
rect 106882 183218 107118 183454
rect 106882 182898 107118 183134
rect 112813 183218 113049 183454
rect 112813 182898 113049 183134
rect 127952 183218 128188 183454
rect 127952 182898 128188 183134
rect 133882 183218 134118 183454
rect 133882 182898 134118 183134
rect 139813 183218 140049 183454
rect 139813 182898 140049 183134
rect 154952 183218 155188 183454
rect 154952 182898 155188 183134
rect 160882 183218 161118 183454
rect 160882 182898 161118 183134
rect 166813 183218 167049 183454
rect 166813 182898 167049 183134
rect 181952 183218 182188 183454
rect 181952 182898 182188 183134
rect 187882 183218 188118 183454
rect 187882 182898 188118 183134
rect 193813 183218 194049 183454
rect 193813 182898 194049 183134
rect 208952 183218 209188 183454
rect 208952 182898 209188 183134
rect 214882 183218 215118 183454
rect 214882 182898 215118 183134
rect 220813 183218 221049 183454
rect 220813 182898 221049 183134
rect 235952 183218 236188 183454
rect 235952 182898 236188 183134
rect 241882 183218 242118 183454
rect 241882 182898 242118 183134
rect 247813 183218 248049 183454
rect 247813 182898 248049 183134
rect 262952 183218 263188 183454
rect 262952 182898 263188 183134
rect 268882 183218 269118 183454
rect 268882 182898 269118 183134
rect 274813 183218 275049 183454
rect 274813 182898 275049 183134
rect 289952 183218 290188 183454
rect 289952 182898 290188 183134
rect 295882 183218 296118 183454
rect 295882 182898 296118 183134
rect 301813 183218 302049 183454
rect 301813 182898 302049 183134
rect 316952 183218 317188 183454
rect 316952 182898 317188 183134
rect 322882 183218 323118 183454
rect 322882 182898 323118 183134
rect 328813 183218 329049 183454
rect 328813 182898 329049 183134
rect 343952 183218 344188 183454
rect 343952 182898 344188 183134
rect 349882 183218 350118 183454
rect 349882 182898 350118 183134
rect 355813 183218 356049 183454
rect 355813 182898 356049 183134
rect 370952 183218 371188 183454
rect 370952 182898 371188 183134
rect 376882 183218 377118 183454
rect 376882 182898 377118 183134
rect 382813 183218 383049 183454
rect 382813 182898 383049 183134
rect 397952 183218 398188 183454
rect 397952 182898 398188 183134
rect 403882 183218 404118 183454
rect 403882 182898 404118 183134
rect 409813 183218 410049 183454
rect 409813 182898 410049 183134
rect 424952 183218 425188 183454
rect 424952 182898 425188 183134
rect 430882 183218 431118 183454
rect 430882 182898 431118 183134
rect 436813 183218 437049 183454
rect 436813 182898 437049 183134
rect 451952 183218 452188 183454
rect 451952 182898 452188 183134
rect 457882 183218 458118 183454
rect 457882 182898 458118 183134
rect 463813 183218 464049 183454
rect 463813 182898 464049 183134
rect 478952 183218 479188 183454
rect 478952 182898 479188 183134
rect 484882 183218 485118 183454
rect 484882 182898 485118 183134
rect 490813 183218 491049 183454
rect 490813 182898 491049 183134
rect 505952 183218 506188 183454
rect 505952 182898 506188 183134
rect 511882 183218 512118 183454
rect 511882 182898 512118 183134
rect 517813 183218 518049 183454
rect 517813 182898 518049 183134
rect 532952 183218 533188 183454
rect 532952 182898 533188 183134
rect 538882 183218 539118 183454
rect 538882 182898 539118 183134
rect 544813 183218 545049 183454
rect 544813 182898 545049 183134
rect 559826 183218 560062 183454
rect 560146 183218 560382 183454
rect 559826 182898 560062 183134
rect 560146 182898 560382 183134
rect 10826 174218 11062 174454
rect 11146 174218 11382 174454
rect 10826 173898 11062 174134
rect 11146 173898 11382 174134
rect 19826 175158 20062 175394
rect 20146 175158 20382 175394
rect 19826 174838 20062 175074
rect 20146 174838 20382 175074
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 37826 175158 38062 175394
rect 38146 175158 38382 175394
rect 37826 174838 38062 175074
rect 38146 174838 38382 175074
rect 46826 174218 47062 174454
rect 47146 174218 47382 174454
rect 46826 173898 47062 174134
rect 47146 173898 47382 174134
rect 55826 175158 56062 175394
rect 56146 175158 56382 175394
rect 55826 174838 56062 175074
rect 56146 174838 56382 175074
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 73826 175158 74062 175394
rect 74146 175158 74382 175394
rect 73826 174838 74062 175074
rect 74146 174838 74382 175074
rect 82826 174218 83062 174454
rect 83146 174218 83382 174454
rect 82826 173898 83062 174134
rect 83146 173898 83382 174134
rect 91826 175158 92062 175394
rect 92146 175158 92382 175394
rect 91826 174838 92062 175074
rect 92146 174838 92382 175074
rect 100826 174218 101062 174454
rect 101146 174218 101382 174454
rect 100826 173898 101062 174134
rect 101146 173898 101382 174134
rect 109826 175158 110062 175394
rect 110146 175158 110382 175394
rect 109826 174838 110062 175074
rect 110146 174838 110382 175074
rect 118826 174218 119062 174454
rect 119146 174218 119382 174454
rect 118826 173898 119062 174134
rect 119146 173898 119382 174134
rect 127826 175158 128062 175394
rect 128146 175158 128382 175394
rect 127826 174838 128062 175074
rect 128146 174838 128382 175074
rect 136826 174218 137062 174454
rect 137146 174218 137382 174454
rect 136826 173898 137062 174134
rect 137146 173898 137382 174134
rect 145826 175158 146062 175394
rect 146146 175158 146382 175394
rect 145826 174838 146062 175074
rect 146146 174838 146382 175074
rect 154826 174218 155062 174454
rect 155146 174218 155382 174454
rect 154826 173898 155062 174134
rect 155146 173898 155382 174134
rect 163826 175158 164062 175394
rect 164146 175158 164382 175394
rect 163826 174838 164062 175074
rect 164146 174838 164382 175074
rect 172826 174218 173062 174454
rect 173146 174218 173382 174454
rect 172826 173898 173062 174134
rect 173146 173898 173382 174134
rect 181826 175158 182062 175394
rect 182146 175158 182382 175394
rect 181826 174838 182062 175074
rect 182146 174838 182382 175074
rect 190826 174218 191062 174454
rect 191146 174218 191382 174454
rect 190826 173898 191062 174134
rect 191146 173898 191382 174134
rect 199826 175158 200062 175394
rect 200146 175158 200382 175394
rect 199826 174838 200062 175074
rect 200146 174838 200382 175074
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 217826 175158 218062 175394
rect 218146 175158 218382 175394
rect 217826 174838 218062 175074
rect 218146 174838 218382 175074
rect 226826 174218 227062 174454
rect 227146 174218 227382 174454
rect 226826 173898 227062 174134
rect 227146 173898 227382 174134
rect 235826 175158 236062 175394
rect 236146 175158 236382 175394
rect 235826 174838 236062 175074
rect 236146 174838 236382 175074
rect 244826 174218 245062 174454
rect 245146 174218 245382 174454
rect 244826 173898 245062 174134
rect 245146 173898 245382 174134
rect 253826 175158 254062 175394
rect 254146 175158 254382 175394
rect 253826 174838 254062 175074
rect 254146 174838 254382 175074
rect 262826 174218 263062 174454
rect 263146 174218 263382 174454
rect 262826 173898 263062 174134
rect 263146 173898 263382 174134
rect 271826 175158 272062 175394
rect 272146 175158 272382 175394
rect 271826 174838 272062 175074
rect 272146 174838 272382 175074
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 289826 175158 290062 175394
rect 290146 175158 290382 175394
rect 289826 174838 290062 175074
rect 290146 174838 290382 175074
rect 298826 174218 299062 174454
rect 299146 174218 299382 174454
rect 298826 173898 299062 174134
rect 299146 173898 299382 174134
rect 307826 175158 308062 175394
rect 308146 175158 308382 175394
rect 307826 174838 308062 175074
rect 308146 174838 308382 175074
rect 316826 174218 317062 174454
rect 317146 174218 317382 174454
rect 316826 173898 317062 174134
rect 317146 173898 317382 174134
rect 325826 175158 326062 175394
rect 326146 175158 326382 175394
rect 325826 174838 326062 175074
rect 326146 174838 326382 175074
rect 334826 174218 335062 174454
rect 335146 174218 335382 174454
rect 334826 173898 335062 174134
rect 335146 173898 335382 174134
rect 343826 175158 344062 175394
rect 344146 175158 344382 175394
rect 343826 174838 344062 175074
rect 344146 174838 344382 175074
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 361826 175158 362062 175394
rect 362146 175158 362382 175394
rect 361826 174838 362062 175074
rect 362146 174838 362382 175074
rect 370826 174218 371062 174454
rect 371146 174218 371382 174454
rect 370826 173898 371062 174134
rect 371146 173898 371382 174134
rect 379826 175158 380062 175394
rect 380146 175158 380382 175394
rect 379826 174838 380062 175074
rect 380146 174838 380382 175074
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 397826 175158 398062 175394
rect 398146 175158 398382 175394
rect 397826 174838 398062 175074
rect 398146 174838 398382 175074
rect 406826 174218 407062 174454
rect 407146 174218 407382 174454
rect 406826 173898 407062 174134
rect 407146 173898 407382 174134
rect 415826 175158 416062 175394
rect 416146 175158 416382 175394
rect 415826 174838 416062 175074
rect 416146 174838 416382 175074
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 433826 175158 434062 175394
rect 434146 175158 434382 175394
rect 433826 174838 434062 175074
rect 434146 174838 434382 175074
rect 442826 174218 443062 174454
rect 443146 174218 443382 174454
rect 442826 173898 443062 174134
rect 443146 173898 443382 174134
rect 451826 175158 452062 175394
rect 452146 175158 452382 175394
rect 451826 174838 452062 175074
rect 452146 174838 452382 175074
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 469826 175158 470062 175394
rect 470146 175158 470382 175394
rect 469826 174838 470062 175074
rect 470146 174838 470382 175074
rect 478826 174218 479062 174454
rect 479146 174218 479382 174454
rect 478826 173898 479062 174134
rect 479146 173898 479382 174134
rect 487826 175158 488062 175394
rect 488146 175158 488382 175394
rect 487826 174838 488062 175074
rect 488146 174838 488382 175074
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 505826 175158 506062 175394
rect 506146 175158 506382 175394
rect 505826 174838 506062 175074
rect 506146 174838 506382 175074
rect 514826 174218 515062 174454
rect 515146 174218 515382 174454
rect 514826 173898 515062 174134
rect 515146 173898 515382 174134
rect 523826 175158 524062 175394
rect 524146 175158 524382 175394
rect 523826 174838 524062 175074
rect 524146 174838 524382 175074
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 541826 175158 542062 175394
rect 542146 175158 542382 175394
rect 541826 174838 542062 175074
rect 542146 174838 542382 175074
rect 550826 174218 551062 174454
rect 551146 174218 551382 174454
rect 550826 173898 551062 174134
rect 551146 173898 551382 174134
rect 19952 165218 20188 165454
rect 19952 164898 20188 165134
rect 25882 165218 26118 165454
rect 25882 164898 26118 165134
rect 31813 165218 32049 165454
rect 31813 164898 32049 165134
rect 46952 165218 47188 165454
rect 46952 164898 47188 165134
rect 52882 165218 53118 165454
rect 52882 164898 53118 165134
rect 58813 165218 59049 165454
rect 58813 164898 59049 165134
rect 73952 165218 74188 165454
rect 73952 164898 74188 165134
rect 79882 165218 80118 165454
rect 79882 164898 80118 165134
rect 85813 165218 86049 165454
rect 85813 164898 86049 165134
rect 100952 165218 101188 165454
rect 100952 164898 101188 165134
rect 106882 165218 107118 165454
rect 106882 164898 107118 165134
rect 112813 165218 113049 165454
rect 112813 164898 113049 165134
rect 127952 165218 128188 165454
rect 127952 164898 128188 165134
rect 133882 165218 134118 165454
rect 133882 164898 134118 165134
rect 139813 165218 140049 165454
rect 139813 164898 140049 165134
rect 154952 165218 155188 165454
rect 154952 164898 155188 165134
rect 160882 165218 161118 165454
rect 160882 164898 161118 165134
rect 166813 165218 167049 165454
rect 166813 164898 167049 165134
rect 181952 165218 182188 165454
rect 181952 164898 182188 165134
rect 187882 165218 188118 165454
rect 187882 164898 188118 165134
rect 193813 165218 194049 165454
rect 193813 164898 194049 165134
rect 208952 165218 209188 165454
rect 208952 164898 209188 165134
rect 214882 165218 215118 165454
rect 214882 164898 215118 165134
rect 220813 165218 221049 165454
rect 220813 164898 221049 165134
rect 235952 165218 236188 165454
rect 235952 164898 236188 165134
rect 241882 165218 242118 165454
rect 241882 164898 242118 165134
rect 247813 165218 248049 165454
rect 247813 164898 248049 165134
rect 262952 165218 263188 165454
rect 262952 164898 263188 165134
rect 268882 165218 269118 165454
rect 268882 164898 269118 165134
rect 274813 165218 275049 165454
rect 274813 164898 275049 165134
rect 289952 165218 290188 165454
rect 289952 164898 290188 165134
rect 295882 165218 296118 165454
rect 295882 164898 296118 165134
rect 301813 165218 302049 165454
rect 301813 164898 302049 165134
rect 316952 165218 317188 165454
rect 316952 164898 317188 165134
rect 322882 165218 323118 165454
rect 322882 164898 323118 165134
rect 328813 165218 329049 165454
rect 328813 164898 329049 165134
rect 343952 165218 344188 165454
rect 343952 164898 344188 165134
rect 349882 165218 350118 165454
rect 349882 164898 350118 165134
rect 355813 165218 356049 165454
rect 355813 164898 356049 165134
rect 370952 165218 371188 165454
rect 370952 164898 371188 165134
rect 376882 165218 377118 165454
rect 376882 164898 377118 165134
rect 382813 165218 383049 165454
rect 382813 164898 383049 165134
rect 397952 165218 398188 165454
rect 397952 164898 398188 165134
rect 403882 165218 404118 165454
rect 403882 164898 404118 165134
rect 409813 165218 410049 165454
rect 409813 164898 410049 165134
rect 424952 165218 425188 165454
rect 424952 164898 425188 165134
rect 430882 165218 431118 165454
rect 430882 164898 431118 165134
rect 436813 165218 437049 165454
rect 436813 164898 437049 165134
rect 451952 165218 452188 165454
rect 451952 164898 452188 165134
rect 457882 165218 458118 165454
rect 457882 164898 458118 165134
rect 463813 165218 464049 165454
rect 463813 164898 464049 165134
rect 478952 165218 479188 165454
rect 478952 164898 479188 165134
rect 484882 165218 485118 165454
rect 484882 164898 485118 165134
rect 490813 165218 491049 165454
rect 490813 164898 491049 165134
rect 505952 165218 506188 165454
rect 505952 164898 506188 165134
rect 511882 165218 512118 165454
rect 511882 164898 512118 165134
rect 517813 165218 518049 165454
rect 517813 164898 518049 165134
rect 532952 165218 533188 165454
rect 532952 164898 533188 165134
rect 538882 165218 539118 165454
rect 538882 164898 539118 165134
rect 544813 165218 545049 165454
rect 544813 164898 545049 165134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 22916 156218 23152 156454
rect 22916 155898 23152 156134
rect 28847 156218 29083 156454
rect 28847 155898 29083 156134
rect 49916 156218 50152 156454
rect 49916 155898 50152 156134
rect 55847 156218 56083 156454
rect 55847 155898 56083 156134
rect 76916 156218 77152 156454
rect 76916 155898 77152 156134
rect 82847 156218 83083 156454
rect 82847 155898 83083 156134
rect 103916 156218 104152 156454
rect 103916 155898 104152 156134
rect 109847 156218 110083 156454
rect 109847 155898 110083 156134
rect 130916 156218 131152 156454
rect 130916 155898 131152 156134
rect 136847 156218 137083 156454
rect 136847 155898 137083 156134
rect 157916 156218 158152 156454
rect 157916 155898 158152 156134
rect 163847 156218 164083 156454
rect 163847 155898 164083 156134
rect 184916 156218 185152 156454
rect 184916 155898 185152 156134
rect 190847 156218 191083 156454
rect 190847 155898 191083 156134
rect 211916 156218 212152 156454
rect 211916 155898 212152 156134
rect 217847 156218 218083 156454
rect 217847 155898 218083 156134
rect 238916 156218 239152 156454
rect 238916 155898 239152 156134
rect 244847 156218 245083 156454
rect 244847 155898 245083 156134
rect 265916 156218 266152 156454
rect 265916 155898 266152 156134
rect 271847 156218 272083 156454
rect 271847 155898 272083 156134
rect 292916 156218 293152 156454
rect 292916 155898 293152 156134
rect 298847 156218 299083 156454
rect 298847 155898 299083 156134
rect 319916 156218 320152 156454
rect 319916 155898 320152 156134
rect 325847 156218 326083 156454
rect 325847 155898 326083 156134
rect 346916 156218 347152 156454
rect 346916 155898 347152 156134
rect 352847 156218 353083 156454
rect 352847 155898 353083 156134
rect 373916 156218 374152 156454
rect 373916 155898 374152 156134
rect 379847 156218 380083 156454
rect 379847 155898 380083 156134
rect 400916 156218 401152 156454
rect 400916 155898 401152 156134
rect 406847 156218 407083 156454
rect 406847 155898 407083 156134
rect 427916 156218 428152 156454
rect 427916 155898 428152 156134
rect 433847 156218 434083 156454
rect 433847 155898 434083 156134
rect 454916 156218 455152 156454
rect 454916 155898 455152 156134
rect 460847 156218 461083 156454
rect 460847 155898 461083 156134
rect 481916 156218 482152 156454
rect 481916 155898 482152 156134
rect 487847 156218 488083 156454
rect 487847 155898 488083 156134
rect 508916 156218 509152 156454
rect 508916 155898 509152 156134
rect 514847 156218 515083 156454
rect 514847 155898 515083 156134
rect 535916 156218 536152 156454
rect 535916 155898 536152 156134
rect 541847 156218 542083 156454
rect 541847 155898 542083 156134
rect 19826 147218 20062 147454
rect 20146 147218 20382 147454
rect 19826 146898 20062 147134
rect 20146 146898 20382 147134
rect 28826 148158 29062 148394
rect 29146 148158 29382 148394
rect 28826 147838 29062 148074
rect 29146 147838 29382 148074
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 46826 148158 47062 148394
rect 47146 148158 47382 148394
rect 46826 147838 47062 148074
rect 47146 147838 47382 148074
rect 55826 147218 56062 147454
rect 56146 147218 56382 147454
rect 55826 146898 56062 147134
rect 56146 146898 56382 147134
rect 64826 148158 65062 148394
rect 65146 148158 65382 148394
rect 64826 147838 65062 148074
rect 65146 147838 65382 148074
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 82826 148158 83062 148394
rect 83146 148158 83382 148394
rect 82826 147838 83062 148074
rect 83146 147838 83382 148074
rect 91826 147218 92062 147454
rect 92146 147218 92382 147454
rect 91826 146898 92062 147134
rect 92146 146898 92382 147134
rect 100826 148158 101062 148394
rect 101146 148158 101382 148394
rect 100826 147838 101062 148074
rect 101146 147838 101382 148074
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 118826 148158 119062 148394
rect 119146 148158 119382 148394
rect 118826 147838 119062 148074
rect 119146 147838 119382 148074
rect 127826 147218 128062 147454
rect 128146 147218 128382 147454
rect 127826 146898 128062 147134
rect 128146 146898 128382 147134
rect 136826 148158 137062 148394
rect 137146 148158 137382 148394
rect 136826 147838 137062 148074
rect 137146 147838 137382 148074
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 154826 148158 155062 148394
rect 155146 148158 155382 148394
rect 154826 147838 155062 148074
rect 155146 147838 155382 148074
rect 163826 147218 164062 147454
rect 164146 147218 164382 147454
rect 163826 146898 164062 147134
rect 164146 146898 164382 147134
rect 172826 148158 173062 148394
rect 173146 148158 173382 148394
rect 172826 147838 173062 148074
rect 173146 147838 173382 148074
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 190826 148158 191062 148394
rect 191146 148158 191382 148394
rect 190826 147838 191062 148074
rect 191146 147838 191382 148074
rect 199826 147218 200062 147454
rect 200146 147218 200382 147454
rect 199826 146898 200062 147134
rect 200146 146898 200382 147134
rect 208826 148158 209062 148394
rect 209146 148158 209382 148394
rect 208826 147838 209062 148074
rect 209146 147838 209382 148074
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 226826 148158 227062 148394
rect 227146 148158 227382 148394
rect 226826 147838 227062 148074
rect 227146 147838 227382 148074
rect 235826 147218 236062 147454
rect 236146 147218 236382 147454
rect 235826 146898 236062 147134
rect 236146 146898 236382 147134
rect 244826 148158 245062 148394
rect 245146 148158 245382 148394
rect 244826 147838 245062 148074
rect 245146 147838 245382 148074
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 262826 148158 263062 148394
rect 263146 148158 263382 148394
rect 262826 147838 263062 148074
rect 263146 147838 263382 148074
rect 271826 147218 272062 147454
rect 272146 147218 272382 147454
rect 271826 146898 272062 147134
rect 272146 146898 272382 147134
rect 280826 148158 281062 148394
rect 281146 148158 281382 148394
rect 280826 147838 281062 148074
rect 281146 147838 281382 148074
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 298826 148158 299062 148394
rect 299146 148158 299382 148394
rect 298826 147838 299062 148074
rect 299146 147838 299382 148074
rect 307826 147218 308062 147454
rect 308146 147218 308382 147454
rect 307826 146898 308062 147134
rect 308146 146898 308382 147134
rect 316826 148158 317062 148394
rect 317146 148158 317382 148394
rect 316826 147838 317062 148074
rect 317146 147838 317382 148074
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 334826 148158 335062 148394
rect 335146 148158 335382 148394
rect 334826 147838 335062 148074
rect 335146 147838 335382 148074
rect 343826 147218 344062 147454
rect 344146 147218 344382 147454
rect 343826 146898 344062 147134
rect 344146 146898 344382 147134
rect 352826 148158 353062 148394
rect 353146 148158 353382 148394
rect 352826 147838 353062 148074
rect 353146 147838 353382 148074
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 370826 148158 371062 148394
rect 371146 148158 371382 148394
rect 370826 147838 371062 148074
rect 371146 147838 371382 148074
rect 379826 147218 380062 147454
rect 380146 147218 380382 147454
rect 379826 146898 380062 147134
rect 380146 146898 380382 147134
rect 388826 148158 389062 148394
rect 389146 148158 389382 148394
rect 388826 147838 389062 148074
rect 389146 147838 389382 148074
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 406826 148158 407062 148394
rect 407146 148158 407382 148394
rect 406826 147838 407062 148074
rect 407146 147838 407382 148074
rect 415826 147218 416062 147454
rect 416146 147218 416382 147454
rect 415826 146898 416062 147134
rect 416146 146898 416382 147134
rect 424826 148158 425062 148394
rect 425146 148158 425382 148394
rect 424826 147838 425062 148074
rect 425146 147838 425382 148074
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 442826 148158 443062 148394
rect 443146 148158 443382 148394
rect 442826 147838 443062 148074
rect 443146 147838 443382 148074
rect 451826 147218 452062 147454
rect 452146 147218 452382 147454
rect 451826 146898 452062 147134
rect 452146 146898 452382 147134
rect 460826 148158 461062 148394
rect 461146 148158 461382 148394
rect 460826 147838 461062 148074
rect 461146 147838 461382 148074
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 478826 148158 479062 148394
rect 479146 148158 479382 148394
rect 478826 147838 479062 148074
rect 479146 147838 479382 148074
rect 487826 147218 488062 147454
rect 488146 147218 488382 147454
rect 487826 146898 488062 147134
rect 488146 146898 488382 147134
rect 496826 148158 497062 148394
rect 497146 148158 497382 148394
rect 496826 147838 497062 148074
rect 497146 147838 497382 148074
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 514826 148158 515062 148394
rect 515146 148158 515382 148394
rect 514826 147838 515062 148074
rect 515146 147838 515382 148074
rect 523826 147218 524062 147454
rect 524146 147218 524382 147454
rect 523826 146898 524062 147134
rect 524146 146898 524382 147134
rect 532826 148158 533062 148394
rect 533146 148158 533382 148394
rect 532826 147838 533062 148074
rect 533146 147838 533382 148074
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 550826 148158 551062 148394
rect 551146 148158 551382 148394
rect 550826 147838 551062 148074
rect 551146 147838 551382 148074
rect 559826 147218 560062 147454
rect 560146 147218 560382 147454
rect 559826 146898 560062 147134
rect 560146 146898 560382 147134
rect 10826 138218 11062 138454
rect 11146 138218 11382 138454
rect 10826 137898 11062 138134
rect 11146 137898 11382 138134
rect 22916 138218 23152 138454
rect 22916 137898 23152 138134
rect 28847 138218 29083 138454
rect 28847 137898 29083 138134
rect 49916 138218 50152 138454
rect 49916 137898 50152 138134
rect 55847 138218 56083 138454
rect 55847 137898 56083 138134
rect 76916 138218 77152 138454
rect 76916 137898 77152 138134
rect 82847 138218 83083 138454
rect 82847 137898 83083 138134
rect 103916 138218 104152 138454
rect 103916 137898 104152 138134
rect 109847 138218 110083 138454
rect 109847 137898 110083 138134
rect 130916 138218 131152 138454
rect 130916 137898 131152 138134
rect 136847 138218 137083 138454
rect 136847 137898 137083 138134
rect 157916 138218 158152 138454
rect 157916 137898 158152 138134
rect 163847 138218 164083 138454
rect 163847 137898 164083 138134
rect 184916 138218 185152 138454
rect 184916 137898 185152 138134
rect 190847 138218 191083 138454
rect 190847 137898 191083 138134
rect 211916 138218 212152 138454
rect 211916 137898 212152 138134
rect 217847 138218 218083 138454
rect 217847 137898 218083 138134
rect 238916 138218 239152 138454
rect 238916 137898 239152 138134
rect 244847 138218 245083 138454
rect 244847 137898 245083 138134
rect 265916 138218 266152 138454
rect 265916 137898 266152 138134
rect 271847 138218 272083 138454
rect 271847 137898 272083 138134
rect 292916 138218 293152 138454
rect 292916 137898 293152 138134
rect 298847 138218 299083 138454
rect 298847 137898 299083 138134
rect 319916 138218 320152 138454
rect 319916 137898 320152 138134
rect 325847 138218 326083 138454
rect 325847 137898 326083 138134
rect 346916 138218 347152 138454
rect 346916 137898 347152 138134
rect 352847 138218 353083 138454
rect 352847 137898 353083 138134
rect 373916 138218 374152 138454
rect 373916 137898 374152 138134
rect 379847 138218 380083 138454
rect 379847 137898 380083 138134
rect 400916 138218 401152 138454
rect 400916 137898 401152 138134
rect 406847 138218 407083 138454
rect 406847 137898 407083 138134
rect 427916 138218 428152 138454
rect 427916 137898 428152 138134
rect 433847 138218 434083 138454
rect 433847 137898 434083 138134
rect 454916 138218 455152 138454
rect 454916 137898 455152 138134
rect 460847 138218 461083 138454
rect 460847 137898 461083 138134
rect 481916 138218 482152 138454
rect 481916 137898 482152 138134
rect 487847 138218 488083 138454
rect 487847 137898 488083 138134
rect 508916 138218 509152 138454
rect 508916 137898 509152 138134
rect 514847 138218 515083 138454
rect 514847 137898 515083 138134
rect 535916 138218 536152 138454
rect 535916 137898 536152 138134
rect 541847 138218 542083 138454
rect 541847 137898 542083 138134
rect 19952 129218 20188 129454
rect 19952 128898 20188 129134
rect 25882 129218 26118 129454
rect 25882 128898 26118 129134
rect 31813 129218 32049 129454
rect 31813 128898 32049 129134
rect 46952 129218 47188 129454
rect 46952 128898 47188 129134
rect 52882 129218 53118 129454
rect 52882 128898 53118 129134
rect 58813 129218 59049 129454
rect 58813 128898 59049 129134
rect 73952 129218 74188 129454
rect 73952 128898 74188 129134
rect 79882 129218 80118 129454
rect 79882 128898 80118 129134
rect 85813 129218 86049 129454
rect 85813 128898 86049 129134
rect 100952 129218 101188 129454
rect 100952 128898 101188 129134
rect 106882 129218 107118 129454
rect 106882 128898 107118 129134
rect 112813 129218 113049 129454
rect 112813 128898 113049 129134
rect 127952 129218 128188 129454
rect 127952 128898 128188 129134
rect 133882 129218 134118 129454
rect 133882 128898 134118 129134
rect 139813 129218 140049 129454
rect 139813 128898 140049 129134
rect 154952 129218 155188 129454
rect 154952 128898 155188 129134
rect 160882 129218 161118 129454
rect 160882 128898 161118 129134
rect 166813 129218 167049 129454
rect 166813 128898 167049 129134
rect 181952 129218 182188 129454
rect 181952 128898 182188 129134
rect 187882 129218 188118 129454
rect 187882 128898 188118 129134
rect 193813 129218 194049 129454
rect 193813 128898 194049 129134
rect 208952 129218 209188 129454
rect 208952 128898 209188 129134
rect 214882 129218 215118 129454
rect 214882 128898 215118 129134
rect 220813 129218 221049 129454
rect 220813 128898 221049 129134
rect 235952 129218 236188 129454
rect 235952 128898 236188 129134
rect 241882 129218 242118 129454
rect 241882 128898 242118 129134
rect 247813 129218 248049 129454
rect 247813 128898 248049 129134
rect 262952 129218 263188 129454
rect 262952 128898 263188 129134
rect 268882 129218 269118 129454
rect 268882 128898 269118 129134
rect 274813 129218 275049 129454
rect 274813 128898 275049 129134
rect 289952 129218 290188 129454
rect 289952 128898 290188 129134
rect 295882 129218 296118 129454
rect 295882 128898 296118 129134
rect 301813 129218 302049 129454
rect 301813 128898 302049 129134
rect 316952 129218 317188 129454
rect 316952 128898 317188 129134
rect 322882 129218 323118 129454
rect 322882 128898 323118 129134
rect 328813 129218 329049 129454
rect 328813 128898 329049 129134
rect 343952 129218 344188 129454
rect 343952 128898 344188 129134
rect 349882 129218 350118 129454
rect 349882 128898 350118 129134
rect 355813 129218 356049 129454
rect 355813 128898 356049 129134
rect 370952 129218 371188 129454
rect 370952 128898 371188 129134
rect 376882 129218 377118 129454
rect 376882 128898 377118 129134
rect 382813 129218 383049 129454
rect 382813 128898 383049 129134
rect 397952 129218 398188 129454
rect 397952 128898 398188 129134
rect 403882 129218 404118 129454
rect 403882 128898 404118 129134
rect 409813 129218 410049 129454
rect 409813 128898 410049 129134
rect 424952 129218 425188 129454
rect 424952 128898 425188 129134
rect 430882 129218 431118 129454
rect 430882 128898 431118 129134
rect 436813 129218 437049 129454
rect 436813 128898 437049 129134
rect 451952 129218 452188 129454
rect 451952 128898 452188 129134
rect 457882 129218 458118 129454
rect 457882 128898 458118 129134
rect 463813 129218 464049 129454
rect 463813 128898 464049 129134
rect 478952 129218 479188 129454
rect 478952 128898 479188 129134
rect 484882 129218 485118 129454
rect 484882 128898 485118 129134
rect 490813 129218 491049 129454
rect 490813 128898 491049 129134
rect 505952 129218 506188 129454
rect 505952 128898 506188 129134
rect 511882 129218 512118 129454
rect 511882 128898 512118 129134
rect 517813 129218 518049 129454
rect 517813 128898 518049 129134
rect 532952 129218 533188 129454
rect 532952 128898 533188 129134
rect 538882 129218 539118 129454
rect 538882 128898 539118 129134
rect 544813 129218 545049 129454
rect 544813 128898 545049 129134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 19826 121158 20062 121394
rect 20146 121158 20382 121394
rect 19826 120838 20062 121074
rect 20146 120838 20382 121074
rect 28826 120218 29062 120454
rect 29146 120218 29382 120454
rect 28826 119898 29062 120134
rect 29146 119898 29382 120134
rect 37826 121158 38062 121394
rect 38146 121158 38382 121394
rect 37826 120838 38062 121074
rect 38146 120838 38382 121074
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 55826 121158 56062 121394
rect 56146 121158 56382 121394
rect 55826 120838 56062 121074
rect 56146 120838 56382 121074
rect 64826 120218 65062 120454
rect 65146 120218 65382 120454
rect 64826 119898 65062 120134
rect 65146 119898 65382 120134
rect 73826 121158 74062 121394
rect 74146 121158 74382 121394
rect 73826 120838 74062 121074
rect 74146 120838 74382 121074
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 91826 121158 92062 121394
rect 92146 121158 92382 121394
rect 91826 120838 92062 121074
rect 92146 120838 92382 121074
rect 100826 120218 101062 120454
rect 101146 120218 101382 120454
rect 100826 119898 101062 120134
rect 101146 119898 101382 120134
rect 109826 121158 110062 121394
rect 110146 121158 110382 121394
rect 109826 120838 110062 121074
rect 110146 120838 110382 121074
rect 118826 120218 119062 120454
rect 119146 120218 119382 120454
rect 118826 119898 119062 120134
rect 119146 119898 119382 120134
rect 127826 121158 128062 121394
rect 128146 121158 128382 121394
rect 127826 120838 128062 121074
rect 128146 120838 128382 121074
rect 136826 120218 137062 120454
rect 137146 120218 137382 120454
rect 136826 119898 137062 120134
rect 137146 119898 137382 120134
rect 145826 121158 146062 121394
rect 146146 121158 146382 121394
rect 145826 120838 146062 121074
rect 146146 120838 146382 121074
rect 154826 120218 155062 120454
rect 155146 120218 155382 120454
rect 154826 119898 155062 120134
rect 155146 119898 155382 120134
rect 163826 121158 164062 121394
rect 164146 121158 164382 121394
rect 163826 120838 164062 121074
rect 164146 120838 164382 121074
rect 172826 120218 173062 120454
rect 173146 120218 173382 120454
rect 172826 119898 173062 120134
rect 173146 119898 173382 120134
rect 181826 121158 182062 121394
rect 182146 121158 182382 121394
rect 181826 120838 182062 121074
rect 182146 120838 182382 121074
rect 190826 120218 191062 120454
rect 191146 120218 191382 120454
rect 190826 119898 191062 120134
rect 191146 119898 191382 120134
rect 199826 121158 200062 121394
rect 200146 121158 200382 121394
rect 199826 120838 200062 121074
rect 200146 120838 200382 121074
rect 208826 120218 209062 120454
rect 209146 120218 209382 120454
rect 208826 119898 209062 120134
rect 209146 119898 209382 120134
rect 217826 121158 218062 121394
rect 218146 121158 218382 121394
rect 217826 120838 218062 121074
rect 218146 120838 218382 121074
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 235826 121158 236062 121394
rect 236146 121158 236382 121394
rect 235826 120838 236062 121074
rect 236146 120838 236382 121074
rect 244826 120218 245062 120454
rect 245146 120218 245382 120454
rect 244826 119898 245062 120134
rect 245146 119898 245382 120134
rect 253826 121158 254062 121394
rect 254146 121158 254382 121394
rect 253826 120838 254062 121074
rect 254146 120838 254382 121074
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 271826 121158 272062 121394
rect 272146 121158 272382 121394
rect 271826 120838 272062 121074
rect 272146 120838 272382 121074
rect 280826 120218 281062 120454
rect 281146 120218 281382 120454
rect 280826 119898 281062 120134
rect 281146 119898 281382 120134
rect 289826 121158 290062 121394
rect 290146 121158 290382 121394
rect 289826 120838 290062 121074
rect 290146 120838 290382 121074
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 307826 121158 308062 121394
rect 308146 121158 308382 121394
rect 307826 120838 308062 121074
rect 308146 120838 308382 121074
rect 316826 120218 317062 120454
rect 317146 120218 317382 120454
rect 316826 119898 317062 120134
rect 317146 119898 317382 120134
rect 325826 121158 326062 121394
rect 326146 121158 326382 121394
rect 325826 120838 326062 121074
rect 326146 120838 326382 121074
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 343826 121158 344062 121394
rect 344146 121158 344382 121394
rect 343826 120838 344062 121074
rect 344146 120838 344382 121074
rect 352826 120218 353062 120454
rect 353146 120218 353382 120454
rect 352826 119898 353062 120134
rect 353146 119898 353382 120134
rect 361826 121158 362062 121394
rect 362146 121158 362382 121394
rect 361826 120838 362062 121074
rect 362146 120838 362382 121074
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 379826 121158 380062 121394
rect 380146 121158 380382 121394
rect 379826 120838 380062 121074
rect 380146 120838 380382 121074
rect 388826 120218 389062 120454
rect 389146 120218 389382 120454
rect 388826 119898 389062 120134
rect 389146 119898 389382 120134
rect 397826 121158 398062 121394
rect 398146 121158 398382 121394
rect 397826 120838 398062 121074
rect 398146 120838 398382 121074
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 415826 121158 416062 121394
rect 416146 121158 416382 121394
rect 415826 120838 416062 121074
rect 416146 120838 416382 121074
rect 424826 120218 425062 120454
rect 425146 120218 425382 120454
rect 424826 119898 425062 120134
rect 425146 119898 425382 120134
rect 433826 121158 434062 121394
rect 434146 121158 434382 121394
rect 433826 120838 434062 121074
rect 434146 120838 434382 121074
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 451826 121158 452062 121394
rect 452146 121158 452382 121394
rect 451826 120838 452062 121074
rect 452146 120838 452382 121074
rect 460826 120218 461062 120454
rect 461146 120218 461382 120454
rect 460826 119898 461062 120134
rect 461146 119898 461382 120134
rect 469826 121158 470062 121394
rect 470146 121158 470382 121394
rect 469826 120838 470062 121074
rect 470146 120838 470382 121074
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 487826 121158 488062 121394
rect 488146 121158 488382 121394
rect 487826 120838 488062 121074
rect 488146 120838 488382 121074
rect 496826 120218 497062 120454
rect 497146 120218 497382 120454
rect 496826 119898 497062 120134
rect 497146 119898 497382 120134
rect 505826 121158 506062 121394
rect 506146 121158 506382 121394
rect 505826 120838 506062 121074
rect 506146 120838 506382 121074
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 523826 121158 524062 121394
rect 524146 121158 524382 121394
rect 523826 120838 524062 121074
rect 524146 120838 524382 121074
rect 532826 120218 533062 120454
rect 533146 120218 533382 120454
rect 532826 119898 533062 120134
rect 533146 119898 533382 120134
rect 541826 121158 542062 121394
rect 542146 121158 542382 121394
rect 541826 120838 542062 121074
rect 542146 120838 542382 121074
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 19952 111218 20188 111454
rect 19952 110898 20188 111134
rect 25882 111218 26118 111454
rect 25882 110898 26118 111134
rect 31813 111218 32049 111454
rect 31813 110898 32049 111134
rect 46952 111218 47188 111454
rect 46952 110898 47188 111134
rect 52882 111218 53118 111454
rect 52882 110898 53118 111134
rect 58813 111218 59049 111454
rect 58813 110898 59049 111134
rect 73952 111218 74188 111454
rect 73952 110898 74188 111134
rect 79882 111218 80118 111454
rect 79882 110898 80118 111134
rect 85813 111218 86049 111454
rect 85813 110898 86049 111134
rect 100952 111218 101188 111454
rect 100952 110898 101188 111134
rect 106882 111218 107118 111454
rect 106882 110898 107118 111134
rect 112813 111218 113049 111454
rect 112813 110898 113049 111134
rect 127952 111218 128188 111454
rect 127952 110898 128188 111134
rect 133882 111218 134118 111454
rect 133882 110898 134118 111134
rect 139813 111218 140049 111454
rect 139813 110898 140049 111134
rect 154952 111218 155188 111454
rect 154952 110898 155188 111134
rect 160882 111218 161118 111454
rect 160882 110898 161118 111134
rect 166813 111218 167049 111454
rect 166813 110898 167049 111134
rect 181952 111218 182188 111454
rect 181952 110898 182188 111134
rect 187882 111218 188118 111454
rect 187882 110898 188118 111134
rect 193813 111218 194049 111454
rect 193813 110898 194049 111134
rect 208952 111218 209188 111454
rect 208952 110898 209188 111134
rect 214882 111218 215118 111454
rect 214882 110898 215118 111134
rect 220813 111218 221049 111454
rect 220813 110898 221049 111134
rect 235952 111218 236188 111454
rect 235952 110898 236188 111134
rect 241882 111218 242118 111454
rect 241882 110898 242118 111134
rect 247813 111218 248049 111454
rect 247813 110898 248049 111134
rect 262952 111218 263188 111454
rect 262952 110898 263188 111134
rect 268882 111218 269118 111454
rect 268882 110898 269118 111134
rect 274813 111218 275049 111454
rect 274813 110898 275049 111134
rect 289952 111218 290188 111454
rect 289952 110898 290188 111134
rect 295882 111218 296118 111454
rect 295882 110898 296118 111134
rect 301813 111218 302049 111454
rect 301813 110898 302049 111134
rect 316952 111218 317188 111454
rect 316952 110898 317188 111134
rect 322882 111218 323118 111454
rect 322882 110898 323118 111134
rect 328813 111218 329049 111454
rect 328813 110898 329049 111134
rect 343952 111218 344188 111454
rect 343952 110898 344188 111134
rect 349882 111218 350118 111454
rect 349882 110898 350118 111134
rect 355813 111218 356049 111454
rect 355813 110898 356049 111134
rect 370952 111218 371188 111454
rect 370952 110898 371188 111134
rect 376882 111218 377118 111454
rect 376882 110898 377118 111134
rect 382813 111218 383049 111454
rect 382813 110898 383049 111134
rect 397952 111218 398188 111454
rect 397952 110898 398188 111134
rect 403882 111218 404118 111454
rect 403882 110898 404118 111134
rect 409813 111218 410049 111454
rect 409813 110898 410049 111134
rect 424952 111218 425188 111454
rect 424952 110898 425188 111134
rect 430882 111218 431118 111454
rect 430882 110898 431118 111134
rect 436813 111218 437049 111454
rect 436813 110898 437049 111134
rect 451952 111218 452188 111454
rect 451952 110898 452188 111134
rect 457882 111218 458118 111454
rect 457882 110898 458118 111134
rect 463813 111218 464049 111454
rect 463813 110898 464049 111134
rect 478952 111218 479188 111454
rect 478952 110898 479188 111134
rect 484882 111218 485118 111454
rect 484882 110898 485118 111134
rect 490813 111218 491049 111454
rect 490813 110898 491049 111134
rect 505952 111218 506188 111454
rect 505952 110898 506188 111134
rect 511882 111218 512118 111454
rect 511882 110898 512118 111134
rect 517813 111218 518049 111454
rect 517813 110898 518049 111134
rect 532952 111218 533188 111454
rect 532952 110898 533188 111134
rect 538882 111218 539118 111454
rect 538882 110898 539118 111134
rect 544813 111218 545049 111454
rect 544813 110898 545049 111134
rect 559826 111218 560062 111454
rect 560146 111218 560382 111454
rect 559826 110898 560062 111134
rect 560146 110898 560382 111134
rect 10826 102218 11062 102454
rect 11146 102218 11382 102454
rect 10826 101898 11062 102134
rect 11146 101898 11382 102134
rect 22916 102218 23152 102454
rect 22916 101898 23152 102134
rect 28847 102218 29083 102454
rect 28847 101898 29083 102134
rect 49916 102218 50152 102454
rect 49916 101898 50152 102134
rect 55847 102218 56083 102454
rect 55847 101898 56083 102134
rect 76916 102218 77152 102454
rect 76916 101898 77152 102134
rect 82847 102218 83083 102454
rect 82847 101898 83083 102134
rect 103916 102218 104152 102454
rect 103916 101898 104152 102134
rect 109847 102218 110083 102454
rect 109847 101898 110083 102134
rect 130916 102218 131152 102454
rect 130916 101898 131152 102134
rect 136847 102218 137083 102454
rect 136847 101898 137083 102134
rect 157916 102218 158152 102454
rect 157916 101898 158152 102134
rect 163847 102218 164083 102454
rect 163847 101898 164083 102134
rect 184916 102218 185152 102454
rect 184916 101898 185152 102134
rect 190847 102218 191083 102454
rect 190847 101898 191083 102134
rect 211916 102218 212152 102454
rect 211916 101898 212152 102134
rect 217847 102218 218083 102454
rect 217847 101898 218083 102134
rect 238916 102218 239152 102454
rect 238916 101898 239152 102134
rect 244847 102218 245083 102454
rect 244847 101898 245083 102134
rect 265916 102218 266152 102454
rect 265916 101898 266152 102134
rect 271847 102218 272083 102454
rect 271847 101898 272083 102134
rect 292916 102218 293152 102454
rect 292916 101898 293152 102134
rect 298847 102218 299083 102454
rect 298847 101898 299083 102134
rect 319916 102218 320152 102454
rect 319916 101898 320152 102134
rect 325847 102218 326083 102454
rect 325847 101898 326083 102134
rect 346916 102218 347152 102454
rect 346916 101898 347152 102134
rect 352847 102218 353083 102454
rect 352847 101898 353083 102134
rect 373916 102218 374152 102454
rect 373916 101898 374152 102134
rect 379847 102218 380083 102454
rect 379847 101898 380083 102134
rect 400916 102218 401152 102454
rect 400916 101898 401152 102134
rect 406847 102218 407083 102454
rect 406847 101898 407083 102134
rect 427916 102218 428152 102454
rect 427916 101898 428152 102134
rect 433847 102218 434083 102454
rect 433847 101898 434083 102134
rect 454916 102218 455152 102454
rect 454916 101898 455152 102134
rect 460847 102218 461083 102454
rect 460847 101898 461083 102134
rect 481916 102218 482152 102454
rect 481916 101898 482152 102134
rect 487847 102218 488083 102454
rect 487847 101898 488083 102134
rect 508916 102218 509152 102454
rect 508916 101898 509152 102134
rect 514847 102218 515083 102454
rect 514847 101898 515083 102134
rect 535916 102218 536152 102454
rect 535916 101898 536152 102134
rect 541847 102218 542083 102454
rect 541847 101898 542083 102134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 28826 94158 29062 94394
rect 29146 94158 29382 94394
rect 28826 93838 29062 94074
rect 29146 93838 29382 94074
rect 37826 93218 38062 93454
rect 38146 93218 38382 93454
rect 37826 92898 38062 93134
rect 38146 92898 38382 93134
rect 46826 94158 47062 94394
rect 47146 94158 47382 94394
rect 46826 93838 47062 94074
rect 47146 93838 47382 94074
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 64826 94158 65062 94394
rect 65146 94158 65382 94394
rect 64826 93838 65062 94074
rect 65146 93838 65382 94074
rect 73826 93218 74062 93454
rect 74146 93218 74382 93454
rect 73826 92898 74062 93134
rect 74146 92898 74382 93134
rect 82826 94158 83062 94394
rect 83146 94158 83382 94394
rect 82826 93838 83062 94074
rect 83146 93838 83382 94074
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 100826 94158 101062 94394
rect 101146 94158 101382 94394
rect 100826 93838 101062 94074
rect 101146 93838 101382 94074
rect 109826 93218 110062 93454
rect 110146 93218 110382 93454
rect 109826 92898 110062 93134
rect 110146 92898 110382 93134
rect 118826 94158 119062 94394
rect 119146 94158 119382 94394
rect 118826 93838 119062 94074
rect 119146 93838 119382 94074
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 136826 94158 137062 94394
rect 137146 94158 137382 94394
rect 136826 93838 137062 94074
rect 137146 93838 137382 94074
rect 145826 93218 146062 93454
rect 146146 93218 146382 93454
rect 145826 92898 146062 93134
rect 146146 92898 146382 93134
rect 154826 94158 155062 94394
rect 155146 94158 155382 94394
rect 154826 93838 155062 94074
rect 155146 93838 155382 94074
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 172826 94158 173062 94394
rect 173146 94158 173382 94394
rect 172826 93838 173062 94074
rect 173146 93838 173382 94074
rect 181826 93218 182062 93454
rect 182146 93218 182382 93454
rect 181826 92898 182062 93134
rect 182146 92898 182382 93134
rect 190826 94158 191062 94394
rect 191146 94158 191382 94394
rect 190826 93838 191062 94074
rect 191146 93838 191382 94074
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 208826 94158 209062 94394
rect 209146 94158 209382 94394
rect 208826 93838 209062 94074
rect 209146 93838 209382 94074
rect 217826 93218 218062 93454
rect 218146 93218 218382 93454
rect 217826 92898 218062 93134
rect 218146 92898 218382 93134
rect 226826 94158 227062 94394
rect 227146 94158 227382 94394
rect 226826 93838 227062 94074
rect 227146 93838 227382 94074
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 244826 94158 245062 94394
rect 245146 94158 245382 94394
rect 244826 93838 245062 94074
rect 245146 93838 245382 94074
rect 253826 93218 254062 93454
rect 254146 93218 254382 93454
rect 253826 92898 254062 93134
rect 254146 92898 254382 93134
rect 262826 94158 263062 94394
rect 263146 94158 263382 94394
rect 262826 93838 263062 94074
rect 263146 93838 263382 94074
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 280826 94158 281062 94394
rect 281146 94158 281382 94394
rect 280826 93838 281062 94074
rect 281146 93838 281382 94074
rect 289826 93218 290062 93454
rect 290146 93218 290382 93454
rect 289826 92898 290062 93134
rect 290146 92898 290382 93134
rect 298826 94158 299062 94394
rect 299146 94158 299382 94394
rect 298826 93838 299062 94074
rect 299146 93838 299382 94074
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 316826 94158 317062 94394
rect 317146 94158 317382 94394
rect 316826 93838 317062 94074
rect 317146 93838 317382 94074
rect 325826 93218 326062 93454
rect 326146 93218 326382 93454
rect 325826 92898 326062 93134
rect 326146 92898 326382 93134
rect 334826 94158 335062 94394
rect 335146 94158 335382 94394
rect 334826 93838 335062 94074
rect 335146 93838 335382 94074
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 352826 94158 353062 94394
rect 353146 94158 353382 94394
rect 352826 93838 353062 94074
rect 353146 93838 353382 94074
rect 361826 93218 362062 93454
rect 362146 93218 362382 93454
rect 361826 92898 362062 93134
rect 362146 92898 362382 93134
rect 370826 94158 371062 94394
rect 371146 94158 371382 94394
rect 370826 93838 371062 94074
rect 371146 93838 371382 94074
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 388826 94158 389062 94394
rect 389146 94158 389382 94394
rect 388826 93838 389062 94074
rect 389146 93838 389382 94074
rect 397826 93218 398062 93454
rect 398146 93218 398382 93454
rect 397826 92898 398062 93134
rect 398146 92898 398382 93134
rect 406826 94158 407062 94394
rect 407146 94158 407382 94394
rect 406826 93838 407062 94074
rect 407146 93838 407382 94074
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 424826 94158 425062 94394
rect 425146 94158 425382 94394
rect 424826 93838 425062 94074
rect 425146 93838 425382 94074
rect 433826 93218 434062 93454
rect 434146 93218 434382 93454
rect 433826 92898 434062 93134
rect 434146 92898 434382 93134
rect 442826 94158 443062 94394
rect 443146 94158 443382 94394
rect 442826 93838 443062 94074
rect 443146 93838 443382 94074
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 460826 94158 461062 94394
rect 461146 94158 461382 94394
rect 460826 93838 461062 94074
rect 461146 93838 461382 94074
rect 469826 93218 470062 93454
rect 470146 93218 470382 93454
rect 469826 92898 470062 93134
rect 470146 92898 470382 93134
rect 478826 94158 479062 94394
rect 479146 94158 479382 94394
rect 478826 93838 479062 94074
rect 479146 93838 479382 94074
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 496826 94158 497062 94394
rect 497146 94158 497382 94394
rect 496826 93838 497062 94074
rect 497146 93838 497382 94074
rect 505826 93218 506062 93454
rect 506146 93218 506382 93454
rect 505826 92898 506062 93134
rect 506146 92898 506382 93134
rect 514826 94158 515062 94394
rect 515146 94158 515382 94394
rect 514826 93838 515062 94074
rect 515146 93838 515382 94074
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 532826 94158 533062 94394
rect 533146 94158 533382 94394
rect 532826 93838 533062 94074
rect 533146 93838 533382 94074
rect 541826 93218 542062 93454
rect 542146 93218 542382 93454
rect 541826 92898 542062 93134
rect 542146 92898 542382 93134
rect 550826 94158 551062 94394
rect 551146 94158 551382 94394
rect 550826 93838 551062 94074
rect 551146 93838 551382 94074
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 22916 84218 23152 84454
rect 22916 83898 23152 84134
rect 28847 84218 29083 84454
rect 28847 83898 29083 84134
rect 49916 84218 50152 84454
rect 49916 83898 50152 84134
rect 55847 84218 56083 84454
rect 55847 83898 56083 84134
rect 76916 84218 77152 84454
rect 76916 83898 77152 84134
rect 82847 84218 83083 84454
rect 82847 83898 83083 84134
rect 103916 84218 104152 84454
rect 103916 83898 104152 84134
rect 109847 84218 110083 84454
rect 109847 83898 110083 84134
rect 130916 84218 131152 84454
rect 130916 83898 131152 84134
rect 136847 84218 137083 84454
rect 136847 83898 137083 84134
rect 157916 84218 158152 84454
rect 157916 83898 158152 84134
rect 163847 84218 164083 84454
rect 163847 83898 164083 84134
rect 184916 84218 185152 84454
rect 184916 83898 185152 84134
rect 190847 84218 191083 84454
rect 190847 83898 191083 84134
rect 211916 84218 212152 84454
rect 211916 83898 212152 84134
rect 217847 84218 218083 84454
rect 217847 83898 218083 84134
rect 238916 84218 239152 84454
rect 238916 83898 239152 84134
rect 244847 84218 245083 84454
rect 244847 83898 245083 84134
rect 265916 84218 266152 84454
rect 265916 83898 266152 84134
rect 271847 84218 272083 84454
rect 271847 83898 272083 84134
rect 292916 84218 293152 84454
rect 292916 83898 293152 84134
rect 298847 84218 299083 84454
rect 298847 83898 299083 84134
rect 319916 84218 320152 84454
rect 319916 83898 320152 84134
rect 325847 84218 326083 84454
rect 325847 83898 326083 84134
rect 346916 84218 347152 84454
rect 346916 83898 347152 84134
rect 352847 84218 353083 84454
rect 352847 83898 353083 84134
rect 373916 84218 374152 84454
rect 373916 83898 374152 84134
rect 379847 84218 380083 84454
rect 379847 83898 380083 84134
rect 400916 84218 401152 84454
rect 400916 83898 401152 84134
rect 406847 84218 407083 84454
rect 406847 83898 407083 84134
rect 427916 84218 428152 84454
rect 427916 83898 428152 84134
rect 433847 84218 434083 84454
rect 433847 83898 434083 84134
rect 454916 84218 455152 84454
rect 454916 83898 455152 84134
rect 460847 84218 461083 84454
rect 460847 83898 461083 84134
rect 481916 84218 482152 84454
rect 481916 83898 482152 84134
rect 487847 84218 488083 84454
rect 487847 83898 488083 84134
rect 508916 84218 509152 84454
rect 508916 83898 509152 84134
rect 514847 84218 515083 84454
rect 514847 83898 515083 84134
rect 535916 84218 536152 84454
rect 535916 83898 536152 84134
rect 541847 84218 542083 84454
rect 541847 83898 542083 84134
rect 19952 75218 20188 75454
rect 19952 74898 20188 75134
rect 25882 75218 26118 75454
rect 25882 74898 26118 75134
rect 31813 75218 32049 75454
rect 31813 74898 32049 75134
rect 46952 75218 47188 75454
rect 46952 74898 47188 75134
rect 52882 75218 53118 75454
rect 52882 74898 53118 75134
rect 58813 75218 59049 75454
rect 58813 74898 59049 75134
rect 73952 75218 74188 75454
rect 73952 74898 74188 75134
rect 79882 75218 80118 75454
rect 79882 74898 80118 75134
rect 85813 75218 86049 75454
rect 85813 74898 86049 75134
rect 100952 75218 101188 75454
rect 100952 74898 101188 75134
rect 106882 75218 107118 75454
rect 106882 74898 107118 75134
rect 112813 75218 113049 75454
rect 112813 74898 113049 75134
rect 127952 75218 128188 75454
rect 127952 74898 128188 75134
rect 133882 75218 134118 75454
rect 133882 74898 134118 75134
rect 139813 75218 140049 75454
rect 139813 74898 140049 75134
rect 154952 75218 155188 75454
rect 154952 74898 155188 75134
rect 160882 75218 161118 75454
rect 160882 74898 161118 75134
rect 166813 75218 167049 75454
rect 166813 74898 167049 75134
rect 181952 75218 182188 75454
rect 181952 74898 182188 75134
rect 187882 75218 188118 75454
rect 187882 74898 188118 75134
rect 193813 75218 194049 75454
rect 193813 74898 194049 75134
rect 208952 75218 209188 75454
rect 208952 74898 209188 75134
rect 214882 75218 215118 75454
rect 214882 74898 215118 75134
rect 220813 75218 221049 75454
rect 220813 74898 221049 75134
rect 235952 75218 236188 75454
rect 235952 74898 236188 75134
rect 241882 75218 242118 75454
rect 241882 74898 242118 75134
rect 247813 75218 248049 75454
rect 247813 74898 248049 75134
rect 262952 75218 263188 75454
rect 262952 74898 263188 75134
rect 268882 75218 269118 75454
rect 268882 74898 269118 75134
rect 274813 75218 275049 75454
rect 274813 74898 275049 75134
rect 289952 75218 290188 75454
rect 289952 74898 290188 75134
rect 295882 75218 296118 75454
rect 295882 74898 296118 75134
rect 301813 75218 302049 75454
rect 301813 74898 302049 75134
rect 316952 75218 317188 75454
rect 316952 74898 317188 75134
rect 322882 75218 323118 75454
rect 322882 74898 323118 75134
rect 328813 75218 329049 75454
rect 328813 74898 329049 75134
rect 343952 75218 344188 75454
rect 343952 74898 344188 75134
rect 349882 75218 350118 75454
rect 349882 74898 350118 75134
rect 355813 75218 356049 75454
rect 355813 74898 356049 75134
rect 370952 75218 371188 75454
rect 370952 74898 371188 75134
rect 376882 75218 377118 75454
rect 376882 74898 377118 75134
rect 382813 75218 383049 75454
rect 382813 74898 383049 75134
rect 397952 75218 398188 75454
rect 397952 74898 398188 75134
rect 403882 75218 404118 75454
rect 403882 74898 404118 75134
rect 409813 75218 410049 75454
rect 409813 74898 410049 75134
rect 424952 75218 425188 75454
rect 424952 74898 425188 75134
rect 430882 75218 431118 75454
rect 430882 74898 431118 75134
rect 436813 75218 437049 75454
rect 436813 74898 437049 75134
rect 451952 75218 452188 75454
rect 451952 74898 452188 75134
rect 457882 75218 458118 75454
rect 457882 74898 458118 75134
rect 463813 75218 464049 75454
rect 463813 74898 464049 75134
rect 478952 75218 479188 75454
rect 478952 74898 479188 75134
rect 484882 75218 485118 75454
rect 484882 74898 485118 75134
rect 490813 75218 491049 75454
rect 490813 74898 491049 75134
rect 505952 75218 506188 75454
rect 505952 74898 506188 75134
rect 511882 75218 512118 75454
rect 511882 74898 512118 75134
rect 517813 75218 518049 75454
rect 517813 74898 518049 75134
rect 532952 75218 533188 75454
rect 532952 74898 533188 75134
rect 538882 75218 539118 75454
rect 538882 74898 539118 75134
rect 544813 75218 545049 75454
rect 544813 74898 545049 75134
rect 559826 75218 560062 75454
rect 560146 75218 560382 75454
rect 559826 74898 560062 75134
rect 560146 74898 560382 75134
rect 10826 66218 11062 66454
rect 11146 66218 11382 66454
rect 10826 65898 11062 66134
rect 11146 65898 11382 66134
rect 19826 67158 20062 67394
rect 20146 67158 20382 67394
rect 19826 66838 20062 67074
rect 20146 66838 20382 67074
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 37826 67158 38062 67394
rect 38146 67158 38382 67394
rect 37826 66838 38062 67074
rect 38146 66838 38382 67074
rect 46826 66218 47062 66454
rect 47146 66218 47382 66454
rect 46826 65898 47062 66134
rect 47146 65898 47382 66134
rect 55826 67158 56062 67394
rect 56146 67158 56382 67394
rect 55826 66838 56062 67074
rect 56146 66838 56382 67074
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 73826 67158 74062 67394
rect 74146 67158 74382 67394
rect 73826 66838 74062 67074
rect 74146 66838 74382 67074
rect 82826 66218 83062 66454
rect 83146 66218 83382 66454
rect 82826 65898 83062 66134
rect 83146 65898 83382 66134
rect 91826 67158 92062 67394
rect 92146 67158 92382 67394
rect 91826 66838 92062 67074
rect 92146 66838 92382 67074
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 109826 67158 110062 67394
rect 110146 67158 110382 67394
rect 109826 66838 110062 67074
rect 110146 66838 110382 67074
rect 118826 66218 119062 66454
rect 119146 66218 119382 66454
rect 118826 65898 119062 66134
rect 119146 65898 119382 66134
rect 127826 67158 128062 67394
rect 128146 67158 128382 67394
rect 127826 66838 128062 67074
rect 128146 66838 128382 67074
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 145826 67158 146062 67394
rect 146146 67158 146382 67394
rect 145826 66838 146062 67074
rect 146146 66838 146382 67074
rect 154826 66218 155062 66454
rect 155146 66218 155382 66454
rect 154826 65898 155062 66134
rect 155146 65898 155382 66134
rect 163826 67158 164062 67394
rect 164146 67158 164382 67394
rect 163826 66838 164062 67074
rect 164146 66838 164382 67074
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 181826 67158 182062 67394
rect 182146 67158 182382 67394
rect 181826 66838 182062 67074
rect 182146 66838 182382 67074
rect 190826 66218 191062 66454
rect 191146 66218 191382 66454
rect 190826 65898 191062 66134
rect 191146 65898 191382 66134
rect 199826 67158 200062 67394
rect 200146 67158 200382 67394
rect 199826 66838 200062 67074
rect 200146 66838 200382 67074
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 217826 67158 218062 67394
rect 218146 67158 218382 67394
rect 217826 66838 218062 67074
rect 218146 66838 218382 67074
rect 226826 66218 227062 66454
rect 227146 66218 227382 66454
rect 226826 65898 227062 66134
rect 227146 65898 227382 66134
rect 235826 67158 236062 67394
rect 236146 67158 236382 67394
rect 235826 66838 236062 67074
rect 236146 66838 236382 67074
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 253826 67158 254062 67394
rect 254146 67158 254382 67394
rect 253826 66838 254062 67074
rect 254146 66838 254382 67074
rect 262826 66218 263062 66454
rect 263146 66218 263382 66454
rect 262826 65898 263062 66134
rect 263146 65898 263382 66134
rect 271826 67158 272062 67394
rect 272146 67158 272382 67394
rect 271826 66838 272062 67074
rect 272146 66838 272382 67074
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 289826 67158 290062 67394
rect 290146 67158 290382 67394
rect 289826 66838 290062 67074
rect 290146 66838 290382 67074
rect 298826 66218 299062 66454
rect 299146 66218 299382 66454
rect 298826 65898 299062 66134
rect 299146 65898 299382 66134
rect 307826 67158 308062 67394
rect 308146 67158 308382 67394
rect 307826 66838 308062 67074
rect 308146 66838 308382 67074
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 325826 67158 326062 67394
rect 326146 67158 326382 67394
rect 325826 66838 326062 67074
rect 326146 66838 326382 67074
rect 334826 66218 335062 66454
rect 335146 66218 335382 66454
rect 334826 65898 335062 66134
rect 335146 65898 335382 66134
rect 343826 67158 344062 67394
rect 344146 67158 344382 67394
rect 343826 66838 344062 67074
rect 344146 66838 344382 67074
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 361826 67158 362062 67394
rect 362146 67158 362382 67394
rect 361826 66838 362062 67074
rect 362146 66838 362382 67074
rect 370826 66218 371062 66454
rect 371146 66218 371382 66454
rect 370826 65898 371062 66134
rect 371146 65898 371382 66134
rect 379826 67158 380062 67394
rect 380146 67158 380382 67394
rect 379826 66838 380062 67074
rect 380146 66838 380382 67074
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 397826 67158 398062 67394
rect 398146 67158 398382 67394
rect 397826 66838 398062 67074
rect 398146 66838 398382 67074
rect 406826 66218 407062 66454
rect 407146 66218 407382 66454
rect 406826 65898 407062 66134
rect 407146 65898 407382 66134
rect 415826 67158 416062 67394
rect 416146 67158 416382 67394
rect 415826 66838 416062 67074
rect 416146 66838 416382 67074
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 433826 67158 434062 67394
rect 434146 67158 434382 67394
rect 433826 66838 434062 67074
rect 434146 66838 434382 67074
rect 442826 66218 443062 66454
rect 443146 66218 443382 66454
rect 442826 65898 443062 66134
rect 443146 65898 443382 66134
rect 451826 67158 452062 67394
rect 452146 67158 452382 67394
rect 451826 66838 452062 67074
rect 452146 66838 452382 67074
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 469826 67158 470062 67394
rect 470146 67158 470382 67394
rect 469826 66838 470062 67074
rect 470146 66838 470382 67074
rect 478826 66218 479062 66454
rect 479146 66218 479382 66454
rect 478826 65898 479062 66134
rect 479146 65898 479382 66134
rect 487826 67158 488062 67394
rect 488146 67158 488382 67394
rect 487826 66838 488062 67074
rect 488146 66838 488382 67074
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 505826 67158 506062 67394
rect 506146 67158 506382 67394
rect 505826 66838 506062 67074
rect 506146 66838 506382 67074
rect 514826 66218 515062 66454
rect 515146 66218 515382 66454
rect 514826 65898 515062 66134
rect 515146 65898 515382 66134
rect 523826 67158 524062 67394
rect 524146 67158 524382 67394
rect 523826 66838 524062 67074
rect 524146 66838 524382 67074
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 541826 67158 542062 67394
rect 542146 67158 542382 67394
rect 541826 66838 542062 67074
rect 542146 66838 542382 67074
rect 550826 66218 551062 66454
rect 551146 66218 551382 66454
rect 550826 65898 551062 66134
rect 551146 65898 551382 66134
rect 19952 57218 20188 57454
rect 19952 56898 20188 57134
rect 25882 57218 26118 57454
rect 25882 56898 26118 57134
rect 31813 57218 32049 57454
rect 31813 56898 32049 57134
rect 46952 57218 47188 57454
rect 46952 56898 47188 57134
rect 52882 57218 53118 57454
rect 52882 56898 53118 57134
rect 58813 57218 59049 57454
rect 58813 56898 59049 57134
rect 73952 57218 74188 57454
rect 73952 56898 74188 57134
rect 79882 57218 80118 57454
rect 79882 56898 80118 57134
rect 85813 57218 86049 57454
rect 85813 56898 86049 57134
rect 100952 57218 101188 57454
rect 100952 56898 101188 57134
rect 106882 57218 107118 57454
rect 106882 56898 107118 57134
rect 112813 57218 113049 57454
rect 112813 56898 113049 57134
rect 127952 57218 128188 57454
rect 127952 56898 128188 57134
rect 133882 57218 134118 57454
rect 133882 56898 134118 57134
rect 139813 57218 140049 57454
rect 139813 56898 140049 57134
rect 154952 57218 155188 57454
rect 154952 56898 155188 57134
rect 160882 57218 161118 57454
rect 160882 56898 161118 57134
rect 166813 57218 167049 57454
rect 166813 56898 167049 57134
rect 181952 57218 182188 57454
rect 181952 56898 182188 57134
rect 187882 57218 188118 57454
rect 187882 56898 188118 57134
rect 193813 57218 194049 57454
rect 193813 56898 194049 57134
rect 208952 57218 209188 57454
rect 208952 56898 209188 57134
rect 214882 57218 215118 57454
rect 214882 56898 215118 57134
rect 220813 57218 221049 57454
rect 220813 56898 221049 57134
rect 235952 57218 236188 57454
rect 235952 56898 236188 57134
rect 241882 57218 242118 57454
rect 241882 56898 242118 57134
rect 247813 57218 248049 57454
rect 247813 56898 248049 57134
rect 262952 57218 263188 57454
rect 262952 56898 263188 57134
rect 268882 57218 269118 57454
rect 268882 56898 269118 57134
rect 274813 57218 275049 57454
rect 274813 56898 275049 57134
rect 289952 57218 290188 57454
rect 289952 56898 290188 57134
rect 295882 57218 296118 57454
rect 295882 56898 296118 57134
rect 301813 57218 302049 57454
rect 301813 56898 302049 57134
rect 316952 57218 317188 57454
rect 316952 56898 317188 57134
rect 322882 57218 323118 57454
rect 322882 56898 323118 57134
rect 328813 57218 329049 57454
rect 328813 56898 329049 57134
rect 343952 57218 344188 57454
rect 343952 56898 344188 57134
rect 349882 57218 350118 57454
rect 349882 56898 350118 57134
rect 355813 57218 356049 57454
rect 355813 56898 356049 57134
rect 370952 57218 371188 57454
rect 370952 56898 371188 57134
rect 376882 57218 377118 57454
rect 376882 56898 377118 57134
rect 382813 57218 383049 57454
rect 382813 56898 383049 57134
rect 397952 57218 398188 57454
rect 397952 56898 398188 57134
rect 403882 57218 404118 57454
rect 403882 56898 404118 57134
rect 409813 57218 410049 57454
rect 409813 56898 410049 57134
rect 424952 57218 425188 57454
rect 424952 56898 425188 57134
rect 430882 57218 431118 57454
rect 430882 56898 431118 57134
rect 436813 57218 437049 57454
rect 436813 56898 437049 57134
rect 451952 57218 452188 57454
rect 451952 56898 452188 57134
rect 457882 57218 458118 57454
rect 457882 56898 458118 57134
rect 463813 57218 464049 57454
rect 463813 56898 464049 57134
rect 478952 57218 479188 57454
rect 478952 56898 479188 57134
rect 484882 57218 485118 57454
rect 484882 56898 485118 57134
rect 490813 57218 491049 57454
rect 490813 56898 491049 57134
rect 505952 57218 506188 57454
rect 505952 56898 506188 57134
rect 511882 57218 512118 57454
rect 511882 56898 512118 57134
rect 517813 57218 518049 57454
rect 517813 56898 518049 57134
rect 532952 57218 533188 57454
rect 532952 56898 533188 57134
rect 538882 57218 539118 57454
rect 538882 56898 539118 57134
rect 544813 57218 545049 57454
rect 544813 56898 545049 57134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 22916 48218 23152 48454
rect 22916 47898 23152 48134
rect 28847 48218 29083 48454
rect 28847 47898 29083 48134
rect 49916 48218 50152 48454
rect 49916 47898 50152 48134
rect 55847 48218 56083 48454
rect 55847 47898 56083 48134
rect 76916 48218 77152 48454
rect 76916 47898 77152 48134
rect 82847 48218 83083 48454
rect 82847 47898 83083 48134
rect 103916 48218 104152 48454
rect 103916 47898 104152 48134
rect 109847 48218 110083 48454
rect 109847 47898 110083 48134
rect 130916 48218 131152 48454
rect 130916 47898 131152 48134
rect 136847 48218 137083 48454
rect 136847 47898 137083 48134
rect 157916 48218 158152 48454
rect 157916 47898 158152 48134
rect 163847 48218 164083 48454
rect 163847 47898 164083 48134
rect 184916 48218 185152 48454
rect 184916 47898 185152 48134
rect 190847 48218 191083 48454
rect 190847 47898 191083 48134
rect 211916 48218 212152 48454
rect 211916 47898 212152 48134
rect 217847 48218 218083 48454
rect 217847 47898 218083 48134
rect 238916 48218 239152 48454
rect 238916 47898 239152 48134
rect 244847 48218 245083 48454
rect 244847 47898 245083 48134
rect 265916 48218 266152 48454
rect 265916 47898 266152 48134
rect 271847 48218 272083 48454
rect 271847 47898 272083 48134
rect 292916 48218 293152 48454
rect 292916 47898 293152 48134
rect 298847 48218 299083 48454
rect 298847 47898 299083 48134
rect 319916 48218 320152 48454
rect 319916 47898 320152 48134
rect 325847 48218 326083 48454
rect 325847 47898 326083 48134
rect 346916 48218 347152 48454
rect 346916 47898 347152 48134
rect 352847 48218 353083 48454
rect 352847 47898 353083 48134
rect 373916 48218 374152 48454
rect 373916 47898 374152 48134
rect 379847 48218 380083 48454
rect 379847 47898 380083 48134
rect 400916 48218 401152 48454
rect 400916 47898 401152 48134
rect 406847 48218 407083 48454
rect 406847 47898 407083 48134
rect 427916 48218 428152 48454
rect 427916 47898 428152 48134
rect 433847 48218 434083 48454
rect 433847 47898 434083 48134
rect 454916 48218 455152 48454
rect 454916 47898 455152 48134
rect 460847 48218 461083 48454
rect 460847 47898 461083 48134
rect 481916 48218 482152 48454
rect 481916 47898 482152 48134
rect 487847 48218 488083 48454
rect 487847 47898 488083 48134
rect 508916 48218 509152 48454
rect 508916 47898 509152 48134
rect 514847 48218 515083 48454
rect 514847 47898 515083 48134
rect 535916 48218 536152 48454
rect 535916 47898 536152 48134
rect 541847 48218 542083 48454
rect 541847 47898 542083 48134
rect 19826 39218 20062 39454
rect 20146 39218 20382 39454
rect 19826 38898 20062 39134
rect 20146 38898 20382 39134
rect 28826 40158 29062 40394
rect 29146 40158 29382 40394
rect 28826 39838 29062 40074
rect 29146 39838 29382 40074
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 46826 40158 47062 40394
rect 47146 40158 47382 40394
rect 46826 39838 47062 40074
rect 47146 39838 47382 40074
rect 55826 39218 56062 39454
rect 56146 39218 56382 39454
rect 55826 38898 56062 39134
rect 56146 38898 56382 39134
rect 64826 40158 65062 40394
rect 65146 40158 65382 40394
rect 64826 39838 65062 40074
rect 65146 39838 65382 40074
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 82826 40158 83062 40394
rect 83146 40158 83382 40394
rect 82826 39838 83062 40074
rect 83146 39838 83382 40074
rect 91826 39218 92062 39454
rect 92146 39218 92382 39454
rect 91826 38898 92062 39134
rect 92146 38898 92382 39134
rect 100826 40158 101062 40394
rect 101146 40158 101382 40394
rect 100826 39838 101062 40074
rect 101146 39838 101382 40074
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 118826 40158 119062 40394
rect 119146 40158 119382 40394
rect 118826 39838 119062 40074
rect 119146 39838 119382 40074
rect 127826 39218 128062 39454
rect 128146 39218 128382 39454
rect 127826 38898 128062 39134
rect 128146 38898 128382 39134
rect 136826 40158 137062 40394
rect 137146 40158 137382 40394
rect 136826 39838 137062 40074
rect 137146 39838 137382 40074
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 154826 40158 155062 40394
rect 155146 40158 155382 40394
rect 154826 39838 155062 40074
rect 155146 39838 155382 40074
rect 163826 39218 164062 39454
rect 164146 39218 164382 39454
rect 163826 38898 164062 39134
rect 164146 38898 164382 39134
rect 172826 40158 173062 40394
rect 173146 40158 173382 40394
rect 172826 39838 173062 40074
rect 173146 39838 173382 40074
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 190826 40158 191062 40394
rect 191146 40158 191382 40394
rect 190826 39838 191062 40074
rect 191146 39838 191382 40074
rect 199826 39218 200062 39454
rect 200146 39218 200382 39454
rect 199826 38898 200062 39134
rect 200146 38898 200382 39134
rect 208826 40158 209062 40394
rect 209146 40158 209382 40394
rect 208826 39838 209062 40074
rect 209146 39838 209382 40074
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 226826 40158 227062 40394
rect 227146 40158 227382 40394
rect 226826 39838 227062 40074
rect 227146 39838 227382 40074
rect 235826 39218 236062 39454
rect 236146 39218 236382 39454
rect 235826 38898 236062 39134
rect 236146 38898 236382 39134
rect 244826 40158 245062 40394
rect 245146 40158 245382 40394
rect 244826 39838 245062 40074
rect 245146 39838 245382 40074
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 262826 40158 263062 40394
rect 263146 40158 263382 40394
rect 262826 39838 263062 40074
rect 263146 39838 263382 40074
rect 271826 39218 272062 39454
rect 272146 39218 272382 39454
rect 271826 38898 272062 39134
rect 272146 38898 272382 39134
rect 280826 40158 281062 40394
rect 281146 40158 281382 40394
rect 280826 39838 281062 40074
rect 281146 39838 281382 40074
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 298826 40158 299062 40394
rect 299146 40158 299382 40394
rect 298826 39838 299062 40074
rect 299146 39838 299382 40074
rect 307826 39218 308062 39454
rect 308146 39218 308382 39454
rect 307826 38898 308062 39134
rect 308146 38898 308382 39134
rect 316826 40158 317062 40394
rect 317146 40158 317382 40394
rect 316826 39838 317062 40074
rect 317146 39838 317382 40074
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 334826 40158 335062 40394
rect 335146 40158 335382 40394
rect 334826 39838 335062 40074
rect 335146 39838 335382 40074
rect 343826 39218 344062 39454
rect 344146 39218 344382 39454
rect 343826 38898 344062 39134
rect 344146 38898 344382 39134
rect 352826 40158 353062 40394
rect 353146 40158 353382 40394
rect 352826 39838 353062 40074
rect 353146 39838 353382 40074
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 370826 40158 371062 40394
rect 371146 40158 371382 40394
rect 370826 39838 371062 40074
rect 371146 39838 371382 40074
rect 379826 39218 380062 39454
rect 380146 39218 380382 39454
rect 379826 38898 380062 39134
rect 380146 38898 380382 39134
rect 388826 40158 389062 40394
rect 389146 40158 389382 40394
rect 388826 39838 389062 40074
rect 389146 39838 389382 40074
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 406826 40158 407062 40394
rect 407146 40158 407382 40394
rect 406826 39838 407062 40074
rect 407146 39838 407382 40074
rect 415826 39218 416062 39454
rect 416146 39218 416382 39454
rect 415826 38898 416062 39134
rect 416146 38898 416382 39134
rect 424826 40158 425062 40394
rect 425146 40158 425382 40394
rect 424826 39838 425062 40074
rect 425146 39838 425382 40074
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 442826 40158 443062 40394
rect 443146 40158 443382 40394
rect 442826 39838 443062 40074
rect 443146 39838 443382 40074
rect 451826 39218 452062 39454
rect 452146 39218 452382 39454
rect 451826 38898 452062 39134
rect 452146 38898 452382 39134
rect 460826 40158 461062 40394
rect 461146 40158 461382 40394
rect 460826 39838 461062 40074
rect 461146 39838 461382 40074
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 478826 40158 479062 40394
rect 479146 40158 479382 40394
rect 478826 39838 479062 40074
rect 479146 39838 479382 40074
rect 487826 39218 488062 39454
rect 488146 39218 488382 39454
rect 487826 38898 488062 39134
rect 488146 38898 488382 39134
rect 496826 40158 497062 40394
rect 497146 40158 497382 40394
rect 496826 39838 497062 40074
rect 497146 39838 497382 40074
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 514826 40158 515062 40394
rect 515146 40158 515382 40394
rect 514826 39838 515062 40074
rect 515146 39838 515382 40074
rect 523826 39218 524062 39454
rect 524146 39218 524382 39454
rect 523826 38898 524062 39134
rect 524146 38898 524382 39134
rect 532826 40158 533062 40394
rect 533146 40158 533382 40394
rect 532826 39838 533062 40074
rect 533146 39838 533382 40074
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 550826 40158 551062 40394
rect 551146 40158 551382 40394
rect 550826 39838 551062 40074
rect 551146 39838 551382 40074
rect 559826 39218 560062 39454
rect 560146 39218 560382 39454
rect 559826 38898 560062 39134
rect 560146 38898 560382 39134
rect 10826 30218 11062 30454
rect 11146 30218 11382 30454
rect 10826 29898 11062 30134
rect 11146 29898 11382 30134
rect 22916 30218 23152 30454
rect 22916 29898 23152 30134
rect 28847 30218 29083 30454
rect 28847 29898 29083 30134
rect 49916 30218 50152 30454
rect 49916 29898 50152 30134
rect 55847 30218 56083 30454
rect 55847 29898 56083 30134
rect 76916 30218 77152 30454
rect 76916 29898 77152 30134
rect 82847 30218 83083 30454
rect 82847 29898 83083 30134
rect 103916 30218 104152 30454
rect 103916 29898 104152 30134
rect 109847 30218 110083 30454
rect 109847 29898 110083 30134
rect 130916 30218 131152 30454
rect 130916 29898 131152 30134
rect 136847 30218 137083 30454
rect 136847 29898 137083 30134
rect 157916 30218 158152 30454
rect 157916 29898 158152 30134
rect 163847 30218 164083 30454
rect 163847 29898 164083 30134
rect 184916 30218 185152 30454
rect 184916 29898 185152 30134
rect 190847 30218 191083 30454
rect 190847 29898 191083 30134
rect 211916 30218 212152 30454
rect 211916 29898 212152 30134
rect 217847 30218 218083 30454
rect 217847 29898 218083 30134
rect 238916 30218 239152 30454
rect 238916 29898 239152 30134
rect 244847 30218 245083 30454
rect 244847 29898 245083 30134
rect 265916 30218 266152 30454
rect 265916 29898 266152 30134
rect 271847 30218 272083 30454
rect 271847 29898 272083 30134
rect 292916 30218 293152 30454
rect 292916 29898 293152 30134
rect 298847 30218 299083 30454
rect 298847 29898 299083 30134
rect 319916 30218 320152 30454
rect 319916 29898 320152 30134
rect 325847 30218 326083 30454
rect 325847 29898 326083 30134
rect 346916 30218 347152 30454
rect 346916 29898 347152 30134
rect 352847 30218 353083 30454
rect 352847 29898 353083 30134
rect 373916 30218 374152 30454
rect 373916 29898 374152 30134
rect 379847 30218 380083 30454
rect 379847 29898 380083 30134
rect 400916 30218 401152 30454
rect 400916 29898 401152 30134
rect 406847 30218 407083 30454
rect 406847 29898 407083 30134
rect 427916 30218 428152 30454
rect 427916 29898 428152 30134
rect 433847 30218 434083 30454
rect 433847 29898 434083 30134
rect 454916 30218 455152 30454
rect 454916 29898 455152 30134
rect 460847 30218 461083 30454
rect 460847 29898 461083 30134
rect 481916 30218 482152 30454
rect 481916 29898 482152 30134
rect 487847 30218 488083 30454
rect 487847 29898 488083 30134
rect 508916 30218 509152 30454
rect 508916 29898 509152 30134
rect 514847 30218 515083 30454
rect 514847 29898 515083 30134
rect 535916 30218 536152 30454
rect 535916 29898 536152 30134
rect 541847 30218 542083 30454
rect 541847 29898 542083 30134
rect 19952 21218 20188 21454
rect 19952 20898 20188 21134
rect 25882 21218 26118 21454
rect 25882 20898 26118 21134
rect 31813 21218 32049 21454
rect 31813 20898 32049 21134
rect 46952 21218 47188 21454
rect 46952 20898 47188 21134
rect 52882 21218 53118 21454
rect 52882 20898 53118 21134
rect 58813 21218 59049 21454
rect 58813 20898 59049 21134
rect 73952 21218 74188 21454
rect 73952 20898 74188 21134
rect 79882 21218 80118 21454
rect 79882 20898 80118 21134
rect 85813 21218 86049 21454
rect 85813 20898 86049 21134
rect 100952 21218 101188 21454
rect 100952 20898 101188 21134
rect 106882 21218 107118 21454
rect 106882 20898 107118 21134
rect 112813 21218 113049 21454
rect 112813 20898 113049 21134
rect 127952 21218 128188 21454
rect 127952 20898 128188 21134
rect 133882 21218 134118 21454
rect 133882 20898 134118 21134
rect 139813 21218 140049 21454
rect 139813 20898 140049 21134
rect 154952 21218 155188 21454
rect 154952 20898 155188 21134
rect 160882 21218 161118 21454
rect 160882 20898 161118 21134
rect 166813 21218 167049 21454
rect 166813 20898 167049 21134
rect 181952 21218 182188 21454
rect 181952 20898 182188 21134
rect 187882 21218 188118 21454
rect 187882 20898 188118 21134
rect 193813 21218 194049 21454
rect 193813 20898 194049 21134
rect 208952 21218 209188 21454
rect 208952 20898 209188 21134
rect 214882 21218 215118 21454
rect 214882 20898 215118 21134
rect 220813 21218 221049 21454
rect 220813 20898 221049 21134
rect 235952 21218 236188 21454
rect 235952 20898 236188 21134
rect 241882 21218 242118 21454
rect 241882 20898 242118 21134
rect 247813 21218 248049 21454
rect 247813 20898 248049 21134
rect 262952 21218 263188 21454
rect 262952 20898 263188 21134
rect 268882 21218 269118 21454
rect 268882 20898 269118 21134
rect 274813 21218 275049 21454
rect 274813 20898 275049 21134
rect 289952 21218 290188 21454
rect 289952 20898 290188 21134
rect 295882 21218 296118 21454
rect 295882 20898 296118 21134
rect 301813 21218 302049 21454
rect 301813 20898 302049 21134
rect 316952 21218 317188 21454
rect 316952 20898 317188 21134
rect 322882 21218 323118 21454
rect 322882 20898 323118 21134
rect 328813 21218 329049 21454
rect 328813 20898 329049 21134
rect 343952 21218 344188 21454
rect 343952 20898 344188 21134
rect 349882 21218 350118 21454
rect 349882 20898 350118 21134
rect 355813 21218 356049 21454
rect 355813 20898 356049 21134
rect 370952 21218 371188 21454
rect 370952 20898 371188 21134
rect 376882 21218 377118 21454
rect 376882 20898 377118 21134
rect 382813 21218 383049 21454
rect 382813 20898 383049 21134
rect 397952 21218 398188 21454
rect 397952 20898 398188 21134
rect 403882 21218 404118 21454
rect 403882 20898 404118 21134
rect 409813 21218 410049 21454
rect 409813 20898 410049 21134
rect 424952 21218 425188 21454
rect 424952 20898 425188 21134
rect 430882 21218 431118 21454
rect 430882 20898 431118 21134
rect 436813 21218 437049 21454
rect 436813 20898 437049 21134
rect 451952 21218 452188 21454
rect 451952 20898 452188 21134
rect 457882 21218 458118 21454
rect 457882 20898 458118 21134
rect 463813 21218 464049 21454
rect 463813 20898 464049 21134
rect 478952 21218 479188 21454
rect 478952 20898 479188 21134
rect 484882 21218 485118 21454
rect 484882 20898 485118 21134
rect 490813 21218 491049 21454
rect 490813 20898 491049 21134
rect 505952 21218 506188 21454
rect 505952 20898 506188 21134
rect 511882 21218 512118 21454
rect 511882 20898 512118 21134
rect 517813 21218 518049 21454
rect 517813 20898 518049 21134
rect 532952 21218 533188 21454
rect 532952 20898 533188 21134
rect 538882 21218 539118 21454
rect 538882 20898 539118 21134
rect 544813 21218 545049 21454
rect 544813 20898 545049 21134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -1542 11062 -1306
rect 11146 -1542 11382 -1306
rect 10826 -1862 11062 -1626
rect 11146 -1862 11382 -1626
rect 19826 3218 20062 3454
rect 20146 3218 20382 3454
rect 19826 2898 20062 3134
rect 20146 2898 20382 3134
rect 19826 -582 20062 -346
rect 20146 -582 20382 -346
rect 19826 -902 20062 -666
rect 20146 -902 20382 -666
rect 28826 12218 29062 12454
rect 29146 12218 29382 12454
rect 28826 11898 29062 12134
rect 29146 11898 29382 12134
rect 28826 -1542 29062 -1306
rect 29146 -1542 29382 -1306
rect 28826 -1862 29062 -1626
rect 29146 -1862 29382 -1626
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -1542 47062 -1306
rect 47146 -1542 47382 -1306
rect 46826 -1862 47062 -1626
rect 47146 -1862 47382 -1626
rect 55826 3218 56062 3454
rect 56146 3218 56382 3454
rect 55826 2898 56062 3134
rect 56146 2898 56382 3134
rect 55826 -582 56062 -346
rect 56146 -582 56382 -346
rect 55826 -902 56062 -666
rect 56146 -902 56382 -666
rect 64826 12218 65062 12454
rect 65146 12218 65382 12454
rect 64826 11898 65062 12134
rect 65146 11898 65382 12134
rect 64826 -1542 65062 -1306
rect 65146 -1542 65382 -1306
rect 64826 -1862 65062 -1626
rect 65146 -1862 65382 -1626
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -1542 83062 -1306
rect 83146 -1542 83382 -1306
rect 82826 -1862 83062 -1626
rect 83146 -1862 83382 -1626
rect 91826 3218 92062 3454
rect 92146 3218 92382 3454
rect 91826 2898 92062 3134
rect 92146 2898 92382 3134
rect 91826 -582 92062 -346
rect 92146 -582 92382 -346
rect 91826 -902 92062 -666
rect 92146 -902 92382 -666
rect 100826 12218 101062 12454
rect 101146 12218 101382 12454
rect 100826 11898 101062 12134
rect 101146 11898 101382 12134
rect 100826 -1542 101062 -1306
rect 101146 -1542 101382 -1306
rect 100826 -1862 101062 -1626
rect 101146 -1862 101382 -1626
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -1542 119062 -1306
rect 119146 -1542 119382 -1306
rect 118826 -1862 119062 -1626
rect 119146 -1862 119382 -1626
rect 127826 3218 128062 3454
rect 128146 3218 128382 3454
rect 127826 2898 128062 3134
rect 128146 2898 128382 3134
rect 127826 -582 128062 -346
rect 128146 -582 128382 -346
rect 127826 -902 128062 -666
rect 128146 -902 128382 -666
rect 136826 12218 137062 12454
rect 137146 12218 137382 12454
rect 136826 11898 137062 12134
rect 137146 11898 137382 12134
rect 136826 -1542 137062 -1306
rect 137146 -1542 137382 -1306
rect 136826 -1862 137062 -1626
rect 137146 -1862 137382 -1626
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -1542 155062 -1306
rect 155146 -1542 155382 -1306
rect 154826 -1862 155062 -1626
rect 155146 -1862 155382 -1626
rect 163826 3218 164062 3454
rect 164146 3218 164382 3454
rect 163826 2898 164062 3134
rect 164146 2898 164382 3134
rect 163826 -582 164062 -346
rect 164146 -582 164382 -346
rect 163826 -902 164062 -666
rect 164146 -902 164382 -666
rect 172826 12218 173062 12454
rect 173146 12218 173382 12454
rect 172826 11898 173062 12134
rect 173146 11898 173382 12134
rect 172826 -1542 173062 -1306
rect 173146 -1542 173382 -1306
rect 172826 -1862 173062 -1626
rect 173146 -1862 173382 -1626
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -1542 191062 -1306
rect 191146 -1542 191382 -1306
rect 190826 -1862 191062 -1626
rect 191146 -1862 191382 -1626
rect 199826 3218 200062 3454
rect 200146 3218 200382 3454
rect 199826 2898 200062 3134
rect 200146 2898 200382 3134
rect 199826 -582 200062 -346
rect 200146 -582 200382 -346
rect 199826 -902 200062 -666
rect 200146 -902 200382 -666
rect 208826 12218 209062 12454
rect 209146 12218 209382 12454
rect 208826 11898 209062 12134
rect 209146 11898 209382 12134
rect 208826 -1542 209062 -1306
rect 209146 -1542 209382 -1306
rect 208826 -1862 209062 -1626
rect 209146 -1862 209382 -1626
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -1542 227062 -1306
rect 227146 -1542 227382 -1306
rect 226826 -1862 227062 -1626
rect 227146 -1862 227382 -1626
rect 235826 3218 236062 3454
rect 236146 3218 236382 3454
rect 235826 2898 236062 3134
rect 236146 2898 236382 3134
rect 235826 -582 236062 -346
rect 236146 -582 236382 -346
rect 235826 -902 236062 -666
rect 236146 -902 236382 -666
rect 244826 12218 245062 12454
rect 245146 12218 245382 12454
rect 244826 11898 245062 12134
rect 245146 11898 245382 12134
rect 244826 -1542 245062 -1306
rect 245146 -1542 245382 -1306
rect 244826 -1862 245062 -1626
rect 245146 -1862 245382 -1626
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -1542 263062 -1306
rect 263146 -1542 263382 -1306
rect 262826 -1862 263062 -1626
rect 263146 -1862 263382 -1626
rect 271826 3218 272062 3454
rect 272146 3218 272382 3454
rect 271826 2898 272062 3134
rect 272146 2898 272382 3134
rect 271826 -582 272062 -346
rect 272146 -582 272382 -346
rect 271826 -902 272062 -666
rect 272146 -902 272382 -666
rect 280826 12218 281062 12454
rect 281146 12218 281382 12454
rect 280826 11898 281062 12134
rect 281146 11898 281382 12134
rect 280826 -1542 281062 -1306
rect 281146 -1542 281382 -1306
rect 280826 -1862 281062 -1626
rect 281146 -1862 281382 -1626
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -1542 299062 -1306
rect 299146 -1542 299382 -1306
rect 298826 -1862 299062 -1626
rect 299146 -1862 299382 -1626
rect 307826 3218 308062 3454
rect 308146 3218 308382 3454
rect 307826 2898 308062 3134
rect 308146 2898 308382 3134
rect 307826 -582 308062 -346
rect 308146 -582 308382 -346
rect 307826 -902 308062 -666
rect 308146 -902 308382 -666
rect 316826 12218 317062 12454
rect 317146 12218 317382 12454
rect 316826 11898 317062 12134
rect 317146 11898 317382 12134
rect 316826 -1542 317062 -1306
rect 317146 -1542 317382 -1306
rect 316826 -1862 317062 -1626
rect 317146 -1862 317382 -1626
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -1542 335062 -1306
rect 335146 -1542 335382 -1306
rect 334826 -1862 335062 -1626
rect 335146 -1862 335382 -1626
rect 343826 3218 344062 3454
rect 344146 3218 344382 3454
rect 343826 2898 344062 3134
rect 344146 2898 344382 3134
rect 343826 -582 344062 -346
rect 344146 -582 344382 -346
rect 343826 -902 344062 -666
rect 344146 -902 344382 -666
rect 352826 12218 353062 12454
rect 353146 12218 353382 12454
rect 352826 11898 353062 12134
rect 353146 11898 353382 12134
rect 352826 -1542 353062 -1306
rect 353146 -1542 353382 -1306
rect 352826 -1862 353062 -1626
rect 353146 -1862 353382 -1626
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -1542 371062 -1306
rect 371146 -1542 371382 -1306
rect 370826 -1862 371062 -1626
rect 371146 -1862 371382 -1626
rect 379826 3218 380062 3454
rect 380146 3218 380382 3454
rect 379826 2898 380062 3134
rect 380146 2898 380382 3134
rect 379826 -582 380062 -346
rect 380146 -582 380382 -346
rect 379826 -902 380062 -666
rect 380146 -902 380382 -666
rect 388826 12218 389062 12454
rect 389146 12218 389382 12454
rect 388826 11898 389062 12134
rect 389146 11898 389382 12134
rect 388826 -1542 389062 -1306
rect 389146 -1542 389382 -1306
rect 388826 -1862 389062 -1626
rect 389146 -1862 389382 -1626
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -1542 407062 -1306
rect 407146 -1542 407382 -1306
rect 406826 -1862 407062 -1626
rect 407146 -1862 407382 -1626
rect 415826 3218 416062 3454
rect 416146 3218 416382 3454
rect 415826 2898 416062 3134
rect 416146 2898 416382 3134
rect 415826 -582 416062 -346
rect 416146 -582 416382 -346
rect 415826 -902 416062 -666
rect 416146 -902 416382 -666
rect 424826 12218 425062 12454
rect 425146 12218 425382 12454
rect 424826 11898 425062 12134
rect 425146 11898 425382 12134
rect 424826 -1542 425062 -1306
rect 425146 -1542 425382 -1306
rect 424826 -1862 425062 -1626
rect 425146 -1862 425382 -1626
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -1542 443062 -1306
rect 443146 -1542 443382 -1306
rect 442826 -1862 443062 -1626
rect 443146 -1862 443382 -1626
rect 451826 3218 452062 3454
rect 452146 3218 452382 3454
rect 451826 2898 452062 3134
rect 452146 2898 452382 3134
rect 451826 -582 452062 -346
rect 452146 -582 452382 -346
rect 451826 -902 452062 -666
rect 452146 -902 452382 -666
rect 460826 12218 461062 12454
rect 461146 12218 461382 12454
rect 460826 11898 461062 12134
rect 461146 11898 461382 12134
rect 460826 -1542 461062 -1306
rect 461146 -1542 461382 -1306
rect 460826 -1862 461062 -1626
rect 461146 -1862 461382 -1626
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -1542 479062 -1306
rect 479146 -1542 479382 -1306
rect 478826 -1862 479062 -1626
rect 479146 -1862 479382 -1626
rect 487826 3218 488062 3454
rect 488146 3218 488382 3454
rect 487826 2898 488062 3134
rect 488146 2898 488382 3134
rect 487826 -582 488062 -346
rect 488146 -582 488382 -346
rect 487826 -902 488062 -666
rect 488146 -902 488382 -666
rect 496826 12218 497062 12454
rect 497146 12218 497382 12454
rect 496826 11898 497062 12134
rect 497146 11898 497382 12134
rect 496826 -1542 497062 -1306
rect 497146 -1542 497382 -1306
rect 496826 -1862 497062 -1626
rect 497146 -1862 497382 -1626
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -1542 515062 -1306
rect 515146 -1542 515382 -1306
rect 514826 -1862 515062 -1626
rect 515146 -1862 515382 -1626
rect 523826 3218 524062 3454
rect 524146 3218 524382 3454
rect 523826 2898 524062 3134
rect 524146 2898 524382 3134
rect 523826 -582 524062 -346
rect 524146 -582 524382 -346
rect 523826 -902 524062 -666
rect 524146 -902 524382 -666
rect 532826 12218 533062 12454
rect 533146 12218 533382 12454
rect 532826 11898 533062 12134
rect 533146 11898 533382 12134
rect 532826 -1542 533062 -1306
rect 533146 -1542 533382 -1306
rect 532826 -1862 533062 -1626
rect 533146 -1862 533382 -1626
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -1542 551062 -1306
rect 551146 -1542 551382 -1306
rect 550826 -1862 551062 -1626
rect 551146 -1862 551382 -1626
rect 559826 3218 560062 3454
rect 560146 3218 560382 3454
rect 559826 2898 560062 3134
rect 560146 2898 560382 3134
rect 559826 -582 560062 -346
rect 560146 -582 560382 -346
rect 559826 -902 560062 -666
rect 560146 -902 560382 -666
rect 568826 705562 569062 705798
rect 569146 705562 569382 705798
rect 568826 705242 569062 705478
rect 569146 705242 569382 705478
rect 568826 696218 569062 696454
rect 569146 696218 569382 696454
rect 568826 695898 569062 696134
rect 569146 695898 569382 696134
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 660218 569062 660454
rect 569146 660218 569382 660454
rect 568826 659898 569062 660134
rect 569146 659898 569382 660134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 624218 569062 624454
rect 569146 624218 569382 624454
rect 568826 623898 569062 624134
rect 569146 623898 569382 624134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 588218 569062 588454
rect 569146 588218 569382 588454
rect 568826 587898 569062 588134
rect 569146 587898 569382 588134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 552218 569062 552454
rect 569146 552218 569382 552454
rect 568826 551898 569062 552134
rect 569146 551898 569382 552134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 516218 569062 516454
rect 569146 516218 569382 516454
rect 568826 515898 569062 516134
rect 569146 515898 569382 516134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 480218 569062 480454
rect 569146 480218 569382 480454
rect 568826 479898 569062 480134
rect 569146 479898 569382 480134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 444218 569062 444454
rect 569146 444218 569382 444454
rect 568826 443898 569062 444134
rect 569146 443898 569382 444134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 408218 569062 408454
rect 569146 408218 569382 408454
rect 568826 407898 569062 408134
rect 569146 407898 569382 408134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 372218 569062 372454
rect 569146 372218 569382 372454
rect 568826 371898 569062 372134
rect 569146 371898 569382 372134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 336218 569062 336454
rect 569146 336218 569382 336454
rect 568826 335898 569062 336134
rect 569146 335898 569382 336134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 300218 569062 300454
rect 569146 300218 569382 300454
rect 568826 299898 569062 300134
rect 569146 299898 569382 300134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 264218 569062 264454
rect 569146 264218 569382 264454
rect 568826 263898 569062 264134
rect 569146 263898 569382 264134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 228218 569062 228454
rect 569146 228218 569382 228454
rect 568826 227898 569062 228134
rect 569146 227898 569382 228134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 192218 569062 192454
rect 569146 192218 569382 192454
rect 568826 191898 569062 192134
rect 569146 191898 569382 192134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 156218 569062 156454
rect 569146 156218 569382 156454
rect 568826 155898 569062 156134
rect 569146 155898 569382 156134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 120218 569062 120454
rect 569146 120218 569382 120454
rect 568826 119898 569062 120134
rect 569146 119898 569382 120134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 84218 569062 84454
rect 569146 84218 569382 84454
rect 568826 83898 569062 84134
rect 569146 83898 569382 84134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 48218 569062 48454
rect 569146 48218 569382 48454
rect 568826 47898 569062 48134
rect 569146 47898 569382 48134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 12218 569062 12454
rect 569146 12218 569382 12454
rect 568826 11898 569062 12134
rect 569146 11898 569382 12134
rect 568826 -1542 569062 -1306
rect 569146 -1542 569382 -1306
rect 568826 -1862 569062 -1626
rect 569146 -1862 569382 -1626
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 669218 578062 669454
rect 578146 669218 578382 669454
rect 577826 668898 578062 669134
rect 578146 668898 578382 669134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 633218 578062 633454
rect 578146 633218 578382 633454
rect 577826 632898 578062 633134
rect 578146 632898 578382 633134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 597218 578062 597454
rect 578146 597218 578382 597454
rect 577826 596898 578062 597134
rect 578146 596898 578382 597134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 561218 578062 561454
rect 578146 561218 578382 561454
rect 577826 560898 578062 561134
rect 578146 560898 578382 561134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 525218 578062 525454
rect 578146 525218 578382 525454
rect 577826 524898 578062 525134
rect 578146 524898 578382 525134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 489218 578062 489454
rect 578146 489218 578382 489454
rect 577826 488898 578062 489134
rect 578146 488898 578382 489134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 453218 578062 453454
rect 578146 453218 578382 453454
rect 577826 452898 578062 453134
rect 578146 452898 578382 453134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 417218 578062 417454
rect 578146 417218 578382 417454
rect 577826 416898 578062 417134
rect 578146 416898 578382 417134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 381218 578062 381454
rect 578146 381218 578382 381454
rect 577826 380898 578062 381134
rect 578146 380898 578382 381134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 345218 578062 345454
rect 578146 345218 578382 345454
rect 577826 344898 578062 345134
rect 578146 344898 578382 345134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 309218 578062 309454
rect 578146 309218 578382 309454
rect 577826 308898 578062 309134
rect 578146 308898 578382 309134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 273218 578062 273454
rect 578146 273218 578382 273454
rect 577826 272898 578062 273134
rect 578146 272898 578382 273134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 237218 578062 237454
rect 578146 237218 578382 237454
rect 577826 236898 578062 237134
rect 578146 236898 578382 237134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 201218 578062 201454
rect 578146 201218 578382 201454
rect 577826 200898 578062 201134
rect 578146 200898 578382 201134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 165218 578062 165454
rect 578146 165218 578382 165454
rect 577826 164898 578062 165134
rect 578146 164898 578382 165134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 129218 578062 129454
rect 578146 129218 578382 129454
rect 577826 128898 578062 129134
rect 578146 128898 578382 129134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 93218 578062 93454
rect 578146 93218 578382 93454
rect 577826 92898 578062 93134
rect 578146 92898 578382 93134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 57218 578062 57454
rect 578146 57218 578382 57454
rect 577826 56898 578062 57134
rect 578146 56898 578382 57134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 21218 578062 21454
rect 578146 21218 578382 21454
rect 577826 20898 578062 21134
rect 578146 20898 578382 21134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 669218 585578 669454
rect 585662 669218 585898 669454
rect 585342 668898 585578 669134
rect 585662 668898 585898 669134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 633218 585578 633454
rect 585662 633218 585898 633454
rect 585342 632898 585578 633134
rect 585662 632898 585898 633134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 597218 585578 597454
rect 585662 597218 585898 597454
rect 585342 596898 585578 597134
rect 585662 596898 585898 597134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 561218 585578 561454
rect 585662 561218 585898 561454
rect 585342 560898 585578 561134
rect 585662 560898 585898 561134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 525218 585578 525454
rect 585662 525218 585898 525454
rect 585342 524898 585578 525134
rect 585662 524898 585898 525134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 489218 585578 489454
rect 585662 489218 585898 489454
rect 585342 488898 585578 489134
rect 585662 488898 585898 489134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 453218 585578 453454
rect 585662 453218 585898 453454
rect 585342 452898 585578 453134
rect 585662 452898 585898 453134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 417218 585578 417454
rect 585662 417218 585898 417454
rect 585342 416898 585578 417134
rect 585662 416898 585898 417134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 381218 585578 381454
rect 585662 381218 585898 381454
rect 585342 380898 585578 381134
rect 585662 380898 585898 381134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 345218 585578 345454
rect 585662 345218 585898 345454
rect 585342 344898 585578 345134
rect 585662 344898 585898 345134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 309218 585578 309454
rect 585662 309218 585898 309454
rect 585342 308898 585578 309134
rect 585662 308898 585898 309134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 273218 585578 273454
rect 585662 273218 585898 273454
rect 585342 272898 585578 273134
rect 585662 272898 585898 273134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 237218 585578 237454
rect 585662 237218 585898 237454
rect 585342 236898 585578 237134
rect 585662 236898 585898 237134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 201218 585578 201454
rect 585662 201218 585898 201454
rect 585342 200898 585578 201134
rect 585662 200898 585898 201134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 165218 585578 165454
rect 585662 165218 585898 165454
rect 585342 164898 585578 165134
rect 585662 164898 585898 165134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 129218 585578 129454
rect 585662 129218 585898 129454
rect 585342 128898 585578 129134
rect 585662 128898 585898 129134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 93218 585578 93454
rect 585662 93218 585898 93454
rect 585342 92898 585578 93134
rect 585662 92898 585898 93134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 57218 585578 57454
rect 585662 57218 585898 57454
rect 585342 56898 585578 57134
rect 585662 56898 585898 57134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 21218 585578 21454
rect 585662 21218 585898 21454
rect 585342 20898 585578 21134
rect 585662 20898 585898 21134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 696218 586538 696454
rect 586622 696218 586858 696454
rect 586302 695898 586538 696134
rect 586622 695898 586858 696134
rect 586302 678218 586538 678454
rect 586622 678218 586858 678454
rect 586302 677898 586538 678134
rect 586622 677898 586858 678134
rect 586302 660218 586538 660454
rect 586622 660218 586858 660454
rect 586302 659898 586538 660134
rect 586622 659898 586858 660134
rect 586302 642218 586538 642454
rect 586622 642218 586858 642454
rect 586302 641898 586538 642134
rect 586622 641898 586858 642134
rect 586302 624218 586538 624454
rect 586622 624218 586858 624454
rect 586302 623898 586538 624134
rect 586622 623898 586858 624134
rect 586302 606218 586538 606454
rect 586622 606218 586858 606454
rect 586302 605898 586538 606134
rect 586622 605898 586858 606134
rect 586302 588218 586538 588454
rect 586622 588218 586858 588454
rect 586302 587898 586538 588134
rect 586622 587898 586858 588134
rect 586302 570218 586538 570454
rect 586622 570218 586858 570454
rect 586302 569898 586538 570134
rect 586622 569898 586858 570134
rect 586302 552218 586538 552454
rect 586622 552218 586858 552454
rect 586302 551898 586538 552134
rect 586622 551898 586858 552134
rect 586302 534218 586538 534454
rect 586622 534218 586858 534454
rect 586302 533898 586538 534134
rect 586622 533898 586858 534134
rect 586302 516218 586538 516454
rect 586622 516218 586858 516454
rect 586302 515898 586538 516134
rect 586622 515898 586858 516134
rect 586302 498218 586538 498454
rect 586622 498218 586858 498454
rect 586302 497898 586538 498134
rect 586622 497898 586858 498134
rect 586302 480218 586538 480454
rect 586622 480218 586858 480454
rect 586302 479898 586538 480134
rect 586622 479898 586858 480134
rect 586302 462218 586538 462454
rect 586622 462218 586858 462454
rect 586302 461898 586538 462134
rect 586622 461898 586858 462134
rect 586302 444218 586538 444454
rect 586622 444218 586858 444454
rect 586302 443898 586538 444134
rect 586622 443898 586858 444134
rect 586302 426218 586538 426454
rect 586622 426218 586858 426454
rect 586302 425898 586538 426134
rect 586622 425898 586858 426134
rect 586302 408218 586538 408454
rect 586622 408218 586858 408454
rect 586302 407898 586538 408134
rect 586622 407898 586858 408134
rect 586302 390218 586538 390454
rect 586622 390218 586858 390454
rect 586302 389898 586538 390134
rect 586622 389898 586858 390134
rect 586302 372218 586538 372454
rect 586622 372218 586858 372454
rect 586302 371898 586538 372134
rect 586622 371898 586858 372134
rect 586302 354218 586538 354454
rect 586622 354218 586858 354454
rect 586302 353898 586538 354134
rect 586622 353898 586858 354134
rect 586302 336218 586538 336454
rect 586622 336218 586858 336454
rect 586302 335898 586538 336134
rect 586622 335898 586858 336134
rect 586302 318218 586538 318454
rect 586622 318218 586858 318454
rect 586302 317898 586538 318134
rect 586622 317898 586858 318134
rect 586302 300218 586538 300454
rect 586622 300218 586858 300454
rect 586302 299898 586538 300134
rect 586622 299898 586858 300134
rect 586302 282218 586538 282454
rect 586622 282218 586858 282454
rect 586302 281898 586538 282134
rect 586622 281898 586858 282134
rect 586302 264218 586538 264454
rect 586622 264218 586858 264454
rect 586302 263898 586538 264134
rect 586622 263898 586858 264134
rect 586302 246218 586538 246454
rect 586622 246218 586858 246454
rect 586302 245898 586538 246134
rect 586622 245898 586858 246134
rect 586302 228218 586538 228454
rect 586622 228218 586858 228454
rect 586302 227898 586538 228134
rect 586622 227898 586858 228134
rect 586302 210218 586538 210454
rect 586622 210218 586858 210454
rect 586302 209898 586538 210134
rect 586622 209898 586858 210134
rect 586302 192218 586538 192454
rect 586622 192218 586858 192454
rect 586302 191898 586538 192134
rect 586622 191898 586858 192134
rect 586302 174218 586538 174454
rect 586622 174218 586858 174454
rect 586302 173898 586538 174134
rect 586622 173898 586858 174134
rect 586302 156218 586538 156454
rect 586622 156218 586858 156454
rect 586302 155898 586538 156134
rect 586622 155898 586858 156134
rect 586302 138218 586538 138454
rect 586622 138218 586858 138454
rect 586302 137898 586538 138134
rect 586622 137898 586858 138134
rect 586302 120218 586538 120454
rect 586622 120218 586858 120454
rect 586302 119898 586538 120134
rect 586622 119898 586858 120134
rect 586302 102218 586538 102454
rect 586622 102218 586858 102454
rect 586302 101898 586538 102134
rect 586622 101898 586858 102134
rect 586302 84218 586538 84454
rect 586622 84218 586858 84454
rect 586302 83898 586538 84134
rect 586622 83898 586858 84134
rect 586302 66218 586538 66454
rect 586622 66218 586858 66454
rect 586302 65898 586538 66134
rect 586622 65898 586858 66134
rect 586302 48218 586538 48454
rect 586622 48218 586858 48454
rect 586302 47898 586538 48134
rect 586622 47898 586858 48134
rect 586302 30218 586538 30454
rect 586622 30218 586858 30454
rect 586302 29898 586538 30134
rect 586622 29898 586858 30134
rect 586302 12218 586538 12454
rect 586622 12218 586858 12454
rect 586302 11898 586538 12134
rect 586622 11898 586858 12134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
<< metal5 >>
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 10826 705798
rect 11062 705562 11146 705798
rect 11382 705562 28826 705798
rect 29062 705562 29146 705798
rect 29382 705562 46826 705798
rect 47062 705562 47146 705798
rect 47382 705562 64826 705798
rect 65062 705562 65146 705798
rect 65382 705562 82826 705798
rect 83062 705562 83146 705798
rect 83382 705562 100826 705798
rect 101062 705562 101146 705798
rect 101382 705562 118826 705798
rect 119062 705562 119146 705798
rect 119382 705562 136826 705798
rect 137062 705562 137146 705798
rect 137382 705562 154826 705798
rect 155062 705562 155146 705798
rect 155382 705562 172826 705798
rect 173062 705562 173146 705798
rect 173382 705562 190826 705798
rect 191062 705562 191146 705798
rect 191382 705562 208826 705798
rect 209062 705562 209146 705798
rect 209382 705562 226826 705798
rect 227062 705562 227146 705798
rect 227382 705562 244826 705798
rect 245062 705562 245146 705798
rect 245382 705562 262826 705798
rect 263062 705562 263146 705798
rect 263382 705562 280826 705798
rect 281062 705562 281146 705798
rect 281382 705562 298826 705798
rect 299062 705562 299146 705798
rect 299382 705562 316826 705798
rect 317062 705562 317146 705798
rect 317382 705562 334826 705798
rect 335062 705562 335146 705798
rect 335382 705562 352826 705798
rect 353062 705562 353146 705798
rect 353382 705562 370826 705798
rect 371062 705562 371146 705798
rect 371382 705562 388826 705798
rect 389062 705562 389146 705798
rect 389382 705562 406826 705798
rect 407062 705562 407146 705798
rect 407382 705562 424826 705798
rect 425062 705562 425146 705798
rect 425382 705562 442826 705798
rect 443062 705562 443146 705798
rect 443382 705562 460826 705798
rect 461062 705562 461146 705798
rect 461382 705562 478826 705798
rect 479062 705562 479146 705798
rect 479382 705562 496826 705798
rect 497062 705562 497146 705798
rect 497382 705562 514826 705798
rect 515062 705562 515146 705798
rect 515382 705562 532826 705798
rect 533062 705562 533146 705798
rect 533382 705562 550826 705798
rect 551062 705562 551146 705798
rect 551382 705562 568826 705798
rect 569062 705562 569146 705798
rect 569382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 10826 705478
rect 11062 705242 11146 705478
rect 11382 705242 28826 705478
rect 29062 705242 29146 705478
rect 29382 705242 46826 705478
rect 47062 705242 47146 705478
rect 47382 705242 64826 705478
rect 65062 705242 65146 705478
rect 65382 705242 82826 705478
rect 83062 705242 83146 705478
rect 83382 705242 100826 705478
rect 101062 705242 101146 705478
rect 101382 705242 118826 705478
rect 119062 705242 119146 705478
rect 119382 705242 136826 705478
rect 137062 705242 137146 705478
rect 137382 705242 154826 705478
rect 155062 705242 155146 705478
rect 155382 705242 172826 705478
rect 173062 705242 173146 705478
rect 173382 705242 190826 705478
rect 191062 705242 191146 705478
rect 191382 705242 208826 705478
rect 209062 705242 209146 705478
rect 209382 705242 226826 705478
rect 227062 705242 227146 705478
rect 227382 705242 244826 705478
rect 245062 705242 245146 705478
rect 245382 705242 262826 705478
rect 263062 705242 263146 705478
rect 263382 705242 280826 705478
rect 281062 705242 281146 705478
rect 281382 705242 298826 705478
rect 299062 705242 299146 705478
rect 299382 705242 316826 705478
rect 317062 705242 317146 705478
rect 317382 705242 334826 705478
rect 335062 705242 335146 705478
rect 335382 705242 352826 705478
rect 353062 705242 353146 705478
rect 353382 705242 370826 705478
rect 371062 705242 371146 705478
rect 371382 705242 388826 705478
rect 389062 705242 389146 705478
rect 389382 705242 406826 705478
rect 407062 705242 407146 705478
rect 407382 705242 424826 705478
rect 425062 705242 425146 705478
rect 425382 705242 442826 705478
rect 443062 705242 443146 705478
rect 443382 705242 460826 705478
rect 461062 705242 461146 705478
rect 461382 705242 478826 705478
rect 479062 705242 479146 705478
rect 479382 705242 496826 705478
rect 497062 705242 497146 705478
rect 497382 705242 514826 705478
rect 515062 705242 515146 705478
rect 515382 705242 532826 705478
rect 533062 705242 533146 705478
rect 533382 705242 550826 705478
rect 551062 705242 551146 705478
rect 551382 705242 568826 705478
rect 569062 705242 569146 705478
rect 569382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 19826 704838
rect 20062 704602 20146 704838
rect 20382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 55826 704838
rect 56062 704602 56146 704838
rect 56382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 91826 704838
rect 92062 704602 92146 704838
rect 92382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 127826 704838
rect 128062 704602 128146 704838
rect 128382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 163826 704838
rect 164062 704602 164146 704838
rect 164382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 199826 704838
rect 200062 704602 200146 704838
rect 200382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 235826 704838
rect 236062 704602 236146 704838
rect 236382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 271826 704838
rect 272062 704602 272146 704838
rect 272382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 307826 704838
rect 308062 704602 308146 704838
rect 308382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 343826 704838
rect 344062 704602 344146 704838
rect 344382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 379826 704838
rect 380062 704602 380146 704838
rect 380382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 415826 704838
rect 416062 704602 416146 704838
rect 416382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 451826 704838
rect 452062 704602 452146 704838
rect 452382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 487826 704838
rect 488062 704602 488146 704838
rect 488382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 523826 704838
rect 524062 704602 524146 704838
rect 524382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 559826 704838
rect 560062 704602 560146 704838
rect 560382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 19826 704518
rect 20062 704282 20146 704518
rect 20382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 55826 704518
rect 56062 704282 56146 704518
rect 56382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 91826 704518
rect 92062 704282 92146 704518
rect 92382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 127826 704518
rect 128062 704282 128146 704518
rect 128382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 163826 704518
rect 164062 704282 164146 704518
rect 164382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 199826 704518
rect 200062 704282 200146 704518
rect 200382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 235826 704518
rect 236062 704282 236146 704518
rect 236382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 271826 704518
rect 272062 704282 272146 704518
rect 272382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 307826 704518
rect 308062 704282 308146 704518
rect 308382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 343826 704518
rect 344062 704282 344146 704518
rect 344382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 379826 704518
rect 380062 704282 380146 704518
rect 380382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 415826 704518
rect 416062 704282 416146 704518
rect 416382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 451826 704518
rect 452062 704282 452146 704518
rect 452382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 487826 704518
rect 488062 704282 488146 704518
rect 488382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 523826 704518
rect 524062 704282 524146 704518
rect 524382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 559826 704518
rect 560062 704282 560146 704518
rect 560382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -2966 696454 586890 696486
rect -2966 696218 -2934 696454
rect -2698 696218 -2614 696454
rect -2378 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 28826 696454
rect 29062 696218 29146 696454
rect 29382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 64826 696454
rect 65062 696218 65146 696454
rect 65382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 100826 696454
rect 101062 696218 101146 696454
rect 101382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 136826 696454
rect 137062 696218 137146 696454
rect 137382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 172826 696454
rect 173062 696218 173146 696454
rect 173382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 208826 696454
rect 209062 696218 209146 696454
rect 209382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 244826 696454
rect 245062 696218 245146 696454
rect 245382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 280826 696454
rect 281062 696218 281146 696454
rect 281382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 316826 696454
rect 317062 696218 317146 696454
rect 317382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 352826 696454
rect 353062 696218 353146 696454
rect 353382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 388826 696454
rect 389062 696218 389146 696454
rect 389382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 424826 696454
rect 425062 696218 425146 696454
rect 425382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 460826 696454
rect 461062 696218 461146 696454
rect 461382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 496826 696454
rect 497062 696218 497146 696454
rect 497382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 532826 696454
rect 533062 696218 533146 696454
rect 533382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 568826 696454
rect 569062 696218 569146 696454
rect 569382 696218 586302 696454
rect 586538 696218 586622 696454
rect 586858 696218 586890 696454
rect -2966 696134 586890 696218
rect -2966 695898 -2934 696134
rect -2698 695898 -2614 696134
rect -2378 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 28826 696134
rect 29062 695898 29146 696134
rect 29382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 64826 696134
rect 65062 695898 65146 696134
rect 65382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 100826 696134
rect 101062 695898 101146 696134
rect 101382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 136826 696134
rect 137062 695898 137146 696134
rect 137382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 172826 696134
rect 173062 695898 173146 696134
rect 173382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 208826 696134
rect 209062 695898 209146 696134
rect 209382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 244826 696134
rect 245062 695898 245146 696134
rect 245382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 280826 696134
rect 281062 695898 281146 696134
rect 281382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 316826 696134
rect 317062 695898 317146 696134
rect 317382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 352826 696134
rect 353062 695898 353146 696134
rect 353382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 388826 696134
rect 389062 695898 389146 696134
rect 389382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 424826 696134
rect 425062 695898 425146 696134
rect 425382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 460826 696134
rect 461062 695898 461146 696134
rect 461382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 496826 696134
rect 497062 695898 497146 696134
rect 497382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 532826 696134
rect 533062 695898 533146 696134
rect 533382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 568826 696134
rect 569062 695898 569146 696134
rect 569382 695898 586302 696134
rect 586538 695898 586622 696134
rect 586858 695898 586890 696134
rect -2966 695866 586890 695898
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 19826 687454
rect 20062 687218 20146 687454
rect 20382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 55826 687454
rect 56062 687218 56146 687454
rect 56382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 91826 687454
rect 92062 687218 92146 687454
rect 92382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 127826 687454
rect 128062 687218 128146 687454
rect 128382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 163826 687454
rect 164062 687218 164146 687454
rect 164382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 199826 687454
rect 200062 687218 200146 687454
rect 200382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 235826 687454
rect 236062 687218 236146 687454
rect 236382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 271826 687454
rect 272062 687218 272146 687454
rect 272382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 307826 687454
rect 308062 687218 308146 687454
rect 308382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 343826 687454
rect 344062 687218 344146 687454
rect 344382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 379826 687454
rect 380062 687218 380146 687454
rect 380382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 415826 687454
rect 416062 687218 416146 687454
rect 416382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 451826 687454
rect 452062 687218 452146 687454
rect 452382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 487826 687454
rect 488062 687218 488146 687454
rect 488382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 523826 687454
rect 524062 687218 524146 687454
rect 524382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 559826 687454
rect 560062 687218 560146 687454
rect 560382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 19826 687134
rect 20062 686898 20146 687134
rect 20382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 55826 687134
rect 56062 686898 56146 687134
rect 56382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 91826 687134
rect 92062 686898 92146 687134
rect 92382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 127826 687134
rect 128062 686898 128146 687134
rect 128382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 163826 687134
rect 164062 686898 164146 687134
rect 164382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 199826 687134
rect 200062 686898 200146 687134
rect 200382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 235826 687134
rect 236062 686898 236146 687134
rect 236382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 271826 687134
rect 272062 686898 272146 687134
rect 272382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 307826 687134
rect 308062 686898 308146 687134
rect 308382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 343826 687134
rect 344062 686898 344146 687134
rect 344382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 379826 687134
rect 380062 686898 380146 687134
rect 380382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 415826 687134
rect 416062 686898 416146 687134
rect 416382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 451826 687134
rect 452062 686898 452146 687134
rect 452382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 487826 687134
rect 488062 686898 488146 687134
rect 488382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 523826 687134
rect 524062 686898 524146 687134
rect 524382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 559826 687134
rect 560062 686898 560146 687134
rect 560382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -2966 678454 586890 678486
rect -2966 678218 -2934 678454
rect -2698 678218 -2614 678454
rect -2378 678218 10826 678454
rect 11062 678218 11146 678454
rect 11382 678218 22916 678454
rect 23152 678218 28847 678454
rect 29083 678218 49916 678454
rect 50152 678218 55847 678454
rect 56083 678218 76916 678454
rect 77152 678218 82847 678454
rect 83083 678218 103916 678454
rect 104152 678218 109847 678454
rect 110083 678218 130916 678454
rect 131152 678218 136847 678454
rect 137083 678218 157916 678454
rect 158152 678218 163847 678454
rect 164083 678218 184916 678454
rect 185152 678218 190847 678454
rect 191083 678218 211916 678454
rect 212152 678218 217847 678454
rect 218083 678218 238916 678454
rect 239152 678218 244847 678454
rect 245083 678218 265916 678454
rect 266152 678218 271847 678454
rect 272083 678218 292916 678454
rect 293152 678218 298847 678454
rect 299083 678218 319916 678454
rect 320152 678218 325847 678454
rect 326083 678218 346916 678454
rect 347152 678218 352847 678454
rect 353083 678218 373916 678454
rect 374152 678218 379847 678454
rect 380083 678218 400916 678454
rect 401152 678218 406847 678454
rect 407083 678218 427916 678454
rect 428152 678218 433847 678454
rect 434083 678218 454916 678454
rect 455152 678218 460847 678454
rect 461083 678218 481916 678454
rect 482152 678218 487847 678454
rect 488083 678218 508916 678454
rect 509152 678218 514847 678454
rect 515083 678218 535916 678454
rect 536152 678218 541847 678454
rect 542083 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 586302 678454
rect 586538 678218 586622 678454
rect 586858 678218 586890 678454
rect -2966 678134 586890 678218
rect -2966 677898 -2934 678134
rect -2698 677898 -2614 678134
rect -2378 677898 10826 678134
rect 11062 677898 11146 678134
rect 11382 677898 22916 678134
rect 23152 677898 28847 678134
rect 29083 677898 49916 678134
rect 50152 677898 55847 678134
rect 56083 677898 76916 678134
rect 77152 677898 82847 678134
rect 83083 677898 103916 678134
rect 104152 677898 109847 678134
rect 110083 677898 130916 678134
rect 131152 677898 136847 678134
rect 137083 677898 157916 678134
rect 158152 677898 163847 678134
rect 164083 677898 184916 678134
rect 185152 677898 190847 678134
rect 191083 677898 211916 678134
rect 212152 677898 217847 678134
rect 218083 677898 238916 678134
rect 239152 677898 244847 678134
rect 245083 677898 265916 678134
rect 266152 677898 271847 678134
rect 272083 677898 292916 678134
rect 293152 677898 298847 678134
rect 299083 677898 319916 678134
rect 320152 677898 325847 678134
rect 326083 677898 346916 678134
rect 347152 677898 352847 678134
rect 353083 677898 373916 678134
rect 374152 677898 379847 678134
rect 380083 677898 400916 678134
rect 401152 677898 406847 678134
rect 407083 677898 427916 678134
rect 428152 677898 433847 678134
rect 434083 677898 454916 678134
rect 455152 677898 460847 678134
rect 461083 677898 481916 678134
rect 482152 677898 487847 678134
rect 488083 677898 508916 678134
rect 509152 677898 514847 678134
rect 515083 677898 535916 678134
rect 536152 677898 541847 678134
rect 542083 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 586302 678134
rect 586538 677898 586622 678134
rect 586858 677898 586890 678134
rect -2966 677866 586890 677898
rect -2966 669454 586890 669486
rect -2966 669218 -1974 669454
rect -1738 669218 -1654 669454
rect -1418 669218 1826 669454
rect 2062 669218 2146 669454
rect 2382 669218 19952 669454
rect 20188 669218 25882 669454
rect 26118 669218 31813 669454
rect 32049 669218 46952 669454
rect 47188 669218 52882 669454
rect 53118 669218 58813 669454
rect 59049 669218 73952 669454
rect 74188 669218 79882 669454
rect 80118 669218 85813 669454
rect 86049 669218 100952 669454
rect 101188 669218 106882 669454
rect 107118 669218 112813 669454
rect 113049 669218 127952 669454
rect 128188 669218 133882 669454
rect 134118 669218 139813 669454
rect 140049 669218 154952 669454
rect 155188 669218 160882 669454
rect 161118 669218 166813 669454
rect 167049 669218 181952 669454
rect 182188 669218 187882 669454
rect 188118 669218 193813 669454
rect 194049 669218 208952 669454
rect 209188 669218 214882 669454
rect 215118 669218 220813 669454
rect 221049 669218 235952 669454
rect 236188 669218 241882 669454
rect 242118 669218 247813 669454
rect 248049 669218 262952 669454
rect 263188 669218 268882 669454
rect 269118 669218 274813 669454
rect 275049 669218 289952 669454
rect 290188 669218 295882 669454
rect 296118 669218 301813 669454
rect 302049 669218 316952 669454
rect 317188 669218 322882 669454
rect 323118 669218 328813 669454
rect 329049 669218 343952 669454
rect 344188 669218 349882 669454
rect 350118 669218 355813 669454
rect 356049 669218 370952 669454
rect 371188 669218 376882 669454
rect 377118 669218 382813 669454
rect 383049 669218 397952 669454
rect 398188 669218 403882 669454
rect 404118 669218 409813 669454
rect 410049 669218 424952 669454
rect 425188 669218 430882 669454
rect 431118 669218 436813 669454
rect 437049 669218 451952 669454
rect 452188 669218 457882 669454
rect 458118 669218 463813 669454
rect 464049 669218 478952 669454
rect 479188 669218 484882 669454
rect 485118 669218 490813 669454
rect 491049 669218 505952 669454
rect 506188 669218 511882 669454
rect 512118 669218 517813 669454
rect 518049 669218 532952 669454
rect 533188 669218 538882 669454
rect 539118 669218 544813 669454
rect 545049 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 577826 669454
rect 578062 669218 578146 669454
rect 578382 669218 585342 669454
rect 585578 669218 585662 669454
rect 585898 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -1974 669134
rect -1738 668898 -1654 669134
rect -1418 668898 1826 669134
rect 2062 668898 2146 669134
rect 2382 668898 19952 669134
rect 20188 668898 25882 669134
rect 26118 668898 31813 669134
rect 32049 668898 46952 669134
rect 47188 668898 52882 669134
rect 53118 668898 58813 669134
rect 59049 668898 73952 669134
rect 74188 668898 79882 669134
rect 80118 668898 85813 669134
rect 86049 668898 100952 669134
rect 101188 668898 106882 669134
rect 107118 668898 112813 669134
rect 113049 668898 127952 669134
rect 128188 668898 133882 669134
rect 134118 668898 139813 669134
rect 140049 668898 154952 669134
rect 155188 668898 160882 669134
rect 161118 668898 166813 669134
rect 167049 668898 181952 669134
rect 182188 668898 187882 669134
rect 188118 668898 193813 669134
rect 194049 668898 208952 669134
rect 209188 668898 214882 669134
rect 215118 668898 220813 669134
rect 221049 668898 235952 669134
rect 236188 668898 241882 669134
rect 242118 668898 247813 669134
rect 248049 668898 262952 669134
rect 263188 668898 268882 669134
rect 269118 668898 274813 669134
rect 275049 668898 289952 669134
rect 290188 668898 295882 669134
rect 296118 668898 301813 669134
rect 302049 668898 316952 669134
rect 317188 668898 322882 669134
rect 323118 668898 328813 669134
rect 329049 668898 343952 669134
rect 344188 668898 349882 669134
rect 350118 668898 355813 669134
rect 356049 668898 370952 669134
rect 371188 668898 376882 669134
rect 377118 668898 382813 669134
rect 383049 668898 397952 669134
rect 398188 668898 403882 669134
rect 404118 668898 409813 669134
rect 410049 668898 424952 669134
rect 425188 668898 430882 669134
rect 431118 668898 436813 669134
rect 437049 668898 451952 669134
rect 452188 668898 457882 669134
rect 458118 668898 463813 669134
rect 464049 668898 478952 669134
rect 479188 668898 484882 669134
rect 485118 668898 490813 669134
rect 491049 668898 505952 669134
rect 506188 668898 511882 669134
rect 512118 668898 517813 669134
rect 518049 668898 532952 669134
rect 533188 668898 538882 669134
rect 539118 668898 544813 669134
rect 545049 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 577826 669134
rect 578062 668898 578146 669134
rect 578382 668898 585342 669134
rect 585578 668898 585662 669134
rect 585898 668898 586890 669134
rect -2966 668866 586890 668898
rect 19794 661394 542414 661426
rect 19794 661158 19826 661394
rect 20062 661158 20146 661394
rect 20382 661158 37826 661394
rect 38062 661158 38146 661394
rect 38382 661158 55826 661394
rect 56062 661158 56146 661394
rect 56382 661158 73826 661394
rect 74062 661158 74146 661394
rect 74382 661158 91826 661394
rect 92062 661158 92146 661394
rect 92382 661158 109826 661394
rect 110062 661158 110146 661394
rect 110382 661158 127826 661394
rect 128062 661158 128146 661394
rect 128382 661158 145826 661394
rect 146062 661158 146146 661394
rect 146382 661158 163826 661394
rect 164062 661158 164146 661394
rect 164382 661158 181826 661394
rect 182062 661158 182146 661394
rect 182382 661158 199826 661394
rect 200062 661158 200146 661394
rect 200382 661158 217826 661394
rect 218062 661158 218146 661394
rect 218382 661158 235826 661394
rect 236062 661158 236146 661394
rect 236382 661158 253826 661394
rect 254062 661158 254146 661394
rect 254382 661158 271826 661394
rect 272062 661158 272146 661394
rect 272382 661158 289826 661394
rect 290062 661158 290146 661394
rect 290382 661158 307826 661394
rect 308062 661158 308146 661394
rect 308382 661158 325826 661394
rect 326062 661158 326146 661394
rect 326382 661158 343826 661394
rect 344062 661158 344146 661394
rect 344382 661158 361826 661394
rect 362062 661158 362146 661394
rect 362382 661158 379826 661394
rect 380062 661158 380146 661394
rect 380382 661158 397826 661394
rect 398062 661158 398146 661394
rect 398382 661158 415826 661394
rect 416062 661158 416146 661394
rect 416382 661158 433826 661394
rect 434062 661158 434146 661394
rect 434382 661158 451826 661394
rect 452062 661158 452146 661394
rect 452382 661158 469826 661394
rect 470062 661158 470146 661394
rect 470382 661158 487826 661394
rect 488062 661158 488146 661394
rect 488382 661158 505826 661394
rect 506062 661158 506146 661394
rect 506382 661158 523826 661394
rect 524062 661158 524146 661394
rect 524382 661158 541826 661394
rect 542062 661158 542146 661394
rect 542382 661158 542414 661394
rect 19794 661074 542414 661158
rect 19794 660838 19826 661074
rect 20062 660838 20146 661074
rect 20382 660838 37826 661074
rect 38062 660838 38146 661074
rect 38382 660838 55826 661074
rect 56062 660838 56146 661074
rect 56382 660838 73826 661074
rect 74062 660838 74146 661074
rect 74382 660838 91826 661074
rect 92062 660838 92146 661074
rect 92382 660838 109826 661074
rect 110062 660838 110146 661074
rect 110382 660838 127826 661074
rect 128062 660838 128146 661074
rect 128382 660838 145826 661074
rect 146062 660838 146146 661074
rect 146382 660838 163826 661074
rect 164062 660838 164146 661074
rect 164382 660838 181826 661074
rect 182062 660838 182146 661074
rect 182382 660838 199826 661074
rect 200062 660838 200146 661074
rect 200382 660838 217826 661074
rect 218062 660838 218146 661074
rect 218382 660838 235826 661074
rect 236062 660838 236146 661074
rect 236382 660838 253826 661074
rect 254062 660838 254146 661074
rect 254382 660838 271826 661074
rect 272062 660838 272146 661074
rect 272382 660838 289826 661074
rect 290062 660838 290146 661074
rect 290382 660838 307826 661074
rect 308062 660838 308146 661074
rect 308382 660838 325826 661074
rect 326062 660838 326146 661074
rect 326382 660838 343826 661074
rect 344062 660838 344146 661074
rect 344382 660838 361826 661074
rect 362062 660838 362146 661074
rect 362382 660838 379826 661074
rect 380062 660838 380146 661074
rect 380382 660838 397826 661074
rect 398062 660838 398146 661074
rect 398382 660838 415826 661074
rect 416062 660838 416146 661074
rect 416382 660838 433826 661074
rect 434062 660838 434146 661074
rect 434382 660838 451826 661074
rect 452062 660838 452146 661074
rect 452382 660838 469826 661074
rect 470062 660838 470146 661074
rect 470382 660838 487826 661074
rect 488062 660838 488146 661074
rect 488382 660838 505826 661074
rect 506062 660838 506146 661074
rect 506382 660838 523826 661074
rect 524062 660838 524146 661074
rect 524382 660838 541826 661074
rect 542062 660838 542146 661074
rect 542382 660838 542414 661074
rect 19794 660806 542414 660838
rect -2966 660454 586890 660486
rect -2966 660218 -2934 660454
rect -2698 660218 -2614 660454
rect -2378 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 28826 660454
rect 29062 660218 29146 660454
rect 29382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 64826 660454
rect 65062 660218 65146 660454
rect 65382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 100826 660454
rect 101062 660218 101146 660454
rect 101382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 136826 660454
rect 137062 660218 137146 660454
rect 137382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 172826 660454
rect 173062 660218 173146 660454
rect 173382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 208826 660454
rect 209062 660218 209146 660454
rect 209382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 244826 660454
rect 245062 660218 245146 660454
rect 245382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 280826 660454
rect 281062 660218 281146 660454
rect 281382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 316826 660454
rect 317062 660218 317146 660454
rect 317382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 352826 660454
rect 353062 660218 353146 660454
rect 353382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 388826 660454
rect 389062 660218 389146 660454
rect 389382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 424826 660454
rect 425062 660218 425146 660454
rect 425382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 460826 660454
rect 461062 660218 461146 660454
rect 461382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 496826 660454
rect 497062 660218 497146 660454
rect 497382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 532826 660454
rect 533062 660218 533146 660454
rect 533382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 568826 660454
rect 569062 660218 569146 660454
rect 569382 660218 586302 660454
rect 586538 660218 586622 660454
rect 586858 660218 586890 660454
rect -2966 660134 586890 660218
rect -2966 659898 -2934 660134
rect -2698 659898 -2614 660134
rect -2378 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 28826 660134
rect 29062 659898 29146 660134
rect 29382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 64826 660134
rect 65062 659898 65146 660134
rect 65382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 100826 660134
rect 101062 659898 101146 660134
rect 101382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 136826 660134
rect 137062 659898 137146 660134
rect 137382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 172826 660134
rect 173062 659898 173146 660134
rect 173382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 208826 660134
rect 209062 659898 209146 660134
rect 209382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 244826 660134
rect 245062 659898 245146 660134
rect 245382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 280826 660134
rect 281062 659898 281146 660134
rect 281382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 316826 660134
rect 317062 659898 317146 660134
rect 317382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 352826 660134
rect 353062 659898 353146 660134
rect 353382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 388826 660134
rect 389062 659898 389146 660134
rect 389382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 424826 660134
rect 425062 659898 425146 660134
rect 425382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 460826 660134
rect 461062 659898 461146 660134
rect 461382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 496826 660134
rect 497062 659898 497146 660134
rect 497382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 532826 660134
rect 533062 659898 533146 660134
rect 533382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 568826 660134
rect 569062 659898 569146 660134
rect 569382 659898 586302 660134
rect 586538 659898 586622 660134
rect 586858 659898 586890 660134
rect -2966 659866 586890 659898
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 19952 651454
rect 20188 651218 25882 651454
rect 26118 651218 31813 651454
rect 32049 651218 46952 651454
rect 47188 651218 52882 651454
rect 53118 651218 58813 651454
rect 59049 651218 73952 651454
rect 74188 651218 79882 651454
rect 80118 651218 85813 651454
rect 86049 651218 100952 651454
rect 101188 651218 106882 651454
rect 107118 651218 112813 651454
rect 113049 651218 127952 651454
rect 128188 651218 133882 651454
rect 134118 651218 139813 651454
rect 140049 651218 154952 651454
rect 155188 651218 160882 651454
rect 161118 651218 166813 651454
rect 167049 651218 181952 651454
rect 182188 651218 187882 651454
rect 188118 651218 193813 651454
rect 194049 651218 208952 651454
rect 209188 651218 214882 651454
rect 215118 651218 220813 651454
rect 221049 651218 235952 651454
rect 236188 651218 241882 651454
rect 242118 651218 247813 651454
rect 248049 651218 262952 651454
rect 263188 651218 268882 651454
rect 269118 651218 274813 651454
rect 275049 651218 289952 651454
rect 290188 651218 295882 651454
rect 296118 651218 301813 651454
rect 302049 651218 316952 651454
rect 317188 651218 322882 651454
rect 323118 651218 328813 651454
rect 329049 651218 343952 651454
rect 344188 651218 349882 651454
rect 350118 651218 355813 651454
rect 356049 651218 370952 651454
rect 371188 651218 376882 651454
rect 377118 651218 382813 651454
rect 383049 651218 397952 651454
rect 398188 651218 403882 651454
rect 404118 651218 409813 651454
rect 410049 651218 424952 651454
rect 425188 651218 430882 651454
rect 431118 651218 436813 651454
rect 437049 651218 451952 651454
rect 452188 651218 457882 651454
rect 458118 651218 463813 651454
rect 464049 651218 478952 651454
rect 479188 651218 484882 651454
rect 485118 651218 490813 651454
rect 491049 651218 505952 651454
rect 506188 651218 511882 651454
rect 512118 651218 517813 651454
rect 518049 651218 532952 651454
rect 533188 651218 538882 651454
rect 539118 651218 544813 651454
rect 545049 651218 559826 651454
rect 560062 651218 560146 651454
rect 560382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 19952 651134
rect 20188 650898 25882 651134
rect 26118 650898 31813 651134
rect 32049 650898 46952 651134
rect 47188 650898 52882 651134
rect 53118 650898 58813 651134
rect 59049 650898 73952 651134
rect 74188 650898 79882 651134
rect 80118 650898 85813 651134
rect 86049 650898 100952 651134
rect 101188 650898 106882 651134
rect 107118 650898 112813 651134
rect 113049 650898 127952 651134
rect 128188 650898 133882 651134
rect 134118 650898 139813 651134
rect 140049 650898 154952 651134
rect 155188 650898 160882 651134
rect 161118 650898 166813 651134
rect 167049 650898 181952 651134
rect 182188 650898 187882 651134
rect 188118 650898 193813 651134
rect 194049 650898 208952 651134
rect 209188 650898 214882 651134
rect 215118 650898 220813 651134
rect 221049 650898 235952 651134
rect 236188 650898 241882 651134
rect 242118 650898 247813 651134
rect 248049 650898 262952 651134
rect 263188 650898 268882 651134
rect 269118 650898 274813 651134
rect 275049 650898 289952 651134
rect 290188 650898 295882 651134
rect 296118 650898 301813 651134
rect 302049 650898 316952 651134
rect 317188 650898 322882 651134
rect 323118 650898 328813 651134
rect 329049 650898 343952 651134
rect 344188 650898 349882 651134
rect 350118 650898 355813 651134
rect 356049 650898 370952 651134
rect 371188 650898 376882 651134
rect 377118 650898 382813 651134
rect 383049 650898 397952 651134
rect 398188 650898 403882 651134
rect 404118 650898 409813 651134
rect 410049 650898 424952 651134
rect 425188 650898 430882 651134
rect 431118 650898 436813 651134
rect 437049 650898 451952 651134
rect 452188 650898 457882 651134
rect 458118 650898 463813 651134
rect 464049 650898 478952 651134
rect 479188 650898 484882 651134
rect 485118 650898 490813 651134
rect 491049 650898 505952 651134
rect 506188 650898 511882 651134
rect 512118 650898 517813 651134
rect 518049 650898 532952 651134
rect 533188 650898 538882 651134
rect 539118 650898 544813 651134
rect 545049 650898 559826 651134
rect 560062 650898 560146 651134
rect 560382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -2966 642454 586890 642486
rect -2966 642218 -2934 642454
rect -2698 642218 -2614 642454
rect -2378 642218 10826 642454
rect 11062 642218 11146 642454
rect 11382 642218 22916 642454
rect 23152 642218 28847 642454
rect 29083 642218 49916 642454
rect 50152 642218 55847 642454
rect 56083 642218 76916 642454
rect 77152 642218 82847 642454
rect 83083 642218 103916 642454
rect 104152 642218 109847 642454
rect 110083 642218 130916 642454
rect 131152 642218 136847 642454
rect 137083 642218 157916 642454
rect 158152 642218 163847 642454
rect 164083 642218 184916 642454
rect 185152 642218 190847 642454
rect 191083 642218 211916 642454
rect 212152 642218 217847 642454
rect 218083 642218 238916 642454
rect 239152 642218 244847 642454
rect 245083 642218 265916 642454
rect 266152 642218 271847 642454
rect 272083 642218 292916 642454
rect 293152 642218 298847 642454
rect 299083 642218 319916 642454
rect 320152 642218 325847 642454
rect 326083 642218 346916 642454
rect 347152 642218 352847 642454
rect 353083 642218 373916 642454
rect 374152 642218 379847 642454
rect 380083 642218 400916 642454
rect 401152 642218 406847 642454
rect 407083 642218 427916 642454
rect 428152 642218 433847 642454
rect 434083 642218 454916 642454
rect 455152 642218 460847 642454
rect 461083 642218 481916 642454
rect 482152 642218 487847 642454
rect 488083 642218 508916 642454
rect 509152 642218 514847 642454
rect 515083 642218 535916 642454
rect 536152 642218 541847 642454
rect 542083 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 586302 642454
rect 586538 642218 586622 642454
rect 586858 642218 586890 642454
rect -2966 642134 586890 642218
rect -2966 641898 -2934 642134
rect -2698 641898 -2614 642134
rect -2378 641898 10826 642134
rect 11062 641898 11146 642134
rect 11382 641898 22916 642134
rect 23152 641898 28847 642134
rect 29083 641898 49916 642134
rect 50152 641898 55847 642134
rect 56083 641898 76916 642134
rect 77152 641898 82847 642134
rect 83083 641898 103916 642134
rect 104152 641898 109847 642134
rect 110083 641898 130916 642134
rect 131152 641898 136847 642134
rect 137083 641898 157916 642134
rect 158152 641898 163847 642134
rect 164083 641898 184916 642134
rect 185152 641898 190847 642134
rect 191083 641898 211916 642134
rect 212152 641898 217847 642134
rect 218083 641898 238916 642134
rect 239152 641898 244847 642134
rect 245083 641898 265916 642134
rect 266152 641898 271847 642134
rect 272083 641898 292916 642134
rect 293152 641898 298847 642134
rect 299083 641898 319916 642134
rect 320152 641898 325847 642134
rect 326083 641898 346916 642134
rect 347152 641898 352847 642134
rect 353083 641898 373916 642134
rect 374152 641898 379847 642134
rect 380083 641898 400916 642134
rect 401152 641898 406847 642134
rect 407083 641898 427916 642134
rect 428152 641898 433847 642134
rect 434083 641898 454916 642134
rect 455152 641898 460847 642134
rect 461083 641898 481916 642134
rect 482152 641898 487847 642134
rect 488083 641898 508916 642134
rect 509152 641898 514847 642134
rect 515083 641898 535916 642134
rect 536152 641898 541847 642134
rect 542083 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 586302 642134
rect 586538 641898 586622 642134
rect 586858 641898 586890 642134
rect -2966 641866 586890 641898
rect 28794 634394 551414 634426
rect 28794 634158 28826 634394
rect 29062 634158 29146 634394
rect 29382 634158 46826 634394
rect 47062 634158 47146 634394
rect 47382 634158 64826 634394
rect 65062 634158 65146 634394
rect 65382 634158 82826 634394
rect 83062 634158 83146 634394
rect 83382 634158 100826 634394
rect 101062 634158 101146 634394
rect 101382 634158 118826 634394
rect 119062 634158 119146 634394
rect 119382 634158 136826 634394
rect 137062 634158 137146 634394
rect 137382 634158 154826 634394
rect 155062 634158 155146 634394
rect 155382 634158 172826 634394
rect 173062 634158 173146 634394
rect 173382 634158 190826 634394
rect 191062 634158 191146 634394
rect 191382 634158 208826 634394
rect 209062 634158 209146 634394
rect 209382 634158 226826 634394
rect 227062 634158 227146 634394
rect 227382 634158 244826 634394
rect 245062 634158 245146 634394
rect 245382 634158 262826 634394
rect 263062 634158 263146 634394
rect 263382 634158 280826 634394
rect 281062 634158 281146 634394
rect 281382 634158 298826 634394
rect 299062 634158 299146 634394
rect 299382 634158 316826 634394
rect 317062 634158 317146 634394
rect 317382 634158 334826 634394
rect 335062 634158 335146 634394
rect 335382 634158 352826 634394
rect 353062 634158 353146 634394
rect 353382 634158 370826 634394
rect 371062 634158 371146 634394
rect 371382 634158 388826 634394
rect 389062 634158 389146 634394
rect 389382 634158 406826 634394
rect 407062 634158 407146 634394
rect 407382 634158 424826 634394
rect 425062 634158 425146 634394
rect 425382 634158 442826 634394
rect 443062 634158 443146 634394
rect 443382 634158 460826 634394
rect 461062 634158 461146 634394
rect 461382 634158 478826 634394
rect 479062 634158 479146 634394
rect 479382 634158 496826 634394
rect 497062 634158 497146 634394
rect 497382 634158 514826 634394
rect 515062 634158 515146 634394
rect 515382 634158 532826 634394
rect 533062 634158 533146 634394
rect 533382 634158 550826 634394
rect 551062 634158 551146 634394
rect 551382 634158 551414 634394
rect 28794 634074 551414 634158
rect 28794 633838 28826 634074
rect 29062 633838 29146 634074
rect 29382 633838 46826 634074
rect 47062 633838 47146 634074
rect 47382 633838 64826 634074
rect 65062 633838 65146 634074
rect 65382 633838 82826 634074
rect 83062 633838 83146 634074
rect 83382 633838 100826 634074
rect 101062 633838 101146 634074
rect 101382 633838 118826 634074
rect 119062 633838 119146 634074
rect 119382 633838 136826 634074
rect 137062 633838 137146 634074
rect 137382 633838 154826 634074
rect 155062 633838 155146 634074
rect 155382 633838 172826 634074
rect 173062 633838 173146 634074
rect 173382 633838 190826 634074
rect 191062 633838 191146 634074
rect 191382 633838 208826 634074
rect 209062 633838 209146 634074
rect 209382 633838 226826 634074
rect 227062 633838 227146 634074
rect 227382 633838 244826 634074
rect 245062 633838 245146 634074
rect 245382 633838 262826 634074
rect 263062 633838 263146 634074
rect 263382 633838 280826 634074
rect 281062 633838 281146 634074
rect 281382 633838 298826 634074
rect 299062 633838 299146 634074
rect 299382 633838 316826 634074
rect 317062 633838 317146 634074
rect 317382 633838 334826 634074
rect 335062 633838 335146 634074
rect 335382 633838 352826 634074
rect 353062 633838 353146 634074
rect 353382 633838 370826 634074
rect 371062 633838 371146 634074
rect 371382 633838 388826 634074
rect 389062 633838 389146 634074
rect 389382 633838 406826 634074
rect 407062 633838 407146 634074
rect 407382 633838 424826 634074
rect 425062 633838 425146 634074
rect 425382 633838 442826 634074
rect 443062 633838 443146 634074
rect 443382 633838 460826 634074
rect 461062 633838 461146 634074
rect 461382 633838 478826 634074
rect 479062 633838 479146 634074
rect 479382 633838 496826 634074
rect 497062 633838 497146 634074
rect 497382 633838 514826 634074
rect 515062 633838 515146 634074
rect 515382 633838 532826 634074
rect 533062 633838 533146 634074
rect 533382 633838 550826 634074
rect 551062 633838 551146 634074
rect 551382 633838 551414 634074
rect 28794 633806 551414 633838
rect -2966 633454 586890 633486
rect -2966 633218 -1974 633454
rect -1738 633218 -1654 633454
rect -1418 633218 1826 633454
rect 2062 633218 2146 633454
rect 2382 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 37826 633454
rect 38062 633218 38146 633454
rect 38382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 73826 633454
rect 74062 633218 74146 633454
rect 74382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 109826 633454
rect 110062 633218 110146 633454
rect 110382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 145826 633454
rect 146062 633218 146146 633454
rect 146382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 181826 633454
rect 182062 633218 182146 633454
rect 182382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 217826 633454
rect 218062 633218 218146 633454
rect 218382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 253826 633454
rect 254062 633218 254146 633454
rect 254382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 289826 633454
rect 290062 633218 290146 633454
rect 290382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 325826 633454
rect 326062 633218 326146 633454
rect 326382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 361826 633454
rect 362062 633218 362146 633454
rect 362382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 397826 633454
rect 398062 633218 398146 633454
rect 398382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 433826 633454
rect 434062 633218 434146 633454
rect 434382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 469826 633454
rect 470062 633218 470146 633454
rect 470382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 505826 633454
rect 506062 633218 506146 633454
rect 506382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 541826 633454
rect 542062 633218 542146 633454
rect 542382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 577826 633454
rect 578062 633218 578146 633454
rect 578382 633218 585342 633454
rect 585578 633218 585662 633454
rect 585898 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -1974 633134
rect -1738 632898 -1654 633134
rect -1418 632898 1826 633134
rect 2062 632898 2146 633134
rect 2382 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 37826 633134
rect 38062 632898 38146 633134
rect 38382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 73826 633134
rect 74062 632898 74146 633134
rect 74382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 109826 633134
rect 110062 632898 110146 633134
rect 110382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 145826 633134
rect 146062 632898 146146 633134
rect 146382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 181826 633134
rect 182062 632898 182146 633134
rect 182382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 217826 633134
rect 218062 632898 218146 633134
rect 218382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 253826 633134
rect 254062 632898 254146 633134
rect 254382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 289826 633134
rect 290062 632898 290146 633134
rect 290382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 325826 633134
rect 326062 632898 326146 633134
rect 326382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 361826 633134
rect 362062 632898 362146 633134
rect 362382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 397826 633134
rect 398062 632898 398146 633134
rect 398382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 433826 633134
rect 434062 632898 434146 633134
rect 434382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 469826 633134
rect 470062 632898 470146 633134
rect 470382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 505826 633134
rect 506062 632898 506146 633134
rect 506382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 541826 633134
rect 542062 632898 542146 633134
rect 542382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 577826 633134
rect 578062 632898 578146 633134
rect 578382 632898 585342 633134
rect 585578 632898 585662 633134
rect 585898 632898 586890 633134
rect -2966 632866 586890 632898
rect -2966 624454 586890 624486
rect -2966 624218 -2934 624454
rect -2698 624218 -2614 624454
rect -2378 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 22916 624454
rect 23152 624218 28847 624454
rect 29083 624218 49916 624454
rect 50152 624218 55847 624454
rect 56083 624218 76916 624454
rect 77152 624218 82847 624454
rect 83083 624218 103916 624454
rect 104152 624218 109847 624454
rect 110083 624218 130916 624454
rect 131152 624218 136847 624454
rect 137083 624218 157916 624454
rect 158152 624218 163847 624454
rect 164083 624218 184916 624454
rect 185152 624218 190847 624454
rect 191083 624218 211916 624454
rect 212152 624218 217847 624454
rect 218083 624218 238916 624454
rect 239152 624218 244847 624454
rect 245083 624218 265916 624454
rect 266152 624218 271847 624454
rect 272083 624218 292916 624454
rect 293152 624218 298847 624454
rect 299083 624218 319916 624454
rect 320152 624218 325847 624454
rect 326083 624218 346916 624454
rect 347152 624218 352847 624454
rect 353083 624218 373916 624454
rect 374152 624218 379847 624454
rect 380083 624218 400916 624454
rect 401152 624218 406847 624454
rect 407083 624218 427916 624454
rect 428152 624218 433847 624454
rect 434083 624218 454916 624454
rect 455152 624218 460847 624454
rect 461083 624218 481916 624454
rect 482152 624218 487847 624454
rect 488083 624218 508916 624454
rect 509152 624218 514847 624454
rect 515083 624218 535916 624454
rect 536152 624218 541847 624454
rect 542083 624218 568826 624454
rect 569062 624218 569146 624454
rect 569382 624218 586302 624454
rect 586538 624218 586622 624454
rect 586858 624218 586890 624454
rect -2966 624134 586890 624218
rect -2966 623898 -2934 624134
rect -2698 623898 -2614 624134
rect -2378 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 22916 624134
rect 23152 623898 28847 624134
rect 29083 623898 49916 624134
rect 50152 623898 55847 624134
rect 56083 623898 76916 624134
rect 77152 623898 82847 624134
rect 83083 623898 103916 624134
rect 104152 623898 109847 624134
rect 110083 623898 130916 624134
rect 131152 623898 136847 624134
rect 137083 623898 157916 624134
rect 158152 623898 163847 624134
rect 164083 623898 184916 624134
rect 185152 623898 190847 624134
rect 191083 623898 211916 624134
rect 212152 623898 217847 624134
rect 218083 623898 238916 624134
rect 239152 623898 244847 624134
rect 245083 623898 265916 624134
rect 266152 623898 271847 624134
rect 272083 623898 292916 624134
rect 293152 623898 298847 624134
rect 299083 623898 319916 624134
rect 320152 623898 325847 624134
rect 326083 623898 346916 624134
rect 347152 623898 352847 624134
rect 353083 623898 373916 624134
rect 374152 623898 379847 624134
rect 380083 623898 400916 624134
rect 401152 623898 406847 624134
rect 407083 623898 427916 624134
rect 428152 623898 433847 624134
rect 434083 623898 454916 624134
rect 455152 623898 460847 624134
rect 461083 623898 481916 624134
rect 482152 623898 487847 624134
rect 488083 623898 508916 624134
rect 509152 623898 514847 624134
rect 515083 623898 535916 624134
rect 536152 623898 541847 624134
rect 542083 623898 568826 624134
rect 569062 623898 569146 624134
rect 569382 623898 586302 624134
rect 586538 623898 586622 624134
rect 586858 623898 586890 624134
rect -2966 623866 586890 623898
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 19952 615454
rect 20188 615218 25882 615454
rect 26118 615218 31813 615454
rect 32049 615218 46952 615454
rect 47188 615218 52882 615454
rect 53118 615218 58813 615454
rect 59049 615218 73952 615454
rect 74188 615218 79882 615454
rect 80118 615218 85813 615454
rect 86049 615218 100952 615454
rect 101188 615218 106882 615454
rect 107118 615218 112813 615454
rect 113049 615218 127952 615454
rect 128188 615218 133882 615454
rect 134118 615218 139813 615454
rect 140049 615218 154952 615454
rect 155188 615218 160882 615454
rect 161118 615218 166813 615454
rect 167049 615218 181952 615454
rect 182188 615218 187882 615454
rect 188118 615218 193813 615454
rect 194049 615218 208952 615454
rect 209188 615218 214882 615454
rect 215118 615218 220813 615454
rect 221049 615218 235952 615454
rect 236188 615218 241882 615454
rect 242118 615218 247813 615454
rect 248049 615218 262952 615454
rect 263188 615218 268882 615454
rect 269118 615218 274813 615454
rect 275049 615218 289952 615454
rect 290188 615218 295882 615454
rect 296118 615218 301813 615454
rect 302049 615218 316952 615454
rect 317188 615218 322882 615454
rect 323118 615218 328813 615454
rect 329049 615218 343952 615454
rect 344188 615218 349882 615454
rect 350118 615218 355813 615454
rect 356049 615218 370952 615454
rect 371188 615218 376882 615454
rect 377118 615218 382813 615454
rect 383049 615218 397952 615454
rect 398188 615218 403882 615454
rect 404118 615218 409813 615454
rect 410049 615218 424952 615454
rect 425188 615218 430882 615454
rect 431118 615218 436813 615454
rect 437049 615218 451952 615454
rect 452188 615218 457882 615454
rect 458118 615218 463813 615454
rect 464049 615218 478952 615454
rect 479188 615218 484882 615454
rect 485118 615218 490813 615454
rect 491049 615218 505952 615454
rect 506188 615218 511882 615454
rect 512118 615218 517813 615454
rect 518049 615218 532952 615454
rect 533188 615218 538882 615454
rect 539118 615218 544813 615454
rect 545049 615218 559826 615454
rect 560062 615218 560146 615454
rect 560382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 19952 615134
rect 20188 614898 25882 615134
rect 26118 614898 31813 615134
rect 32049 614898 46952 615134
rect 47188 614898 52882 615134
rect 53118 614898 58813 615134
rect 59049 614898 73952 615134
rect 74188 614898 79882 615134
rect 80118 614898 85813 615134
rect 86049 614898 100952 615134
rect 101188 614898 106882 615134
rect 107118 614898 112813 615134
rect 113049 614898 127952 615134
rect 128188 614898 133882 615134
rect 134118 614898 139813 615134
rect 140049 614898 154952 615134
rect 155188 614898 160882 615134
rect 161118 614898 166813 615134
rect 167049 614898 181952 615134
rect 182188 614898 187882 615134
rect 188118 614898 193813 615134
rect 194049 614898 208952 615134
rect 209188 614898 214882 615134
rect 215118 614898 220813 615134
rect 221049 614898 235952 615134
rect 236188 614898 241882 615134
rect 242118 614898 247813 615134
rect 248049 614898 262952 615134
rect 263188 614898 268882 615134
rect 269118 614898 274813 615134
rect 275049 614898 289952 615134
rect 290188 614898 295882 615134
rect 296118 614898 301813 615134
rect 302049 614898 316952 615134
rect 317188 614898 322882 615134
rect 323118 614898 328813 615134
rect 329049 614898 343952 615134
rect 344188 614898 349882 615134
rect 350118 614898 355813 615134
rect 356049 614898 370952 615134
rect 371188 614898 376882 615134
rect 377118 614898 382813 615134
rect 383049 614898 397952 615134
rect 398188 614898 403882 615134
rect 404118 614898 409813 615134
rect 410049 614898 424952 615134
rect 425188 614898 430882 615134
rect 431118 614898 436813 615134
rect 437049 614898 451952 615134
rect 452188 614898 457882 615134
rect 458118 614898 463813 615134
rect 464049 614898 478952 615134
rect 479188 614898 484882 615134
rect 485118 614898 490813 615134
rect 491049 614898 505952 615134
rect 506188 614898 511882 615134
rect 512118 614898 517813 615134
rect 518049 614898 532952 615134
rect 533188 614898 538882 615134
rect 539118 614898 544813 615134
rect 545049 614898 559826 615134
rect 560062 614898 560146 615134
rect 560382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect 19794 607394 542414 607426
rect 19794 607158 19826 607394
rect 20062 607158 20146 607394
rect 20382 607158 37826 607394
rect 38062 607158 38146 607394
rect 38382 607158 55826 607394
rect 56062 607158 56146 607394
rect 56382 607158 73826 607394
rect 74062 607158 74146 607394
rect 74382 607158 91826 607394
rect 92062 607158 92146 607394
rect 92382 607158 109826 607394
rect 110062 607158 110146 607394
rect 110382 607158 127826 607394
rect 128062 607158 128146 607394
rect 128382 607158 145826 607394
rect 146062 607158 146146 607394
rect 146382 607158 163826 607394
rect 164062 607158 164146 607394
rect 164382 607158 181826 607394
rect 182062 607158 182146 607394
rect 182382 607158 199826 607394
rect 200062 607158 200146 607394
rect 200382 607158 217826 607394
rect 218062 607158 218146 607394
rect 218382 607158 235826 607394
rect 236062 607158 236146 607394
rect 236382 607158 253826 607394
rect 254062 607158 254146 607394
rect 254382 607158 271826 607394
rect 272062 607158 272146 607394
rect 272382 607158 289826 607394
rect 290062 607158 290146 607394
rect 290382 607158 307826 607394
rect 308062 607158 308146 607394
rect 308382 607158 325826 607394
rect 326062 607158 326146 607394
rect 326382 607158 343826 607394
rect 344062 607158 344146 607394
rect 344382 607158 361826 607394
rect 362062 607158 362146 607394
rect 362382 607158 379826 607394
rect 380062 607158 380146 607394
rect 380382 607158 397826 607394
rect 398062 607158 398146 607394
rect 398382 607158 415826 607394
rect 416062 607158 416146 607394
rect 416382 607158 433826 607394
rect 434062 607158 434146 607394
rect 434382 607158 451826 607394
rect 452062 607158 452146 607394
rect 452382 607158 469826 607394
rect 470062 607158 470146 607394
rect 470382 607158 487826 607394
rect 488062 607158 488146 607394
rect 488382 607158 505826 607394
rect 506062 607158 506146 607394
rect 506382 607158 523826 607394
rect 524062 607158 524146 607394
rect 524382 607158 541826 607394
rect 542062 607158 542146 607394
rect 542382 607158 542414 607394
rect 19794 607074 542414 607158
rect 19794 606838 19826 607074
rect 20062 606838 20146 607074
rect 20382 606838 37826 607074
rect 38062 606838 38146 607074
rect 38382 606838 55826 607074
rect 56062 606838 56146 607074
rect 56382 606838 73826 607074
rect 74062 606838 74146 607074
rect 74382 606838 91826 607074
rect 92062 606838 92146 607074
rect 92382 606838 109826 607074
rect 110062 606838 110146 607074
rect 110382 606838 127826 607074
rect 128062 606838 128146 607074
rect 128382 606838 145826 607074
rect 146062 606838 146146 607074
rect 146382 606838 163826 607074
rect 164062 606838 164146 607074
rect 164382 606838 181826 607074
rect 182062 606838 182146 607074
rect 182382 606838 199826 607074
rect 200062 606838 200146 607074
rect 200382 606838 217826 607074
rect 218062 606838 218146 607074
rect 218382 606838 235826 607074
rect 236062 606838 236146 607074
rect 236382 606838 253826 607074
rect 254062 606838 254146 607074
rect 254382 606838 271826 607074
rect 272062 606838 272146 607074
rect 272382 606838 289826 607074
rect 290062 606838 290146 607074
rect 290382 606838 307826 607074
rect 308062 606838 308146 607074
rect 308382 606838 325826 607074
rect 326062 606838 326146 607074
rect 326382 606838 343826 607074
rect 344062 606838 344146 607074
rect 344382 606838 361826 607074
rect 362062 606838 362146 607074
rect 362382 606838 379826 607074
rect 380062 606838 380146 607074
rect 380382 606838 397826 607074
rect 398062 606838 398146 607074
rect 398382 606838 415826 607074
rect 416062 606838 416146 607074
rect 416382 606838 433826 607074
rect 434062 606838 434146 607074
rect 434382 606838 451826 607074
rect 452062 606838 452146 607074
rect 452382 606838 469826 607074
rect 470062 606838 470146 607074
rect 470382 606838 487826 607074
rect 488062 606838 488146 607074
rect 488382 606838 505826 607074
rect 506062 606838 506146 607074
rect 506382 606838 523826 607074
rect 524062 606838 524146 607074
rect 524382 606838 541826 607074
rect 542062 606838 542146 607074
rect 542382 606838 542414 607074
rect 19794 606806 542414 606838
rect -2966 606454 586890 606486
rect -2966 606218 -2934 606454
rect -2698 606218 -2614 606454
rect -2378 606218 10826 606454
rect 11062 606218 11146 606454
rect 11382 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 46826 606454
rect 47062 606218 47146 606454
rect 47382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 82826 606454
rect 83062 606218 83146 606454
rect 83382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 118826 606454
rect 119062 606218 119146 606454
rect 119382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 154826 606454
rect 155062 606218 155146 606454
rect 155382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 190826 606454
rect 191062 606218 191146 606454
rect 191382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 226826 606454
rect 227062 606218 227146 606454
rect 227382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 262826 606454
rect 263062 606218 263146 606454
rect 263382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 298826 606454
rect 299062 606218 299146 606454
rect 299382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 334826 606454
rect 335062 606218 335146 606454
rect 335382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 370826 606454
rect 371062 606218 371146 606454
rect 371382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 406826 606454
rect 407062 606218 407146 606454
rect 407382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 442826 606454
rect 443062 606218 443146 606454
rect 443382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 478826 606454
rect 479062 606218 479146 606454
rect 479382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 514826 606454
rect 515062 606218 515146 606454
rect 515382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 550826 606454
rect 551062 606218 551146 606454
rect 551382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 586302 606454
rect 586538 606218 586622 606454
rect 586858 606218 586890 606454
rect -2966 606134 586890 606218
rect -2966 605898 -2934 606134
rect -2698 605898 -2614 606134
rect -2378 605898 10826 606134
rect 11062 605898 11146 606134
rect 11382 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 46826 606134
rect 47062 605898 47146 606134
rect 47382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 82826 606134
rect 83062 605898 83146 606134
rect 83382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 118826 606134
rect 119062 605898 119146 606134
rect 119382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 154826 606134
rect 155062 605898 155146 606134
rect 155382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 190826 606134
rect 191062 605898 191146 606134
rect 191382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 226826 606134
rect 227062 605898 227146 606134
rect 227382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 262826 606134
rect 263062 605898 263146 606134
rect 263382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 298826 606134
rect 299062 605898 299146 606134
rect 299382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 334826 606134
rect 335062 605898 335146 606134
rect 335382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 370826 606134
rect 371062 605898 371146 606134
rect 371382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 406826 606134
rect 407062 605898 407146 606134
rect 407382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 442826 606134
rect 443062 605898 443146 606134
rect 443382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 478826 606134
rect 479062 605898 479146 606134
rect 479382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 514826 606134
rect 515062 605898 515146 606134
rect 515382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 550826 606134
rect 551062 605898 551146 606134
rect 551382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 586302 606134
rect 586538 605898 586622 606134
rect 586858 605898 586890 606134
rect -2966 605866 586890 605898
rect -2966 597454 586890 597486
rect -2966 597218 -1974 597454
rect -1738 597218 -1654 597454
rect -1418 597218 1826 597454
rect 2062 597218 2146 597454
rect 2382 597218 19952 597454
rect 20188 597218 25882 597454
rect 26118 597218 31813 597454
rect 32049 597218 46952 597454
rect 47188 597218 52882 597454
rect 53118 597218 58813 597454
rect 59049 597218 73952 597454
rect 74188 597218 79882 597454
rect 80118 597218 85813 597454
rect 86049 597218 100952 597454
rect 101188 597218 106882 597454
rect 107118 597218 112813 597454
rect 113049 597218 127952 597454
rect 128188 597218 133882 597454
rect 134118 597218 139813 597454
rect 140049 597218 154952 597454
rect 155188 597218 160882 597454
rect 161118 597218 166813 597454
rect 167049 597218 181952 597454
rect 182188 597218 187882 597454
rect 188118 597218 193813 597454
rect 194049 597218 208952 597454
rect 209188 597218 214882 597454
rect 215118 597218 220813 597454
rect 221049 597218 235952 597454
rect 236188 597218 241882 597454
rect 242118 597218 247813 597454
rect 248049 597218 262952 597454
rect 263188 597218 268882 597454
rect 269118 597218 274813 597454
rect 275049 597218 289952 597454
rect 290188 597218 295882 597454
rect 296118 597218 301813 597454
rect 302049 597218 316952 597454
rect 317188 597218 322882 597454
rect 323118 597218 328813 597454
rect 329049 597218 343952 597454
rect 344188 597218 349882 597454
rect 350118 597218 355813 597454
rect 356049 597218 370952 597454
rect 371188 597218 376882 597454
rect 377118 597218 382813 597454
rect 383049 597218 397952 597454
rect 398188 597218 403882 597454
rect 404118 597218 409813 597454
rect 410049 597218 424952 597454
rect 425188 597218 430882 597454
rect 431118 597218 436813 597454
rect 437049 597218 451952 597454
rect 452188 597218 457882 597454
rect 458118 597218 463813 597454
rect 464049 597218 478952 597454
rect 479188 597218 484882 597454
rect 485118 597218 490813 597454
rect 491049 597218 505952 597454
rect 506188 597218 511882 597454
rect 512118 597218 517813 597454
rect 518049 597218 532952 597454
rect 533188 597218 538882 597454
rect 539118 597218 544813 597454
rect 545049 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 577826 597454
rect 578062 597218 578146 597454
rect 578382 597218 585342 597454
rect 585578 597218 585662 597454
rect 585898 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -1974 597134
rect -1738 596898 -1654 597134
rect -1418 596898 1826 597134
rect 2062 596898 2146 597134
rect 2382 596898 19952 597134
rect 20188 596898 25882 597134
rect 26118 596898 31813 597134
rect 32049 596898 46952 597134
rect 47188 596898 52882 597134
rect 53118 596898 58813 597134
rect 59049 596898 73952 597134
rect 74188 596898 79882 597134
rect 80118 596898 85813 597134
rect 86049 596898 100952 597134
rect 101188 596898 106882 597134
rect 107118 596898 112813 597134
rect 113049 596898 127952 597134
rect 128188 596898 133882 597134
rect 134118 596898 139813 597134
rect 140049 596898 154952 597134
rect 155188 596898 160882 597134
rect 161118 596898 166813 597134
rect 167049 596898 181952 597134
rect 182188 596898 187882 597134
rect 188118 596898 193813 597134
rect 194049 596898 208952 597134
rect 209188 596898 214882 597134
rect 215118 596898 220813 597134
rect 221049 596898 235952 597134
rect 236188 596898 241882 597134
rect 242118 596898 247813 597134
rect 248049 596898 262952 597134
rect 263188 596898 268882 597134
rect 269118 596898 274813 597134
rect 275049 596898 289952 597134
rect 290188 596898 295882 597134
rect 296118 596898 301813 597134
rect 302049 596898 316952 597134
rect 317188 596898 322882 597134
rect 323118 596898 328813 597134
rect 329049 596898 343952 597134
rect 344188 596898 349882 597134
rect 350118 596898 355813 597134
rect 356049 596898 370952 597134
rect 371188 596898 376882 597134
rect 377118 596898 382813 597134
rect 383049 596898 397952 597134
rect 398188 596898 403882 597134
rect 404118 596898 409813 597134
rect 410049 596898 424952 597134
rect 425188 596898 430882 597134
rect 431118 596898 436813 597134
rect 437049 596898 451952 597134
rect 452188 596898 457882 597134
rect 458118 596898 463813 597134
rect 464049 596898 478952 597134
rect 479188 596898 484882 597134
rect 485118 596898 490813 597134
rect 491049 596898 505952 597134
rect 506188 596898 511882 597134
rect 512118 596898 517813 597134
rect 518049 596898 532952 597134
rect 533188 596898 538882 597134
rect 539118 596898 544813 597134
rect 545049 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 577826 597134
rect 578062 596898 578146 597134
rect 578382 596898 585342 597134
rect 585578 596898 585662 597134
rect 585898 596898 586890 597134
rect -2966 596866 586890 596898
rect -2966 588454 586890 588486
rect -2966 588218 -2934 588454
rect -2698 588218 -2614 588454
rect -2378 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 22916 588454
rect 23152 588218 28847 588454
rect 29083 588218 49916 588454
rect 50152 588218 55847 588454
rect 56083 588218 76916 588454
rect 77152 588218 82847 588454
rect 83083 588218 103916 588454
rect 104152 588218 109847 588454
rect 110083 588218 130916 588454
rect 131152 588218 136847 588454
rect 137083 588218 157916 588454
rect 158152 588218 163847 588454
rect 164083 588218 184916 588454
rect 185152 588218 190847 588454
rect 191083 588218 211916 588454
rect 212152 588218 217847 588454
rect 218083 588218 238916 588454
rect 239152 588218 244847 588454
rect 245083 588218 265916 588454
rect 266152 588218 271847 588454
rect 272083 588218 292916 588454
rect 293152 588218 298847 588454
rect 299083 588218 319916 588454
rect 320152 588218 325847 588454
rect 326083 588218 346916 588454
rect 347152 588218 352847 588454
rect 353083 588218 373916 588454
rect 374152 588218 379847 588454
rect 380083 588218 400916 588454
rect 401152 588218 406847 588454
rect 407083 588218 427916 588454
rect 428152 588218 433847 588454
rect 434083 588218 454916 588454
rect 455152 588218 460847 588454
rect 461083 588218 481916 588454
rect 482152 588218 487847 588454
rect 488083 588218 508916 588454
rect 509152 588218 514847 588454
rect 515083 588218 535916 588454
rect 536152 588218 541847 588454
rect 542083 588218 568826 588454
rect 569062 588218 569146 588454
rect 569382 588218 586302 588454
rect 586538 588218 586622 588454
rect 586858 588218 586890 588454
rect -2966 588134 586890 588218
rect -2966 587898 -2934 588134
rect -2698 587898 -2614 588134
rect -2378 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 22916 588134
rect 23152 587898 28847 588134
rect 29083 587898 49916 588134
rect 50152 587898 55847 588134
rect 56083 587898 76916 588134
rect 77152 587898 82847 588134
rect 83083 587898 103916 588134
rect 104152 587898 109847 588134
rect 110083 587898 130916 588134
rect 131152 587898 136847 588134
rect 137083 587898 157916 588134
rect 158152 587898 163847 588134
rect 164083 587898 184916 588134
rect 185152 587898 190847 588134
rect 191083 587898 211916 588134
rect 212152 587898 217847 588134
rect 218083 587898 238916 588134
rect 239152 587898 244847 588134
rect 245083 587898 265916 588134
rect 266152 587898 271847 588134
rect 272083 587898 292916 588134
rect 293152 587898 298847 588134
rect 299083 587898 319916 588134
rect 320152 587898 325847 588134
rect 326083 587898 346916 588134
rect 347152 587898 352847 588134
rect 353083 587898 373916 588134
rect 374152 587898 379847 588134
rect 380083 587898 400916 588134
rect 401152 587898 406847 588134
rect 407083 587898 427916 588134
rect 428152 587898 433847 588134
rect 434083 587898 454916 588134
rect 455152 587898 460847 588134
rect 461083 587898 481916 588134
rect 482152 587898 487847 588134
rect 488083 587898 508916 588134
rect 509152 587898 514847 588134
rect 515083 587898 535916 588134
rect 536152 587898 541847 588134
rect 542083 587898 568826 588134
rect 569062 587898 569146 588134
rect 569382 587898 586302 588134
rect 586538 587898 586622 588134
rect 586858 587898 586890 588134
rect -2966 587866 586890 587898
rect 28794 580394 551414 580426
rect 28794 580158 28826 580394
rect 29062 580158 29146 580394
rect 29382 580158 46826 580394
rect 47062 580158 47146 580394
rect 47382 580158 64826 580394
rect 65062 580158 65146 580394
rect 65382 580158 82826 580394
rect 83062 580158 83146 580394
rect 83382 580158 100826 580394
rect 101062 580158 101146 580394
rect 101382 580158 118826 580394
rect 119062 580158 119146 580394
rect 119382 580158 136826 580394
rect 137062 580158 137146 580394
rect 137382 580158 154826 580394
rect 155062 580158 155146 580394
rect 155382 580158 172826 580394
rect 173062 580158 173146 580394
rect 173382 580158 190826 580394
rect 191062 580158 191146 580394
rect 191382 580158 208826 580394
rect 209062 580158 209146 580394
rect 209382 580158 226826 580394
rect 227062 580158 227146 580394
rect 227382 580158 244826 580394
rect 245062 580158 245146 580394
rect 245382 580158 262826 580394
rect 263062 580158 263146 580394
rect 263382 580158 280826 580394
rect 281062 580158 281146 580394
rect 281382 580158 298826 580394
rect 299062 580158 299146 580394
rect 299382 580158 316826 580394
rect 317062 580158 317146 580394
rect 317382 580158 334826 580394
rect 335062 580158 335146 580394
rect 335382 580158 352826 580394
rect 353062 580158 353146 580394
rect 353382 580158 370826 580394
rect 371062 580158 371146 580394
rect 371382 580158 388826 580394
rect 389062 580158 389146 580394
rect 389382 580158 406826 580394
rect 407062 580158 407146 580394
rect 407382 580158 424826 580394
rect 425062 580158 425146 580394
rect 425382 580158 442826 580394
rect 443062 580158 443146 580394
rect 443382 580158 460826 580394
rect 461062 580158 461146 580394
rect 461382 580158 478826 580394
rect 479062 580158 479146 580394
rect 479382 580158 496826 580394
rect 497062 580158 497146 580394
rect 497382 580158 514826 580394
rect 515062 580158 515146 580394
rect 515382 580158 532826 580394
rect 533062 580158 533146 580394
rect 533382 580158 550826 580394
rect 551062 580158 551146 580394
rect 551382 580158 551414 580394
rect 28794 580074 551414 580158
rect 28794 579838 28826 580074
rect 29062 579838 29146 580074
rect 29382 579838 46826 580074
rect 47062 579838 47146 580074
rect 47382 579838 64826 580074
rect 65062 579838 65146 580074
rect 65382 579838 82826 580074
rect 83062 579838 83146 580074
rect 83382 579838 100826 580074
rect 101062 579838 101146 580074
rect 101382 579838 118826 580074
rect 119062 579838 119146 580074
rect 119382 579838 136826 580074
rect 137062 579838 137146 580074
rect 137382 579838 154826 580074
rect 155062 579838 155146 580074
rect 155382 579838 172826 580074
rect 173062 579838 173146 580074
rect 173382 579838 190826 580074
rect 191062 579838 191146 580074
rect 191382 579838 208826 580074
rect 209062 579838 209146 580074
rect 209382 579838 226826 580074
rect 227062 579838 227146 580074
rect 227382 579838 244826 580074
rect 245062 579838 245146 580074
rect 245382 579838 262826 580074
rect 263062 579838 263146 580074
rect 263382 579838 280826 580074
rect 281062 579838 281146 580074
rect 281382 579838 298826 580074
rect 299062 579838 299146 580074
rect 299382 579838 316826 580074
rect 317062 579838 317146 580074
rect 317382 579838 334826 580074
rect 335062 579838 335146 580074
rect 335382 579838 352826 580074
rect 353062 579838 353146 580074
rect 353382 579838 370826 580074
rect 371062 579838 371146 580074
rect 371382 579838 388826 580074
rect 389062 579838 389146 580074
rect 389382 579838 406826 580074
rect 407062 579838 407146 580074
rect 407382 579838 424826 580074
rect 425062 579838 425146 580074
rect 425382 579838 442826 580074
rect 443062 579838 443146 580074
rect 443382 579838 460826 580074
rect 461062 579838 461146 580074
rect 461382 579838 478826 580074
rect 479062 579838 479146 580074
rect 479382 579838 496826 580074
rect 497062 579838 497146 580074
rect 497382 579838 514826 580074
rect 515062 579838 515146 580074
rect 515382 579838 532826 580074
rect 533062 579838 533146 580074
rect 533382 579838 550826 580074
rect 551062 579838 551146 580074
rect 551382 579838 551414 580074
rect 28794 579806 551414 579838
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 19826 579454
rect 20062 579218 20146 579454
rect 20382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 55826 579454
rect 56062 579218 56146 579454
rect 56382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 91826 579454
rect 92062 579218 92146 579454
rect 92382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 127826 579454
rect 128062 579218 128146 579454
rect 128382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 163826 579454
rect 164062 579218 164146 579454
rect 164382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 199826 579454
rect 200062 579218 200146 579454
rect 200382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 235826 579454
rect 236062 579218 236146 579454
rect 236382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 271826 579454
rect 272062 579218 272146 579454
rect 272382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 307826 579454
rect 308062 579218 308146 579454
rect 308382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 343826 579454
rect 344062 579218 344146 579454
rect 344382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 379826 579454
rect 380062 579218 380146 579454
rect 380382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 415826 579454
rect 416062 579218 416146 579454
rect 416382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 451826 579454
rect 452062 579218 452146 579454
rect 452382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 487826 579454
rect 488062 579218 488146 579454
rect 488382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 523826 579454
rect 524062 579218 524146 579454
rect 524382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 559826 579454
rect 560062 579218 560146 579454
rect 560382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 19826 579134
rect 20062 578898 20146 579134
rect 20382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 55826 579134
rect 56062 578898 56146 579134
rect 56382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 91826 579134
rect 92062 578898 92146 579134
rect 92382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 127826 579134
rect 128062 578898 128146 579134
rect 128382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 163826 579134
rect 164062 578898 164146 579134
rect 164382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 199826 579134
rect 200062 578898 200146 579134
rect 200382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 235826 579134
rect 236062 578898 236146 579134
rect 236382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 271826 579134
rect 272062 578898 272146 579134
rect 272382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 307826 579134
rect 308062 578898 308146 579134
rect 308382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 343826 579134
rect 344062 578898 344146 579134
rect 344382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 379826 579134
rect 380062 578898 380146 579134
rect 380382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 415826 579134
rect 416062 578898 416146 579134
rect 416382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 451826 579134
rect 452062 578898 452146 579134
rect 452382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 487826 579134
rect 488062 578898 488146 579134
rect 488382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 523826 579134
rect 524062 578898 524146 579134
rect 524382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 559826 579134
rect 560062 578898 560146 579134
rect 560382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -2966 570454 586890 570486
rect -2966 570218 -2934 570454
rect -2698 570218 -2614 570454
rect -2378 570218 10826 570454
rect 11062 570218 11146 570454
rect 11382 570218 22916 570454
rect 23152 570218 28847 570454
rect 29083 570218 49916 570454
rect 50152 570218 55847 570454
rect 56083 570218 76916 570454
rect 77152 570218 82847 570454
rect 83083 570218 103916 570454
rect 104152 570218 109847 570454
rect 110083 570218 130916 570454
rect 131152 570218 136847 570454
rect 137083 570218 157916 570454
rect 158152 570218 163847 570454
rect 164083 570218 184916 570454
rect 185152 570218 190847 570454
rect 191083 570218 211916 570454
rect 212152 570218 217847 570454
rect 218083 570218 238916 570454
rect 239152 570218 244847 570454
rect 245083 570218 265916 570454
rect 266152 570218 271847 570454
rect 272083 570218 292916 570454
rect 293152 570218 298847 570454
rect 299083 570218 319916 570454
rect 320152 570218 325847 570454
rect 326083 570218 346916 570454
rect 347152 570218 352847 570454
rect 353083 570218 373916 570454
rect 374152 570218 379847 570454
rect 380083 570218 400916 570454
rect 401152 570218 406847 570454
rect 407083 570218 427916 570454
rect 428152 570218 433847 570454
rect 434083 570218 454916 570454
rect 455152 570218 460847 570454
rect 461083 570218 481916 570454
rect 482152 570218 487847 570454
rect 488083 570218 508916 570454
rect 509152 570218 514847 570454
rect 515083 570218 535916 570454
rect 536152 570218 541847 570454
rect 542083 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 586302 570454
rect 586538 570218 586622 570454
rect 586858 570218 586890 570454
rect -2966 570134 586890 570218
rect -2966 569898 -2934 570134
rect -2698 569898 -2614 570134
rect -2378 569898 10826 570134
rect 11062 569898 11146 570134
rect 11382 569898 22916 570134
rect 23152 569898 28847 570134
rect 29083 569898 49916 570134
rect 50152 569898 55847 570134
rect 56083 569898 76916 570134
rect 77152 569898 82847 570134
rect 83083 569898 103916 570134
rect 104152 569898 109847 570134
rect 110083 569898 130916 570134
rect 131152 569898 136847 570134
rect 137083 569898 157916 570134
rect 158152 569898 163847 570134
rect 164083 569898 184916 570134
rect 185152 569898 190847 570134
rect 191083 569898 211916 570134
rect 212152 569898 217847 570134
rect 218083 569898 238916 570134
rect 239152 569898 244847 570134
rect 245083 569898 265916 570134
rect 266152 569898 271847 570134
rect 272083 569898 292916 570134
rect 293152 569898 298847 570134
rect 299083 569898 319916 570134
rect 320152 569898 325847 570134
rect 326083 569898 346916 570134
rect 347152 569898 352847 570134
rect 353083 569898 373916 570134
rect 374152 569898 379847 570134
rect 380083 569898 400916 570134
rect 401152 569898 406847 570134
rect 407083 569898 427916 570134
rect 428152 569898 433847 570134
rect 434083 569898 454916 570134
rect 455152 569898 460847 570134
rect 461083 569898 481916 570134
rect 482152 569898 487847 570134
rect 488083 569898 508916 570134
rect 509152 569898 514847 570134
rect 515083 569898 535916 570134
rect 536152 569898 541847 570134
rect 542083 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 586302 570134
rect 586538 569898 586622 570134
rect 586858 569898 586890 570134
rect -2966 569866 586890 569898
rect -2966 561454 586890 561486
rect -2966 561218 -1974 561454
rect -1738 561218 -1654 561454
rect -1418 561218 1826 561454
rect 2062 561218 2146 561454
rect 2382 561218 19952 561454
rect 20188 561218 25882 561454
rect 26118 561218 31813 561454
rect 32049 561218 46952 561454
rect 47188 561218 52882 561454
rect 53118 561218 58813 561454
rect 59049 561218 73952 561454
rect 74188 561218 79882 561454
rect 80118 561218 85813 561454
rect 86049 561218 100952 561454
rect 101188 561218 106882 561454
rect 107118 561218 112813 561454
rect 113049 561218 127952 561454
rect 128188 561218 133882 561454
rect 134118 561218 139813 561454
rect 140049 561218 154952 561454
rect 155188 561218 160882 561454
rect 161118 561218 166813 561454
rect 167049 561218 181952 561454
rect 182188 561218 187882 561454
rect 188118 561218 193813 561454
rect 194049 561218 208952 561454
rect 209188 561218 214882 561454
rect 215118 561218 220813 561454
rect 221049 561218 235952 561454
rect 236188 561218 241882 561454
rect 242118 561218 247813 561454
rect 248049 561218 262952 561454
rect 263188 561218 268882 561454
rect 269118 561218 274813 561454
rect 275049 561218 289952 561454
rect 290188 561218 295882 561454
rect 296118 561218 301813 561454
rect 302049 561218 316952 561454
rect 317188 561218 322882 561454
rect 323118 561218 328813 561454
rect 329049 561218 343952 561454
rect 344188 561218 349882 561454
rect 350118 561218 355813 561454
rect 356049 561218 370952 561454
rect 371188 561218 376882 561454
rect 377118 561218 382813 561454
rect 383049 561218 397952 561454
rect 398188 561218 403882 561454
rect 404118 561218 409813 561454
rect 410049 561218 424952 561454
rect 425188 561218 430882 561454
rect 431118 561218 436813 561454
rect 437049 561218 451952 561454
rect 452188 561218 457882 561454
rect 458118 561218 463813 561454
rect 464049 561218 478952 561454
rect 479188 561218 484882 561454
rect 485118 561218 490813 561454
rect 491049 561218 505952 561454
rect 506188 561218 511882 561454
rect 512118 561218 517813 561454
rect 518049 561218 532952 561454
rect 533188 561218 538882 561454
rect 539118 561218 544813 561454
rect 545049 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 577826 561454
rect 578062 561218 578146 561454
rect 578382 561218 585342 561454
rect 585578 561218 585662 561454
rect 585898 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -1974 561134
rect -1738 560898 -1654 561134
rect -1418 560898 1826 561134
rect 2062 560898 2146 561134
rect 2382 560898 19952 561134
rect 20188 560898 25882 561134
rect 26118 560898 31813 561134
rect 32049 560898 46952 561134
rect 47188 560898 52882 561134
rect 53118 560898 58813 561134
rect 59049 560898 73952 561134
rect 74188 560898 79882 561134
rect 80118 560898 85813 561134
rect 86049 560898 100952 561134
rect 101188 560898 106882 561134
rect 107118 560898 112813 561134
rect 113049 560898 127952 561134
rect 128188 560898 133882 561134
rect 134118 560898 139813 561134
rect 140049 560898 154952 561134
rect 155188 560898 160882 561134
rect 161118 560898 166813 561134
rect 167049 560898 181952 561134
rect 182188 560898 187882 561134
rect 188118 560898 193813 561134
rect 194049 560898 208952 561134
rect 209188 560898 214882 561134
rect 215118 560898 220813 561134
rect 221049 560898 235952 561134
rect 236188 560898 241882 561134
rect 242118 560898 247813 561134
rect 248049 560898 262952 561134
rect 263188 560898 268882 561134
rect 269118 560898 274813 561134
rect 275049 560898 289952 561134
rect 290188 560898 295882 561134
rect 296118 560898 301813 561134
rect 302049 560898 316952 561134
rect 317188 560898 322882 561134
rect 323118 560898 328813 561134
rect 329049 560898 343952 561134
rect 344188 560898 349882 561134
rect 350118 560898 355813 561134
rect 356049 560898 370952 561134
rect 371188 560898 376882 561134
rect 377118 560898 382813 561134
rect 383049 560898 397952 561134
rect 398188 560898 403882 561134
rect 404118 560898 409813 561134
rect 410049 560898 424952 561134
rect 425188 560898 430882 561134
rect 431118 560898 436813 561134
rect 437049 560898 451952 561134
rect 452188 560898 457882 561134
rect 458118 560898 463813 561134
rect 464049 560898 478952 561134
rect 479188 560898 484882 561134
rect 485118 560898 490813 561134
rect 491049 560898 505952 561134
rect 506188 560898 511882 561134
rect 512118 560898 517813 561134
rect 518049 560898 532952 561134
rect 533188 560898 538882 561134
rect 539118 560898 544813 561134
rect 545049 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 577826 561134
rect 578062 560898 578146 561134
rect 578382 560898 585342 561134
rect 585578 560898 585662 561134
rect 585898 560898 586890 561134
rect -2966 560866 586890 560898
rect 19794 553394 542414 553426
rect 19794 553158 19826 553394
rect 20062 553158 20146 553394
rect 20382 553158 37826 553394
rect 38062 553158 38146 553394
rect 38382 553158 55826 553394
rect 56062 553158 56146 553394
rect 56382 553158 73826 553394
rect 74062 553158 74146 553394
rect 74382 553158 91826 553394
rect 92062 553158 92146 553394
rect 92382 553158 109826 553394
rect 110062 553158 110146 553394
rect 110382 553158 127826 553394
rect 128062 553158 128146 553394
rect 128382 553158 145826 553394
rect 146062 553158 146146 553394
rect 146382 553158 163826 553394
rect 164062 553158 164146 553394
rect 164382 553158 181826 553394
rect 182062 553158 182146 553394
rect 182382 553158 199826 553394
rect 200062 553158 200146 553394
rect 200382 553158 217826 553394
rect 218062 553158 218146 553394
rect 218382 553158 235826 553394
rect 236062 553158 236146 553394
rect 236382 553158 253826 553394
rect 254062 553158 254146 553394
rect 254382 553158 271826 553394
rect 272062 553158 272146 553394
rect 272382 553158 289826 553394
rect 290062 553158 290146 553394
rect 290382 553158 307826 553394
rect 308062 553158 308146 553394
rect 308382 553158 325826 553394
rect 326062 553158 326146 553394
rect 326382 553158 343826 553394
rect 344062 553158 344146 553394
rect 344382 553158 361826 553394
rect 362062 553158 362146 553394
rect 362382 553158 379826 553394
rect 380062 553158 380146 553394
rect 380382 553158 397826 553394
rect 398062 553158 398146 553394
rect 398382 553158 415826 553394
rect 416062 553158 416146 553394
rect 416382 553158 433826 553394
rect 434062 553158 434146 553394
rect 434382 553158 451826 553394
rect 452062 553158 452146 553394
rect 452382 553158 469826 553394
rect 470062 553158 470146 553394
rect 470382 553158 487826 553394
rect 488062 553158 488146 553394
rect 488382 553158 505826 553394
rect 506062 553158 506146 553394
rect 506382 553158 523826 553394
rect 524062 553158 524146 553394
rect 524382 553158 541826 553394
rect 542062 553158 542146 553394
rect 542382 553158 542414 553394
rect 19794 553074 542414 553158
rect 19794 552838 19826 553074
rect 20062 552838 20146 553074
rect 20382 552838 37826 553074
rect 38062 552838 38146 553074
rect 38382 552838 55826 553074
rect 56062 552838 56146 553074
rect 56382 552838 73826 553074
rect 74062 552838 74146 553074
rect 74382 552838 91826 553074
rect 92062 552838 92146 553074
rect 92382 552838 109826 553074
rect 110062 552838 110146 553074
rect 110382 552838 127826 553074
rect 128062 552838 128146 553074
rect 128382 552838 145826 553074
rect 146062 552838 146146 553074
rect 146382 552838 163826 553074
rect 164062 552838 164146 553074
rect 164382 552838 181826 553074
rect 182062 552838 182146 553074
rect 182382 552838 199826 553074
rect 200062 552838 200146 553074
rect 200382 552838 217826 553074
rect 218062 552838 218146 553074
rect 218382 552838 235826 553074
rect 236062 552838 236146 553074
rect 236382 552838 253826 553074
rect 254062 552838 254146 553074
rect 254382 552838 271826 553074
rect 272062 552838 272146 553074
rect 272382 552838 289826 553074
rect 290062 552838 290146 553074
rect 290382 552838 307826 553074
rect 308062 552838 308146 553074
rect 308382 552838 325826 553074
rect 326062 552838 326146 553074
rect 326382 552838 343826 553074
rect 344062 552838 344146 553074
rect 344382 552838 361826 553074
rect 362062 552838 362146 553074
rect 362382 552838 379826 553074
rect 380062 552838 380146 553074
rect 380382 552838 397826 553074
rect 398062 552838 398146 553074
rect 398382 552838 415826 553074
rect 416062 552838 416146 553074
rect 416382 552838 433826 553074
rect 434062 552838 434146 553074
rect 434382 552838 451826 553074
rect 452062 552838 452146 553074
rect 452382 552838 469826 553074
rect 470062 552838 470146 553074
rect 470382 552838 487826 553074
rect 488062 552838 488146 553074
rect 488382 552838 505826 553074
rect 506062 552838 506146 553074
rect 506382 552838 523826 553074
rect 524062 552838 524146 553074
rect 524382 552838 541826 553074
rect 542062 552838 542146 553074
rect 542382 552838 542414 553074
rect 19794 552806 542414 552838
rect -2966 552454 586890 552486
rect -2966 552218 -2934 552454
rect -2698 552218 -2614 552454
rect -2378 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 28826 552454
rect 29062 552218 29146 552454
rect 29382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 64826 552454
rect 65062 552218 65146 552454
rect 65382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 100826 552454
rect 101062 552218 101146 552454
rect 101382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 136826 552454
rect 137062 552218 137146 552454
rect 137382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 172826 552454
rect 173062 552218 173146 552454
rect 173382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 208826 552454
rect 209062 552218 209146 552454
rect 209382 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 244826 552454
rect 245062 552218 245146 552454
rect 245382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 280826 552454
rect 281062 552218 281146 552454
rect 281382 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 316826 552454
rect 317062 552218 317146 552454
rect 317382 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 352826 552454
rect 353062 552218 353146 552454
rect 353382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 388826 552454
rect 389062 552218 389146 552454
rect 389382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 424826 552454
rect 425062 552218 425146 552454
rect 425382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 460826 552454
rect 461062 552218 461146 552454
rect 461382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 496826 552454
rect 497062 552218 497146 552454
rect 497382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 532826 552454
rect 533062 552218 533146 552454
rect 533382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 568826 552454
rect 569062 552218 569146 552454
rect 569382 552218 586302 552454
rect 586538 552218 586622 552454
rect 586858 552218 586890 552454
rect -2966 552134 586890 552218
rect -2966 551898 -2934 552134
rect -2698 551898 -2614 552134
rect -2378 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 28826 552134
rect 29062 551898 29146 552134
rect 29382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 64826 552134
rect 65062 551898 65146 552134
rect 65382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 100826 552134
rect 101062 551898 101146 552134
rect 101382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 136826 552134
rect 137062 551898 137146 552134
rect 137382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 172826 552134
rect 173062 551898 173146 552134
rect 173382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 208826 552134
rect 209062 551898 209146 552134
rect 209382 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 244826 552134
rect 245062 551898 245146 552134
rect 245382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 280826 552134
rect 281062 551898 281146 552134
rect 281382 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 316826 552134
rect 317062 551898 317146 552134
rect 317382 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 352826 552134
rect 353062 551898 353146 552134
rect 353382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 388826 552134
rect 389062 551898 389146 552134
rect 389382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 424826 552134
rect 425062 551898 425146 552134
rect 425382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 460826 552134
rect 461062 551898 461146 552134
rect 461382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 496826 552134
rect 497062 551898 497146 552134
rect 497382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 532826 552134
rect 533062 551898 533146 552134
rect 533382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 568826 552134
rect 569062 551898 569146 552134
rect 569382 551898 586302 552134
rect 586538 551898 586622 552134
rect 586858 551898 586890 552134
rect -2966 551866 586890 551898
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 19952 543454
rect 20188 543218 25882 543454
rect 26118 543218 31813 543454
rect 32049 543218 46952 543454
rect 47188 543218 52882 543454
rect 53118 543218 58813 543454
rect 59049 543218 73952 543454
rect 74188 543218 79882 543454
rect 80118 543218 85813 543454
rect 86049 543218 100952 543454
rect 101188 543218 106882 543454
rect 107118 543218 112813 543454
rect 113049 543218 127952 543454
rect 128188 543218 133882 543454
rect 134118 543218 139813 543454
rect 140049 543218 154952 543454
rect 155188 543218 160882 543454
rect 161118 543218 166813 543454
rect 167049 543218 181952 543454
rect 182188 543218 187882 543454
rect 188118 543218 193813 543454
rect 194049 543218 208952 543454
rect 209188 543218 214882 543454
rect 215118 543218 220813 543454
rect 221049 543218 235952 543454
rect 236188 543218 241882 543454
rect 242118 543218 247813 543454
rect 248049 543218 262952 543454
rect 263188 543218 268882 543454
rect 269118 543218 274813 543454
rect 275049 543218 289952 543454
rect 290188 543218 295882 543454
rect 296118 543218 301813 543454
rect 302049 543218 316952 543454
rect 317188 543218 322882 543454
rect 323118 543218 328813 543454
rect 329049 543218 343952 543454
rect 344188 543218 349882 543454
rect 350118 543218 355813 543454
rect 356049 543218 370952 543454
rect 371188 543218 376882 543454
rect 377118 543218 382813 543454
rect 383049 543218 397952 543454
rect 398188 543218 403882 543454
rect 404118 543218 409813 543454
rect 410049 543218 424952 543454
rect 425188 543218 430882 543454
rect 431118 543218 436813 543454
rect 437049 543218 451952 543454
rect 452188 543218 457882 543454
rect 458118 543218 463813 543454
rect 464049 543218 478952 543454
rect 479188 543218 484882 543454
rect 485118 543218 490813 543454
rect 491049 543218 505952 543454
rect 506188 543218 511882 543454
rect 512118 543218 517813 543454
rect 518049 543218 532952 543454
rect 533188 543218 538882 543454
rect 539118 543218 544813 543454
rect 545049 543218 559826 543454
rect 560062 543218 560146 543454
rect 560382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 19952 543134
rect 20188 542898 25882 543134
rect 26118 542898 31813 543134
rect 32049 542898 46952 543134
rect 47188 542898 52882 543134
rect 53118 542898 58813 543134
rect 59049 542898 73952 543134
rect 74188 542898 79882 543134
rect 80118 542898 85813 543134
rect 86049 542898 100952 543134
rect 101188 542898 106882 543134
rect 107118 542898 112813 543134
rect 113049 542898 127952 543134
rect 128188 542898 133882 543134
rect 134118 542898 139813 543134
rect 140049 542898 154952 543134
rect 155188 542898 160882 543134
rect 161118 542898 166813 543134
rect 167049 542898 181952 543134
rect 182188 542898 187882 543134
rect 188118 542898 193813 543134
rect 194049 542898 208952 543134
rect 209188 542898 214882 543134
rect 215118 542898 220813 543134
rect 221049 542898 235952 543134
rect 236188 542898 241882 543134
rect 242118 542898 247813 543134
rect 248049 542898 262952 543134
rect 263188 542898 268882 543134
rect 269118 542898 274813 543134
rect 275049 542898 289952 543134
rect 290188 542898 295882 543134
rect 296118 542898 301813 543134
rect 302049 542898 316952 543134
rect 317188 542898 322882 543134
rect 323118 542898 328813 543134
rect 329049 542898 343952 543134
rect 344188 542898 349882 543134
rect 350118 542898 355813 543134
rect 356049 542898 370952 543134
rect 371188 542898 376882 543134
rect 377118 542898 382813 543134
rect 383049 542898 397952 543134
rect 398188 542898 403882 543134
rect 404118 542898 409813 543134
rect 410049 542898 424952 543134
rect 425188 542898 430882 543134
rect 431118 542898 436813 543134
rect 437049 542898 451952 543134
rect 452188 542898 457882 543134
rect 458118 542898 463813 543134
rect 464049 542898 478952 543134
rect 479188 542898 484882 543134
rect 485118 542898 490813 543134
rect 491049 542898 505952 543134
rect 506188 542898 511882 543134
rect 512118 542898 517813 543134
rect 518049 542898 532952 543134
rect 533188 542898 538882 543134
rect 539118 542898 544813 543134
rect 545049 542898 559826 543134
rect 560062 542898 560146 543134
rect 560382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -2966 534454 586890 534486
rect -2966 534218 -2934 534454
rect -2698 534218 -2614 534454
rect -2378 534218 10826 534454
rect 11062 534218 11146 534454
rect 11382 534218 22916 534454
rect 23152 534218 28847 534454
rect 29083 534218 49916 534454
rect 50152 534218 55847 534454
rect 56083 534218 76916 534454
rect 77152 534218 82847 534454
rect 83083 534218 103916 534454
rect 104152 534218 109847 534454
rect 110083 534218 130916 534454
rect 131152 534218 136847 534454
rect 137083 534218 157916 534454
rect 158152 534218 163847 534454
rect 164083 534218 184916 534454
rect 185152 534218 190847 534454
rect 191083 534218 211916 534454
rect 212152 534218 217847 534454
rect 218083 534218 238916 534454
rect 239152 534218 244847 534454
rect 245083 534218 265916 534454
rect 266152 534218 271847 534454
rect 272083 534218 292916 534454
rect 293152 534218 298847 534454
rect 299083 534218 319916 534454
rect 320152 534218 325847 534454
rect 326083 534218 346916 534454
rect 347152 534218 352847 534454
rect 353083 534218 373916 534454
rect 374152 534218 379847 534454
rect 380083 534218 400916 534454
rect 401152 534218 406847 534454
rect 407083 534218 427916 534454
rect 428152 534218 433847 534454
rect 434083 534218 454916 534454
rect 455152 534218 460847 534454
rect 461083 534218 481916 534454
rect 482152 534218 487847 534454
rect 488083 534218 508916 534454
rect 509152 534218 514847 534454
rect 515083 534218 535916 534454
rect 536152 534218 541847 534454
rect 542083 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 586302 534454
rect 586538 534218 586622 534454
rect 586858 534218 586890 534454
rect -2966 534134 586890 534218
rect -2966 533898 -2934 534134
rect -2698 533898 -2614 534134
rect -2378 533898 10826 534134
rect 11062 533898 11146 534134
rect 11382 533898 22916 534134
rect 23152 533898 28847 534134
rect 29083 533898 49916 534134
rect 50152 533898 55847 534134
rect 56083 533898 76916 534134
rect 77152 533898 82847 534134
rect 83083 533898 103916 534134
rect 104152 533898 109847 534134
rect 110083 533898 130916 534134
rect 131152 533898 136847 534134
rect 137083 533898 157916 534134
rect 158152 533898 163847 534134
rect 164083 533898 184916 534134
rect 185152 533898 190847 534134
rect 191083 533898 211916 534134
rect 212152 533898 217847 534134
rect 218083 533898 238916 534134
rect 239152 533898 244847 534134
rect 245083 533898 265916 534134
rect 266152 533898 271847 534134
rect 272083 533898 292916 534134
rect 293152 533898 298847 534134
rect 299083 533898 319916 534134
rect 320152 533898 325847 534134
rect 326083 533898 346916 534134
rect 347152 533898 352847 534134
rect 353083 533898 373916 534134
rect 374152 533898 379847 534134
rect 380083 533898 400916 534134
rect 401152 533898 406847 534134
rect 407083 533898 427916 534134
rect 428152 533898 433847 534134
rect 434083 533898 454916 534134
rect 455152 533898 460847 534134
rect 461083 533898 481916 534134
rect 482152 533898 487847 534134
rect 488083 533898 508916 534134
rect 509152 533898 514847 534134
rect 515083 533898 535916 534134
rect 536152 533898 541847 534134
rect 542083 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 586302 534134
rect 586538 533898 586622 534134
rect 586858 533898 586890 534134
rect -2966 533866 586890 533898
rect 28794 526394 551414 526426
rect 28794 526158 28826 526394
rect 29062 526158 29146 526394
rect 29382 526158 46826 526394
rect 47062 526158 47146 526394
rect 47382 526158 64826 526394
rect 65062 526158 65146 526394
rect 65382 526158 82826 526394
rect 83062 526158 83146 526394
rect 83382 526158 100826 526394
rect 101062 526158 101146 526394
rect 101382 526158 118826 526394
rect 119062 526158 119146 526394
rect 119382 526158 136826 526394
rect 137062 526158 137146 526394
rect 137382 526158 154826 526394
rect 155062 526158 155146 526394
rect 155382 526158 172826 526394
rect 173062 526158 173146 526394
rect 173382 526158 190826 526394
rect 191062 526158 191146 526394
rect 191382 526158 208826 526394
rect 209062 526158 209146 526394
rect 209382 526158 226826 526394
rect 227062 526158 227146 526394
rect 227382 526158 244826 526394
rect 245062 526158 245146 526394
rect 245382 526158 262826 526394
rect 263062 526158 263146 526394
rect 263382 526158 280826 526394
rect 281062 526158 281146 526394
rect 281382 526158 298826 526394
rect 299062 526158 299146 526394
rect 299382 526158 316826 526394
rect 317062 526158 317146 526394
rect 317382 526158 334826 526394
rect 335062 526158 335146 526394
rect 335382 526158 352826 526394
rect 353062 526158 353146 526394
rect 353382 526158 370826 526394
rect 371062 526158 371146 526394
rect 371382 526158 388826 526394
rect 389062 526158 389146 526394
rect 389382 526158 406826 526394
rect 407062 526158 407146 526394
rect 407382 526158 424826 526394
rect 425062 526158 425146 526394
rect 425382 526158 442826 526394
rect 443062 526158 443146 526394
rect 443382 526158 460826 526394
rect 461062 526158 461146 526394
rect 461382 526158 478826 526394
rect 479062 526158 479146 526394
rect 479382 526158 496826 526394
rect 497062 526158 497146 526394
rect 497382 526158 514826 526394
rect 515062 526158 515146 526394
rect 515382 526158 532826 526394
rect 533062 526158 533146 526394
rect 533382 526158 550826 526394
rect 551062 526158 551146 526394
rect 551382 526158 551414 526394
rect 28794 526074 551414 526158
rect 28794 525838 28826 526074
rect 29062 525838 29146 526074
rect 29382 525838 46826 526074
rect 47062 525838 47146 526074
rect 47382 525838 64826 526074
rect 65062 525838 65146 526074
rect 65382 525838 82826 526074
rect 83062 525838 83146 526074
rect 83382 525838 100826 526074
rect 101062 525838 101146 526074
rect 101382 525838 118826 526074
rect 119062 525838 119146 526074
rect 119382 525838 136826 526074
rect 137062 525838 137146 526074
rect 137382 525838 154826 526074
rect 155062 525838 155146 526074
rect 155382 525838 172826 526074
rect 173062 525838 173146 526074
rect 173382 525838 190826 526074
rect 191062 525838 191146 526074
rect 191382 525838 208826 526074
rect 209062 525838 209146 526074
rect 209382 525838 226826 526074
rect 227062 525838 227146 526074
rect 227382 525838 244826 526074
rect 245062 525838 245146 526074
rect 245382 525838 262826 526074
rect 263062 525838 263146 526074
rect 263382 525838 280826 526074
rect 281062 525838 281146 526074
rect 281382 525838 298826 526074
rect 299062 525838 299146 526074
rect 299382 525838 316826 526074
rect 317062 525838 317146 526074
rect 317382 525838 334826 526074
rect 335062 525838 335146 526074
rect 335382 525838 352826 526074
rect 353062 525838 353146 526074
rect 353382 525838 370826 526074
rect 371062 525838 371146 526074
rect 371382 525838 388826 526074
rect 389062 525838 389146 526074
rect 389382 525838 406826 526074
rect 407062 525838 407146 526074
rect 407382 525838 424826 526074
rect 425062 525838 425146 526074
rect 425382 525838 442826 526074
rect 443062 525838 443146 526074
rect 443382 525838 460826 526074
rect 461062 525838 461146 526074
rect 461382 525838 478826 526074
rect 479062 525838 479146 526074
rect 479382 525838 496826 526074
rect 497062 525838 497146 526074
rect 497382 525838 514826 526074
rect 515062 525838 515146 526074
rect 515382 525838 532826 526074
rect 533062 525838 533146 526074
rect 533382 525838 550826 526074
rect 551062 525838 551146 526074
rect 551382 525838 551414 526074
rect 28794 525806 551414 525838
rect -2966 525454 586890 525486
rect -2966 525218 -1974 525454
rect -1738 525218 -1654 525454
rect -1418 525218 1826 525454
rect 2062 525218 2146 525454
rect 2382 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 37826 525454
rect 38062 525218 38146 525454
rect 38382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 73826 525454
rect 74062 525218 74146 525454
rect 74382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 109826 525454
rect 110062 525218 110146 525454
rect 110382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 145826 525454
rect 146062 525218 146146 525454
rect 146382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 181826 525454
rect 182062 525218 182146 525454
rect 182382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 217826 525454
rect 218062 525218 218146 525454
rect 218382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 253826 525454
rect 254062 525218 254146 525454
rect 254382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 289826 525454
rect 290062 525218 290146 525454
rect 290382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 325826 525454
rect 326062 525218 326146 525454
rect 326382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 361826 525454
rect 362062 525218 362146 525454
rect 362382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 397826 525454
rect 398062 525218 398146 525454
rect 398382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 433826 525454
rect 434062 525218 434146 525454
rect 434382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 469826 525454
rect 470062 525218 470146 525454
rect 470382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 505826 525454
rect 506062 525218 506146 525454
rect 506382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 541826 525454
rect 542062 525218 542146 525454
rect 542382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 577826 525454
rect 578062 525218 578146 525454
rect 578382 525218 585342 525454
rect 585578 525218 585662 525454
rect 585898 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -1974 525134
rect -1738 524898 -1654 525134
rect -1418 524898 1826 525134
rect 2062 524898 2146 525134
rect 2382 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 37826 525134
rect 38062 524898 38146 525134
rect 38382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 73826 525134
rect 74062 524898 74146 525134
rect 74382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 109826 525134
rect 110062 524898 110146 525134
rect 110382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 145826 525134
rect 146062 524898 146146 525134
rect 146382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 181826 525134
rect 182062 524898 182146 525134
rect 182382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 217826 525134
rect 218062 524898 218146 525134
rect 218382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 253826 525134
rect 254062 524898 254146 525134
rect 254382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 289826 525134
rect 290062 524898 290146 525134
rect 290382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 325826 525134
rect 326062 524898 326146 525134
rect 326382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 361826 525134
rect 362062 524898 362146 525134
rect 362382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 397826 525134
rect 398062 524898 398146 525134
rect 398382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 433826 525134
rect 434062 524898 434146 525134
rect 434382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 469826 525134
rect 470062 524898 470146 525134
rect 470382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 505826 525134
rect 506062 524898 506146 525134
rect 506382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 541826 525134
rect 542062 524898 542146 525134
rect 542382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 577826 525134
rect 578062 524898 578146 525134
rect 578382 524898 585342 525134
rect 585578 524898 585662 525134
rect 585898 524898 586890 525134
rect -2966 524866 586890 524898
rect -2966 516454 586890 516486
rect -2966 516218 -2934 516454
rect -2698 516218 -2614 516454
rect -2378 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 22916 516454
rect 23152 516218 28847 516454
rect 29083 516218 49916 516454
rect 50152 516218 55847 516454
rect 56083 516218 76916 516454
rect 77152 516218 82847 516454
rect 83083 516218 103916 516454
rect 104152 516218 109847 516454
rect 110083 516218 130916 516454
rect 131152 516218 136847 516454
rect 137083 516218 157916 516454
rect 158152 516218 163847 516454
rect 164083 516218 184916 516454
rect 185152 516218 190847 516454
rect 191083 516218 211916 516454
rect 212152 516218 217847 516454
rect 218083 516218 238916 516454
rect 239152 516218 244847 516454
rect 245083 516218 265916 516454
rect 266152 516218 271847 516454
rect 272083 516218 292916 516454
rect 293152 516218 298847 516454
rect 299083 516218 319916 516454
rect 320152 516218 325847 516454
rect 326083 516218 346916 516454
rect 347152 516218 352847 516454
rect 353083 516218 373916 516454
rect 374152 516218 379847 516454
rect 380083 516218 400916 516454
rect 401152 516218 406847 516454
rect 407083 516218 427916 516454
rect 428152 516218 433847 516454
rect 434083 516218 454916 516454
rect 455152 516218 460847 516454
rect 461083 516218 481916 516454
rect 482152 516218 487847 516454
rect 488083 516218 508916 516454
rect 509152 516218 514847 516454
rect 515083 516218 535916 516454
rect 536152 516218 541847 516454
rect 542083 516218 568826 516454
rect 569062 516218 569146 516454
rect 569382 516218 586302 516454
rect 586538 516218 586622 516454
rect 586858 516218 586890 516454
rect -2966 516134 586890 516218
rect -2966 515898 -2934 516134
rect -2698 515898 -2614 516134
rect -2378 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 22916 516134
rect 23152 515898 28847 516134
rect 29083 515898 49916 516134
rect 50152 515898 55847 516134
rect 56083 515898 76916 516134
rect 77152 515898 82847 516134
rect 83083 515898 103916 516134
rect 104152 515898 109847 516134
rect 110083 515898 130916 516134
rect 131152 515898 136847 516134
rect 137083 515898 157916 516134
rect 158152 515898 163847 516134
rect 164083 515898 184916 516134
rect 185152 515898 190847 516134
rect 191083 515898 211916 516134
rect 212152 515898 217847 516134
rect 218083 515898 238916 516134
rect 239152 515898 244847 516134
rect 245083 515898 265916 516134
rect 266152 515898 271847 516134
rect 272083 515898 292916 516134
rect 293152 515898 298847 516134
rect 299083 515898 319916 516134
rect 320152 515898 325847 516134
rect 326083 515898 346916 516134
rect 347152 515898 352847 516134
rect 353083 515898 373916 516134
rect 374152 515898 379847 516134
rect 380083 515898 400916 516134
rect 401152 515898 406847 516134
rect 407083 515898 427916 516134
rect 428152 515898 433847 516134
rect 434083 515898 454916 516134
rect 455152 515898 460847 516134
rect 461083 515898 481916 516134
rect 482152 515898 487847 516134
rect 488083 515898 508916 516134
rect 509152 515898 514847 516134
rect 515083 515898 535916 516134
rect 536152 515898 541847 516134
rect 542083 515898 568826 516134
rect 569062 515898 569146 516134
rect 569382 515898 586302 516134
rect 586538 515898 586622 516134
rect 586858 515898 586890 516134
rect -2966 515866 586890 515898
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 19952 507454
rect 20188 507218 25882 507454
rect 26118 507218 31813 507454
rect 32049 507218 46952 507454
rect 47188 507218 52882 507454
rect 53118 507218 58813 507454
rect 59049 507218 73952 507454
rect 74188 507218 79882 507454
rect 80118 507218 85813 507454
rect 86049 507218 100952 507454
rect 101188 507218 106882 507454
rect 107118 507218 112813 507454
rect 113049 507218 127952 507454
rect 128188 507218 133882 507454
rect 134118 507218 139813 507454
rect 140049 507218 154952 507454
rect 155188 507218 160882 507454
rect 161118 507218 166813 507454
rect 167049 507218 181952 507454
rect 182188 507218 187882 507454
rect 188118 507218 193813 507454
rect 194049 507218 208952 507454
rect 209188 507218 214882 507454
rect 215118 507218 220813 507454
rect 221049 507218 235952 507454
rect 236188 507218 241882 507454
rect 242118 507218 247813 507454
rect 248049 507218 262952 507454
rect 263188 507218 268882 507454
rect 269118 507218 274813 507454
rect 275049 507218 289952 507454
rect 290188 507218 295882 507454
rect 296118 507218 301813 507454
rect 302049 507218 316952 507454
rect 317188 507218 322882 507454
rect 323118 507218 328813 507454
rect 329049 507218 343952 507454
rect 344188 507218 349882 507454
rect 350118 507218 355813 507454
rect 356049 507218 370952 507454
rect 371188 507218 376882 507454
rect 377118 507218 382813 507454
rect 383049 507218 397952 507454
rect 398188 507218 403882 507454
rect 404118 507218 409813 507454
rect 410049 507218 424952 507454
rect 425188 507218 430882 507454
rect 431118 507218 436813 507454
rect 437049 507218 451952 507454
rect 452188 507218 457882 507454
rect 458118 507218 463813 507454
rect 464049 507218 478952 507454
rect 479188 507218 484882 507454
rect 485118 507218 490813 507454
rect 491049 507218 505952 507454
rect 506188 507218 511882 507454
rect 512118 507218 517813 507454
rect 518049 507218 532952 507454
rect 533188 507218 538882 507454
rect 539118 507218 544813 507454
rect 545049 507218 559826 507454
rect 560062 507218 560146 507454
rect 560382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 19952 507134
rect 20188 506898 25882 507134
rect 26118 506898 31813 507134
rect 32049 506898 46952 507134
rect 47188 506898 52882 507134
rect 53118 506898 58813 507134
rect 59049 506898 73952 507134
rect 74188 506898 79882 507134
rect 80118 506898 85813 507134
rect 86049 506898 100952 507134
rect 101188 506898 106882 507134
rect 107118 506898 112813 507134
rect 113049 506898 127952 507134
rect 128188 506898 133882 507134
rect 134118 506898 139813 507134
rect 140049 506898 154952 507134
rect 155188 506898 160882 507134
rect 161118 506898 166813 507134
rect 167049 506898 181952 507134
rect 182188 506898 187882 507134
rect 188118 506898 193813 507134
rect 194049 506898 208952 507134
rect 209188 506898 214882 507134
rect 215118 506898 220813 507134
rect 221049 506898 235952 507134
rect 236188 506898 241882 507134
rect 242118 506898 247813 507134
rect 248049 506898 262952 507134
rect 263188 506898 268882 507134
rect 269118 506898 274813 507134
rect 275049 506898 289952 507134
rect 290188 506898 295882 507134
rect 296118 506898 301813 507134
rect 302049 506898 316952 507134
rect 317188 506898 322882 507134
rect 323118 506898 328813 507134
rect 329049 506898 343952 507134
rect 344188 506898 349882 507134
rect 350118 506898 355813 507134
rect 356049 506898 370952 507134
rect 371188 506898 376882 507134
rect 377118 506898 382813 507134
rect 383049 506898 397952 507134
rect 398188 506898 403882 507134
rect 404118 506898 409813 507134
rect 410049 506898 424952 507134
rect 425188 506898 430882 507134
rect 431118 506898 436813 507134
rect 437049 506898 451952 507134
rect 452188 506898 457882 507134
rect 458118 506898 463813 507134
rect 464049 506898 478952 507134
rect 479188 506898 484882 507134
rect 485118 506898 490813 507134
rect 491049 506898 505952 507134
rect 506188 506898 511882 507134
rect 512118 506898 517813 507134
rect 518049 506898 532952 507134
rect 533188 506898 538882 507134
rect 539118 506898 544813 507134
rect 545049 506898 559826 507134
rect 560062 506898 560146 507134
rect 560382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect 19794 499394 542414 499426
rect 19794 499158 19826 499394
rect 20062 499158 20146 499394
rect 20382 499158 37826 499394
rect 38062 499158 38146 499394
rect 38382 499158 55826 499394
rect 56062 499158 56146 499394
rect 56382 499158 73826 499394
rect 74062 499158 74146 499394
rect 74382 499158 91826 499394
rect 92062 499158 92146 499394
rect 92382 499158 109826 499394
rect 110062 499158 110146 499394
rect 110382 499158 127826 499394
rect 128062 499158 128146 499394
rect 128382 499158 145826 499394
rect 146062 499158 146146 499394
rect 146382 499158 163826 499394
rect 164062 499158 164146 499394
rect 164382 499158 181826 499394
rect 182062 499158 182146 499394
rect 182382 499158 199826 499394
rect 200062 499158 200146 499394
rect 200382 499158 217826 499394
rect 218062 499158 218146 499394
rect 218382 499158 235826 499394
rect 236062 499158 236146 499394
rect 236382 499158 253826 499394
rect 254062 499158 254146 499394
rect 254382 499158 271826 499394
rect 272062 499158 272146 499394
rect 272382 499158 289826 499394
rect 290062 499158 290146 499394
rect 290382 499158 307826 499394
rect 308062 499158 308146 499394
rect 308382 499158 325826 499394
rect 326062 499158 326146 499394
rect 326382 499158 343826 499394
rect 344062 499158 344146 499394
rect 344382 499158 361826 499394
rect 362062 499158 362146 499394
rect 362382 499158 379826 499394
rect 380062 499158 380146 499394
rect 380382 499158 397826 499394
rect 398062 499158 398146 499394
rect 398382 499158 415826 499394
rect 416062 499158 416146 499394
rect 416382 499158 433826 499394
rect 434062 499158 434146 499394
rect 434382 499158 451826 499394
rect 452062 499158 452146 499394
rect 452382 499158 469826 499394
rect 470062 499158 470146 499394
rect 470382 499158 487826 499394
rect 488062 499158 488146 499394
rect 488382 499158 505826 499394
rect 506062 499158 506146 499394
rect 506382 499158 523826 499394
rect 524062 499158 524146 499394
rect 524382 499158 541826 499394
rect 542062 499158 542146 499394
rect 542382 499158 542414 499394
rect 19794 499074 542414 499158
rect 19794 498838 19826 499074
rect 20062 498838 20146 499074
rect 20382 498838 37826 499074
rect 38062 498838 38146 499074
rect 38382 498838 55826 499074
rect 56062 498838 56146 499074
rect 56382 498838 73826 499074
rect 74062 498838 74146 499074
rect 74382 498838 91826 499074
rect 92062 498838 92146 499074
rect 92382 498838 109826 499074
rect 110062 498838 110146 499074
rect 110382 498838 127826 499074
rect 128062 498838 128146 499074
rect 128382 498838 145826 499074
rect 146062 498838 146146 499074
rect 146382 498838 163826 499074
rect 164062 498838 164146 499074
rect 164382 498838 181826 499074
rect 182062 498838 182146 499074
rect 182382 498838 199826 499074
rect 200062 498838 200146 499074
rect 200382 498838 217826 499074
rect 218062 498838 218146 499074
rect 218382 498838 235826 499074
rect 236062 498838 236146 499074
rect 236382 498838 253826 499074
rect 254062 498838 254146 499074
rect 254382 498838 271826 499074
rect 272062 498838 272146 499074
rect 272382 498838 289826 499074
rect 290062 498838 290146 499074
rect 290382 498838 307826 499074
rect 308062 498838 308146 499074
rect 308382 498838 325826 499074
rect 326062 498838 326146 499074
rect 326382 498838 343826 499074
rect 344062 498838 344146 499074
rect 344382 498838 361826 499074
rect 362062 498838 362146 499074
rect 362382 498838 379826 499074
rect 380062 498838 380146 499074
rect 380382 498838 397826 499074
rect 398062 498838 398146 499074
rect 398382 498838 415826 499074
rect 416062 498838 416146 499074
rect 416382 498838 433826 499074
rect 434062 498838 434146 499074
rect 434382 498838 451826 499074
rect 452062 498838 452146 499074
rect 452382 498838 469826 499074
rect 470062 498838 470146 499074
rect 470382 498838 487826 499074
rect 488062 498838 488146 499074
rect 488382 498838 505826 499074
rect 506062 498838 506146 499074
rect 506382 498838 523826 499074
rect 524062 498838 524146 499074
rect 524382 498838 541826 499074
rect 542062 498838 542146 499074
rect 542382 498838 542414 499074
rect 19794 498806 542414 498838
rect -2966 498454 586890 498486
rect -2966 498218 -2934 498454
rect -2698 498218 -2614 498454
rect -2378 498218 10826 498454
rect 11062 498218 11146 498454
rect 11382 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 46826 498454
rect 47062 498218 47146 498454
rect 47382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 82826 498454
rect 83062 498218 83146 498454
rect 83382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 118826 498454
rect 119062 498218 119146 498454
rect 119382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 154826 498454
rect 155062 498218 155146 498454
rect 155382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 190826 498454
rect 191062 498218 191146 498454
rect 191382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 226826 498454
rect 227062 498218 227146 498454
rect 227382 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 262826 498454
rect 263062 498218 263146 498454
rect 263382 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 298826 498454
rect 299062 498218 299146 498454
rect 299382 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 334826 498454
rect 335062 498218 335146 498454
rect 335382 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 370826 498454
rect 371062 498218 371146 498454
rect 371382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 406826 498454
rect 407062 498218 407146 498454
rect 407382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 442826 498454
rect 443062 498218 443146 498454
rect 443382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 478826 498454
rect 479062 498218 479146 498454
rect 479382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 514826 498454
rect 515062 498218 515146 498454
rect 515382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 550826 498454
rect 551062 498218 551146 498454
rect 551382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 586302 498454
rect 586538 498218 586622 498454
rect 586858 498218 586890 498454
rect -2966 498134 586890 498218
rect -2966 497898 -2934 498134
rect -2698 497898 -2614 498134
rect -2378 497898 10826 498134
rect 11062 497898 11146 498134
rect 11382 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 46826 498134
rect 47062 497898 47146 498134
rect 47382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 82826 498134
rect 83062 497898 83146 498134
rect 83382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 118826 498134
rect 119062 497898 119146 498134
rect 119382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 154826 498134
rect 155062 497898 155146 498134
rect 155382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 190826 498134
rect 191062 497898 191146 498134
rect 191382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 226826 498134
rect 227062 497898 227146 498134
rect 227382 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 262826 498134
rect 263062 497898 263146 498134
rect 263382 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 298826 498134
rect 299062 497898 299146 498134
rect 299382 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 334826 498134
rect 335062 497898 335146 498134
rect 335382 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 370826 498134
rect 371062 497898 371146 498134
rect 371382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 406826 498134
rect 407062 497898 407146 498134
rect 407382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 442826 498134
rect 443062 497898 443146 498134
rect 443382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 478826 498134
rect 479062 497898 479146 498134
rect 479382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 514826 498134
rect 515062 497898 515146 498134
rect 515382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 550826 498134
rect 551062 497898 551146 498134
rect 551382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 586302 498134
rect 586538 497898 586622 498134
rect 586858 497898 586890 498134
rect -2966 497866 586890 497898
rect -2966 489454 586890 489486
rect -2966 489218 -1974 489454
rect -1738 489218 -1654 489454
rect -1418 489218 1826 489454
rect 2062 489218 2146 489454
rect 2382 489218 19952 489454
rect 20188 489218 25882 489454
rect 26118 489218 31813 489454
rect 32049 489218 46952 489454
rect 47188 489218 52882 489454
rect 53118 489218 58813 489454
rect 59049 489218 73952 489454
rect 74188 489218 79882 489454
rect 80118 489218 85813 489454
rect 86049 489218 100952 489454
rect 101188 489218 106882 489454
rect 107118 489218 112813 489454
rect 113049 489218 127952 489454
rect 128188 489218 133882 489454
rect 134118 489218 139813 489454
rect 140049 489218 154952 489454
rect 155188 489218 160882 489454
rect 161118 489218 166813 489454
rect 167049 489218 181952 489454
rect 182188 489218 187882 489454
rect 188118 489218 193813 489454
rect 194049 489218 208952 489454
rect 209188 489218 214882 489454
rect 215118 489218 220813 489454
rect 221049 489218 235952 489454
rect 236188 489218 241882 489454
rect 242118 489218 247813 489454
rect 248049 489218 262952 489454
rect 263188 489218 268882 489454
rect 269118 489218 274813 489454
rect 275049 489218 289952 489454
rect 290188 489218 295882 489454
rect 296118 489218 301813 489454
rect 302049 489218 316952 489454
rect 317188 489218 322882 489454
rect 323118 489218 328813 489454
rect 329049 489218 343952 489454
rect 344188 489218 349882 489454
rect 350118 489218 355813 489454
rect 356049 489218 370952 489454
rect 371188 489218 376882 489454
rect 377118 489218 382813 489454
rect 383049 489218 397952 489454
rect 398188 489218 403882 489454
rect 404118 489218 409813 489454
rect 410049 489218 424952 489454
rect 425188 489218 430882 489454
rect 431118 489218 436813 489454
rect 437049 489218 451952 489454
rect 452188 489218 457882 489454
rect 458118 489218 463813 489454
rect 464049 489218 478952 489454
rect 479188 489218 484882 489454
rect 485118 489218 490813 489454
rect 491049 489218 505952 489454
rect 506188 489218 511882 489454
rect 512118 489218 517813 489454
rect 518049 489218 532952 489454
rect 533188 489218 538882 489454
rect 539118 489218 544813 489454
rect 545049 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 577826 489454
rect 578062 489218 578146 489454
rect 578382 489218 585342 489454
rect 585578 489218 585662 489454
rect 585898 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -1974 489134
rect -1738 488898 -1654 489134
rect -1418 488898 1826 489134
rect 2062 488898 2146 489134
rect 2382 488898 19952 489134
rect 20188 488898 25882 489134
rect 26118 488898 31813 489134
rect 32049 488898 46952 489134
rect 47188 488898 52882 489134
rect 53118 488898 58813 489134
rect 59049 488898 73952 489134
rect 74188 488898 79882 489134
rect 80118 488898 85813 489134
rect 86049 488898 100952 489134
rect 101188 488898 106882 489134
rect 107118 488898 112813 489134
rect 113049 488898 127952 489134
rect 128188 488898 133882 489134
rect 134118 488898 139813 489134
rect 140049 488898 154952 489134
rect 155188 488898 160882 489134
rect 161118 488898 166813 489134
rect 167049 488898 181952 489134
rect 182188 488898 187882 489134
rect 188118 488898 193813 489134
rect 194049 488898 208952 489134
rect 209188 488898 214882 489134
rect 215118 488898 220813 489134
rect 221049 488898 235952 489134
rect 236188 488898 241882 489134
rect 242118 488898 247813 489134
rect 248049 488898 262952 489134
rect 263188 488898 268882 489134
rect 269118 488898 274813 489134
rect 275049 488898 289952 489134
rect 290188 488898 295882 489134
rect 296118 488898 301813 489134
rect 302049 488898 316952 489134
rect 317188 488898 322882 489134
rect 323118 488898 328813 489134
rect 329049 488898 343952 489134
rect 344188 488898 349882 489134
rect 350118 488898 355813 489134
rect 356049 488898 370952 489134
rect 371188 488898 376882 489134
rect 377118 488898 382813 489134
rect 383049 488898 397952 489134
rect 398188 488898 403882 489134
rect 404118 488898 409813 489134
rect 410049 488898 424952 489134
rect 425188 488898 430882 489134
rect 431118 488898 436813 489134
rect 437049 488898 451952 489134
rect 452188 488898 457882 489134
rect 458118 488898 463813 489134
rect 464049 488898 478952 489134
rect 479188 488898 484882 489134
rect 485118 488898 490813 489134
rect 491049 488898 505952 489134
rect 506188 488898 511882 489134
rect 512118 488898 517813 489134
rect 518049 488898 532952 489134
rect 533188 488898 538882 489134
rect 539118 488898 544813 489134
rect 545049 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 577826 489134
rect 578062 488898 578146 489134
rect 578382 488898 585342 489134
rect 585578 488898 585662 489134
rect 585898 488898 586890 489134
rect -2966 488866 586890 488898
rect -2966 480454 586890 480486
rect -2966 480218 -2934 480454
rect -2698 480218 -2614 480454
rect -2378 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 22916 480454
rect 23152 480218 28847 480454
rect 29083 480218 49916 480454
rect 50152 480218 55847 480454
rect 56083 480218 76916 480454
rect 77152 480218 82847 480454
rect 83083 480218 103916 480454
rect 104152 480218 109847 480454
rect 110083 480218 130916 480454
rect 131152 480218 136847 480454
rect 137083 480218 157916 480454
rect 158152 480218 163847 480454
rect 164083 480218 184916 480454
rect 185152 480218 190847 480454
rect 191083 480218 211916 480454
rect 212152 480218 217847 480454
rect 218083 480218 238916 480454
rect 239152 480218 244847 480454
rect 245083 480218 265916 480454
rect 266152 480218 271847 480454
rect 272083 480218 292916 480454
rect 293152 480218 298847 480454
rect 299083 480218 319916 480454
rect 320152 480218 325847 480454
rect 326083 480218 346916 480454
rect 347152 480218 352847 480454
rect 353083 480218 373916 480454
rect 374152 480218 379847 480454
rect 380083 480218 400916 480454
rect 401152 480218 406847 480454
rect 407083 480218 427916 480454
rect 428152 480218 433847 480454
rect 434083 480218 454916 480454
rect 455152 480218 460847 480454
rect 461083 480218 481916 480454
rect 482152 480218 487847 480454
rect 488083 480218 508916 480454
rect 509152 480218 514847 480454
rect 515083 480218 535916 480454
rect 536152 480218 541847 480454
rect 542083 480218 568826 480454
rect 569062 480218 569146 480454
rect 569382 480218 586302 480454
rect 586538 480218 586622 480454
rect 586858 480218 586890 480454
rect -2966 480134 586890 480218
rect -2966 479898 -2934 480134
rect -2698 479898 -2614 480134
rect -2378 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 22916 480134
rect 23152 479898 28847 480134
rect 29083 479898 49916 480134
rect 50152 479898 55847 480134
rect 56083 479898 76916 480134
rect 77152 479898 82847 480134
rect 83083 479898 103916 480134
rect 104152 479898 109847 480134
rect 110083 479898 130916 480134
rect 131152 479898 136847 480134
rect 137083 479898 157916 480134
rect 158152 479898 163847 480134
rect 164083 479898 184916 480134
rect 185152 479898 190847 480134
rect 191083 479898 211916 480134
rect 212152 479898 217847 480134
rect 218083 479898 238916 480134
rect 239152 479898 244847 480134
rect 245083 479898 265916 480134
rect 266152 479898 271847 480134
rect 272083 479898 292916 480134
rect 293152 479898 298847 480134
rect 299083 479898 319916 480134
rect 320152 479898 325847 480134
rect 326083 479898 346916 480134
rect 347152 479898 352847 480134
rect 353083 479898 373916 480134
rect 374152 479898 379847 480134
rect 380083 479898 400916 480134
rect 401152 479898 406847 480134
rect 407083 479898 427916 480134
rect 428152 479898 433847 480134
rect 434083 479898 454916 480134
rect 455152 479898 460847 480134
rect 461083 479898 481916 480134
rect 482152 479898 487847 480134
rect 488083 479898 508916 480134
rect 509152 479898 514847 480134
rect 515083 479898 535916 480134
rect 536152 479898 541847 480134
rect 542083 479898 568826 480134
rect 569062 479898 569146 480134
rect 569382 479898 586302 480134
rect 586538 479898 586622 480134
rect 586858 479898 586890 480134
rect -2966 479866 586890 479898
rect 28794 472394 551414 472426
rect 28794 472158 28826 472394
rect 29062 472158 29146 472394
rect 29382 472158 46826 472394
rect 47062 472158 47146 472394
rect 47382 472158 64826 472394
rect 65062 472158 65146 472394
rect 65382 472158 82826 472394
rect 83062 472158 83146 472394
rect 83382 472158 100826 472394
rect 101062 472158 101146 472394
rect 101382 472158 118826 472394
rect 119062 472158 119146 472394
rect 119382 472158 136826 472394
rect 137062 472158 137146 472394
rect 137382 472158 154826 472394
rect 155062 472158 155146 472394
rect 155382 472158 172826 472394
rect 173062 472158 173146 472394
rect 173382 472158 190826 472394
rect 191062 472158 191146 472394
rect 191382 472158 208826 472394
rect 209062 472158 209146 472394
rect 209382 472158 226826 472394
rect 227062 472158 227146 472394
rect 227382 472158 244826 472394
rect 245062 472158 245146 472394
rect 245382 472158 262826 472394
rect 263062 472158 263146 472394
rect 263382 472158 280826 472394
rect 281062 472158 281146 472394
rect 281382 472158 298826 472394
rect 299062 472158 299146 472394
rect 299382 472158 316826 472394
rect 317062 472158 317146 472394
rect 317382 472158 334826 472394
rect 335062 472158 335146 472394
rect 335382 472158 352826 472394
rect 353062 472158 353146 472394
rect 353382 472158 370826 472394
rect 371062 472158 371146 472394
rect 371382 472158 388826 472394
rect 389062 472158 389146 472394
rect 389382 472158 406826 472394
rect 407062 472158 407146 472394
rect 407382 472158 424826 472394
rect 425062 472158 425146 472394
rect 425382 472158 442826 472394
rect 443062 472158 443146 472394
rect 443382 472158 460826 472394
rect 461062 472158 461146 472394
rect 461382 472158 478826 472394
rect 479062 472158 479146 472394
rect 479382 472158 496826 472394
rect 497062 472158 497146 472394
rect 497382 472158 514826 472394
rect 515062 472158 515146 472394
rect 515382 472158 532826 472394
rect 533062 472158 533146 472394
rect 533382 472158 550826 472394
rect 551062 472158 551146 472394
rect 551382 472158 551414 472394
rect 28794 472074 551414 472158
rect 28794 471838 28826 472074
rect 29062 471838 29146 472074
rect 29382 471838 46826 472074
rect 47062 471838 47146 472074
rect 47382 471838 64826 472074
rect 65062 471838 65146 472074
rect 65382 471838 82826 472074
rect 83062 471838 83146 472074
rect 83382 471838 100826 472074
rect 101062 471838 101146 472074
rect 101382 471838 118826 472074
rect 119062 471838 119146 472074
rect 119382 471838 136826 472074
rect 137062 471838 137146 472074
rect 137382 471838 154826 472074
rect 155062 471838 155146 472074
rect 155382 471838 172826 472074
rect 173062 471838 173146 472074
rect 173382 471838 190826 472074
rect 191062 471838 191146 472074
rect 191382 471838 208826 472074
rect 209062 471838 209146 472074
rect 209382 471838 226826 472074
rect 227062 471838 227146 472074
rect 227382 471838 244826 472074
rect 245062 471838 245146 472074
rect 245382 471838 262826 472074
rect 263062 471838 263146 472074
rect 263382 471838 280826 472074
rect 281062 471838 281146 472074
rect 281382 471838 298826 472074
rect 299062 471838 299146 472074
rect 299382 471838 316826 472074
rect 317062 471838 317146 472074
rect 317382 471838 334826 472074
rect 335062 471838 335146 472074
rect 335382 471838 352826 472074
rect 353062 471838 353146 472074
rect 353382 471838 370826 472074
rect 371062 471838 371146 472074
rect 371382 471838 388826 472074
rect 389062 471838 389146 472074
rect 389382 471838 406826 472074
rect 407062 471838 407146 472074
rect 407382 471838 424826 472074
rect 425062 471838 425146 472074
rect 425382 471838 442826 472074
rect 443062 471838 443146 472074
rect 443382 471838 460826 472074
rect 461062 471838 461146 472074
rect 461382 471838 478826 472074
rect 479062 471838 479146 472074
rect 479382 471838 496826 472074
rect 497062 471838 497146 472074
rect 497382 471838 514826 472074
rect 515062 471838 515146 472074
rect 515382 471838 532826 472074
rect 533062 471838 533146 472074
rect 533382 471838 550826 472074
rect 551062 471838 551146 472074
rect 551382 471838 551414 472074
rect 28794 471806 551414 471838
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 19826 471454
rect 20062 471218 20146 471454
rect 20382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 55826 471454
rect 56062 471218 56146 471454
rect 56382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 91826 471454
rect 92062 471218 92146 471454
rect 92382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 127826 471454
rect 128062 471218 128146 471454
rect 128382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 163826 471454
rect 164062 471218 164146 471454
rect 164382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 199826 471454
rect 200062 471218 200146 471454
rect 200382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 235826 471454
rect 236062 471218 236146 471454
rect 236382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 271826 471454
rect 272062 471218 272146 471454
rect 272382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 307826 471454
rect 308062 471218 308146 471454
rect 308382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 343826 471454
rect 344062 471218 344146 471454
rect 344382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 379826 471454
rect 380062 471218 380146 471454
rect 380382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 415826 471454
rect 416062 471218 416146 471454
rect 416382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 451826 471454
rect 452062 471218 452146 471454
rect 452382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 487826 471454
rect 488062 471218 488146 471454
rect 488382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 523826 471454
rect 524062 471218 524146 471454
rect 524382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 559826 471454
rect 560062 471218 560146 471454
rect 560382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 19826 471134
rect 20062 470898 20146 471134
rect 20382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 55826 471134
rect 56062 470898 56146 471134
rect 56382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 91826 471134
rect 92062 470898 92146 471134
rect 92382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 127826 471134
rect 128062 470898 128146 471134
rect 128382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 163826 471134
rect 164062 470898 164146 471134
rect 164382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 199826 471134
rect 200062 470898 200146 471134
rect 200382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 235826 471134
rect 236062 470898 236146 471134
rect 236382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 271826 471134
rect 272062 470898 272146 471134
rect 272382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 307826 471134
rect 308062 470898 308146 471134
rect 308382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 343826 471134
rect 344062 470898 344146 471134
rect 344382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 379826 471134
rect 380062 470898 380146 471134
rect 380382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 415826 471134
rect 416062 470898 416146 471134
rect 416382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 451826 471134
rect 452062 470898 452146 471134
rect 452382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 487826 471134
rect 488062 470898 488146 471134
rect 488382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 523826 471134
rect 524062 470898 524146 471134
rect 524382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 559826 471134
rect 560062 470898 560146 471134
rect 560382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -2966 462454 586890 462486
rect -2966 462218 -2934 462454
rect -2698 462218 -2614 462454
rect -2378 462218 10826 462454
rect 11062 462218 11146 462454
rect 11382 462218 22916 462454
rect 23152 462218 28847 462454
rect 29083 462218 49916 462454
rect 50152 462218 55847 462454
rect 56083 462218 76916 462454
rect 77152 462218 82847 462454
rect 83083 462218 103916 462454
rect 104152 462218 109847 462454
rect 110083 462218 130916 462454
rect 131152 462218 136847 462454
rect 137083 462218 157916 462454
rect 158152 462218 163847 462454
rect 164083 462218 184916 462454
rect 185152 462218 190847 462454
rect 191083 462218 211916 462454
rect 212152 462218 217847 462454
rect 218083 462218 238916 462454
rect 239152 462218 244847 462454
rect 245083 462218 265916 462454
rect 266152 462218 271847 462454
rect 272083 462218 292916 462454
rect 293152 462218 298847 462454
rect 299083 462218 319916 462454
rect 320152 462218 325847 462454
rect 326083 462218 346916 462454
rect 347152 462218 352847 462454
rect 353083 462218 373916 462454
rect 374152 462218 379847 462454
rect 380083 462218 400916 462454
rect 401152 462218 406847 462454
rect 407083 462218 427916 462454
rect 428152 462218 433847 462454
rect 434083 462218 454916 462454
rect 455152 462218 460847 462454
rect 461083 462218 481916 462454
rect 482152 462218 487847 462454
rect 488083 462218 508916 462454
rect 509152 462218 514847 462454
rect 515083 462218 535916 462454
rect 536152 462218 541847 462454
rect 542083 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 586302 462454
rect 586538 462218 586622 462454
rect 586858 462218 586890 462454
rect -2966 462134 586890 462218
rect -2966 461898 -2934 462134
rect -2698 461898 -2614 462134
rect -2378 461898 10826 462134
rect 11062 461898 11146 462134
rect 11382 461898 22916 462134
rect 23152 461898 28847 462134
rect 29083 461898 49916 462134
rect 50152 461898 55847 462134
rect 56083 461898 76916 462134
rect 77152 461898 82847 462134
rect 83083 461898 103916 462134
rect 104152 461898 109847 462134
rect 110083 461898 130916 462134
rect 131152 461898 136847 462134
rect 137083 461898 157916 462134
rect 158152 461898 163847 462134
rect 164083 461898 184916 462134
rect 185152 461898 190847 462134
rect 191083 461898 211916 462134
rect 212152 461898 217847 462134
rect 218083 461898 238916 462134
rect 239152 461898 244847 462134
rect 245083 461898 265916 462134
rect 266152 461898 271847 462134
rect 272083 461898 292916 462134
rect 293152 461898 298847 462134
rect 299083 461898 319916 462134
rect 320152 461898 325847 462134
rect 326083 461898 346916 462134
rect 347152 461898 352847 462134
rect 353083 461898 373916 462134
rect 374152 461898 379847 462134
rect 380083 461898 400916 462134
rect 401152 461898 406847 462134
rect 407083 461898 427916 462134
rect 428152 461898 433847 462134
rect 434083 461898 454916 462134
rect 455152 461898 460847 462134
rect 461083 461898 481916 462134
rect 482152 461898 487847 462134
rect 488083 461898 508916 462134
rect 509152 461898 514847 462134
rect 515083 461898 535916 462134
rect 536152 461898 541847 462134
rect 542083 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 586302 462134
rect 586538 461898 586622 462134
rect 586858 461898 586890 462134
rect -2966 461866 586890 461898
rect -2966 453454 586890 453486
rect -2966 453218 -1974 453454
rect -1738 453218 -1654 453454
rect -1418 453218 1826 453454
rect 2062 453218 2146 453454
rect 2382 453218 19952 453454
rect 20188 453218 25882 453454
rect 26118 453218 31813 453454
rect 32049 453218 46952 453454
rect 47188 453218 52882 453454
rect 53118 453218 58813 453454
rect 59049 453218 73952 453454
rect 74188 453218 79882 453454
rect 80118 453218 85813 453454
rect 86049 453218 100952 453454
rect 101188 453218 106882 453454
rect 107118 453218 112813 453454
rect 113049 453218 127952 453454
rect 128188 453218 133882 453454
rect 134118 453218 139813 453454
rect 140049 453218 154952 453454
rect 155188 453218 160882 453454
rect 161118 453218 166813 453454
rect 167049 453218 181952 453454
rect 182188 453218 187882 453454
rect 188118 453218 193813 453454
rect 194049 453218 208952 453454
rect 209188 453218 214882 453454
rect 215118 453218 220813 453454
rect 221049 453218 235952 453454
rect 236188 453218 241882 453454
rect 242118 453218 247813 453454
rect 248049 453218 262952 453454
rect 263188 453218 268882 453454
rect 269118 453218 274813 453454
rect 275049 453218 289952 453454
rect 290188 453218 295882 453454
rect 296118 453218 301813 453454
rect 302049 453218 316952 453454
rect 317188 453218 322882 453454
rect 323118 453218 328813 453454
rect 329049 453218 343952 453454
rect 344188 453218 349882 453454
rect 350118 453218 355813 453454
rect 356049 453218 370952 453454
rect 371188 453218 376882 453454
rect 377118 453218 382813 453454
rect 383049 453218 397952 453454
rect 398188 453218 403882 453454
rect 404118 453218 409813 453454
rect 410049 453218 424952 453454
rect 425188 453218 430882 453454
rect 431118 453218 436813 453454
rect 437049 453218 451952 453454
rect 452188 453218 457882 453454
rect 458118 453218 463813 453454
rect 464049 453218 478952 453454
rect 479188 453218 484882 453454
rect 485118 453218 490813 453454
rect 491049 453218 505952 453454
rect 506188 453218 511882 453454
rect 512118 453218 517813 453454
rect 518049 453218 532952 453454
rect 533188 453218 538882 453454
rect 539118 453218 544813 453454
rect 545049 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 577826 453454
rect 578062 453218 578146 453454
rect 578382 453218 585342 453454
rect 585578 453218 585662 453454
rect 585898 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -1974 453134
rect -1738 452898 -1654 453134
rect -1418 452898 1826 453134
rect 2062 452898 2146 453134
rect 2382 452898 19952 453134
rect 20188 452898 25882 453134
rect 26118 452898 31813 453134
rect 32049 452898 46952 453134
rect 47188 452898 52882 453134
rect 53118 452898 58813 453134
rect 59049 452898 73952 453134
rect 74188 452898 79882 453134
rect 80118 452898 85813 453134
rect 86049 452898 100952 453134
rect 101188 452898 106882 453134
rect 107118 452898 112813 453134
rect 113049 452898 127952 453134
rect 128188 452898 133882 453134
rect 134118 452898 139813 453134
rect 140049 452898 154952 453134
rect 155188 452898 160882 453134
rect 161118 452898 166813 453134
rect 167049 452898 181952 453134
rect 182188 452898 187882 453134
rect 188118 452898 193813 453134
rect 194049 452898 208952 453134
rect 209188 452898 214882 453134
rect 215118 452898 220813 453134
rect 221049 452898 235952 453134
rect 236188 452898 241882 453134
rect 242118 452898 247813 453134
rect 248049 452898 262952 453134
rect 263188 452898 268882 453134
rect 269118 452898 274813 453134
rect 275049 452898 289952 453134
rect 290188 452898 295882 453134
rect 296118 452898 301813 453134
rect 302049 452898 316952 453134
rect 317188 452898 322882 453134
rect 323118 452898 328813 453134
rect 329049 452898 343952 453134
rect 344188 452898 349882 453134
rect 350118 452898 355813 453134
rect 356049 452898 370952 453134
rect 371188 452898 376882 453134
rect 377118 452898 382813 453134
rect 383049 452898 397952 453134
rect 398188 452898 403882 453134
rect 404118 452898 409813 453134
rect 410049 452898 424952 453134
rect 425188 452898 430882 453134
rect 431118 452898 436813 453134
rect 437049 452898 451952 453134
rect 452188 452898 457882 453134
rect 458118 452898 463813 453134
rect 464049 452898 478952 453134
rect 479188 452898 484882 453134
rect 485118 452898 490813 453134
rect 491049 452898 505952 453134
rect 506188 452898 511882 453134
rect 512118 452898 517813 453134
rect 518049 452898 532952 453134
rect 533188 452898 538882 453134
rect 539118 452898 544813 453134
rect 545049 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 577826 453134
rect 578062 452898 578146 453134
rect 578382 452898 585342 453134
rect 585578 452898 585662 453134
rect 585898 452898 586890 453134
rect -2966 452866 586890 452898
rect 19794 445394 542414 445426
rect 19794 445158 19826 445394
rect 20062 445158 20146 445394
rect 20382 445158 37826 445394
rect 38062 445158 38146 445394
rect 38382 445158 55826 445394
rect 56062 445158 56146 445394
rect 56382 445158 73826 445394
rect 74062 445158 74146 445394
rect 74382 445158 91826 445394
rect 92062 445158 92146 445394
rect 92382 445158 109826 445394
rect 110062 445158 110146 445394
rect 110382 445158 127826 445394
rect 128062 445158 128146 445394
rect 128382 445158 145826 445394
rect 146062 445158 146146 445394
rect 146382 445158 163826 445394
rect 164062 445158 164146 445394
rect 164382 445158 181826 445394
rect 182062 445158 182146 445394
rect 182382 445158 199826 445394
rect 200062 445158 200146 445394
rect 200382 445158 217826 445394
rect 218062 445158 218146 445394
rect 218382 445158 235826 445394
rect 236062 445158 236146 445394
rect 236382 445158 253826 445394
rect 254062 445158 254146 445394
rect 254382 445158 271826 445394
rect 272062 445158 272146 445394
rect 272382 445158 289826 445394
rect 290062 445158 290146 445394
rect 290382 445158 307826 445394
rect 308062 445158 308146 445394
rect 308382 445158 325826 445394
rect 326062 445158 326146 445394
rect 326382 445158 343826 445394
rect 344062 445158 344146 445394
rect 344382 445158 361826 445394
rect 362062 445158 362146 445394
rect 362382 445158 379826 445394
rect 380062 445158 380146 445394
rect 380382 445158 397826 445394
rect 398062 445158 398146 445394
rect 398382 445158 415826 445394
rect 416062 445158 416146 445394
rect 416382 445158 433826 445394
rect 434062 445158 434146 445394
rect 434382 445158 451826 445394
rect 452062 445158 452146 445394
rect 452382 445158 469826 445394
rect 470062 445158 470146 445394
rect 470382 445158 487826 445394
rect 488062 445158 488146 445394
rect 488382 445158 505826 445394
rect 506062 445158 506146 445394
rect 506382 445158 523826 445394
rect 524062 445158 524146 445394
rect 524382 445158 541826 445394
rect 542062 445158 542146 445394
rect 542382 445158 542414 445394
rect 19794 445074 542414 445158
rect 19794 444838 19826 445074
rect 20062 444838 20146 445074
rect 20382 444838 37826 445074
rect 38062 444838 38146 445074
rect 38382 444838 55826 445074
rect 56062 444838 56146 445074
rect 56382 444838 73826 445074
rect 74062 444838 74146 445074
rect 74382 444838 91826 445074
rect 92062 444838 92146 445074
rect 92382 444838 109826 445074
rect 110062 444838 110146 445074
rect 110382 444838 127826 445074
rect 128062 444838 128146 445074
rect 128382 444838 145826 445074
rect 146062 444838 146146 445074
rect 146382 444838 163826 445074
rect 164062 444838 164146 445074
rect 164382 444838 181826 445074
rect 182062 444838 182146 445074
rect 182382 444838 199826 445074
rect 200062 444838 200146 445074
rect 200382 444838 217826 445074
rect 218062 444838 218146 445074
rect 218382 444838 235826 445074
rect 236062 444838 236146 445074
rect 236382 444838 253826 445074
rect 254062 444838 254146 445074
rect 254382 444838 271826 445074
rect 272062 444838 272146 445074
rect 272382 444838 289826 445074
rect 290062 444838 290146 445074
rect 290382 444838 307826 445074
rect 308062 444838 308146 445074
rect 308382 444838 325826 445074
rect 326062 444838 326146 445074
rect 326382 444838 343826 445074
rect 344062 444838 344146 445074
rect 344382 444838 361826 445074
rect 362062 444838 362146 445074
rect 362382 444838 379826 445074
rect 380062 444838 380146 445074
rect 380382 444838 397826 445074
rect 398062 444838 398146 445074
rect 398382 444838 415826 445074
rect 416062 444838 416146 445074
rect 416382 444838 433826 445074
rect 434062 444838 434146 445074
rect 434382 444838 451826 445074
rect 452062 444838 452146 445074
rect 452382 444838 469826 445074
rect 470062 444838 470146 445074
rect 470382 444838 487826 445074
rect 488062 444838 488146 445074
rect 488382 444838 505826 445074
rect 506062 444838 506146 445074
rect 506382 444838 523826 445074
rect 524062 444838 524146 445074
rect 524382 444838 541826 445074
rect 542062 444838 542146 445074
rect 542382 444838 542414 445074
rect 19794 444806 542414 444838
rect -2966 444454 586890 444486
rect -2966 444218 -2934 444454
rect -2698 444218 -2614 444454
rect -2378 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 28826 444454
rect 29062 444218 29146 444454
rect 29382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 64826 444454
rect 65062 444218 65146 444454
rect 65382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 100826 444454
rect 101062 444218 101146 444454
rect 101382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 136826 444454
rect 137062 444218 137146 444454
rect 137382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 172826 444454
rect 173062 444218 173146 444454
rect 173382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 208826 444454
rect 209062 444218 209146 444454
rect 209382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 244826 444454
rect 245062 444218 245146 444454
rect 245382 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 280826 444454
rect 281062 444218 281146 444454
rect 281382 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 316826 444454
rect 317062 444218 317146 444454
rect 317382 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 352826 444454
rect 353062 444218 353146 444454
rect 353382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 388826 444454
rect 389062 444218 389146 444454
rect 389382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 424826 444454
rect 425062 444218 425146 444454
rect 425382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 460826 444454
rect 461062 444218 461146 444454
rect 461382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 496826 444454
rect 497062 444218 497146 444454
rect 497382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 532826 444454
rect 533062 444218 533146 444454
rect 533382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 568826 444454
rect 569062 444218 569146 444454
rect 569382 444218 586302 444454
rect 586538 444218 586622 444454
rect 586858 444218 586890 444454
rect -2966 444134 586890 444218
rect -2966 443898 -2934 444134
rect -2698 443898 -2614 444134
rect -2378 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 28826 444134
rect 29062 443898 29146 444134
rect 29382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 64826 444134
rect 65062 443898 65146 444134
rect 65382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 100826 444134
rect 101062 443898 101146 444134
rect 101382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 136826 444134
rect 137062 443898 137146 444134
rect 137382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 172826 444134
rect 173062 443898 173146 444134
rect 173382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 208826 444134
rect 209062 443898 209146 444134
rect 209382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 244826 444134
rect 245062 443898 245146 444134
rect 245382 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 280826 444134
rect 281062 443898 281146 444134
rect 281382 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 316826 444134
rect 317062 443898 317146 444134
rect 317382 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 352826 444134
rect 353062 443898 353146 444134
rect 353382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 388826 444134
rect 389062 443898 389146 444134
rect 389382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 424826 444134
rect 425062 443898 425146 444134
rect 425382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 460826 444134
rect 461062 443898 461146 444134
rect 461382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 496826 444134
rect 497062 443898 497146 444134
rect 497382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 532826 444134
rect 533062 443898 533146 444134
rect 533382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 568826 444134
rect 569062 443898 569146 444134
rect 569382 443898 586302 444134
rect 586538 443898 586622 444134
rect 586858 443898 586890 444134
rect -2966 443866 586890 443898
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 19952 435454
rect 20188 435218 25882 435454
rect 26118 435218 31813 435454
rect 32049 435218 46952 435454
rect 47188 435218 52882 435454
rect 53118 435218 58813 435454
rect 59049 435218 73952 435454
rect 74188 435218 79882 435454
rect 80118 435218 85813 435454
rect 86049 435218 100952 435454
rect 101188 435218 106882 435454
rect 107118 435218 112813 435454
rect 113049 435218 127952 435454
rect 128188 435218 133882 435454
rect 134118 435218 139813 435454
rect 140049 435218 154952 435454
rect 155188 435218 160882 435454
rect 161118 435218 166813 435454
rect 167049 435218 181952 435454
rect 182188 435218 187882 435454
rect 188118 435218 193813 435454
rect 194049 435218 208952 435454
rect 209188 435218 214882 435454
rect 215118 435218 220813 435454
rect 221049 435218 235952 435454
rect 236188 435218 241882 435454
rect 242118 435218 247813 435454
rect 248049 435218 262952 435454
rect 263188 435218 268882 435454
rect 269118 435218 274813 435454
rect 275049 435218 289952 435454
rect 290188 435218 295882 435454
rect 296118 435218 301813 435454
rect 302049 435218 316952 435454
rect 317188 435218 322882 435454
rect 323118 435218 328813 435454
rect 329049 435218 343952 435454
rect 344188 435218 349882 435454
rect 350118 435218 355813 435454
rect 356049 435218 370952 435454
rect 371188 435218 376882 435454
rect 377118 435218 382813 435454
rect 383049 435218 397952 435454
rect 398188 435218 403882 435454
rect 404118 435218 409813 435454
rect 410049 435218 424952 435454
rect 425188 435218 430882 435454
rect 431118 435218 436813 435454
rect 437049 435218 451952 435454
rect 452188 435218 457882 435454
rect 458118 435218 463813 435454
rect 464049 435218 478952 435454
rect 479188 435218 484882 435454
rect 485118 435218 490813 435454
rect 491049 435218 505952 435454
rect 506188 435218 511882 435454
rect 512118 435218 517813 435454
rect 518049 435218 532952 435454
rect 533188 435218 538882 435454
rect 539118 435218 544813 435454
rect 545049 435218 559826 435454
rect 560062 435218 560146 435454
rect 560382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 19952 435134
rect 20188 434898 25882 435134
rect 26118 434898 31813 435134
rect 32049 434898 46952 435134
rect 47188 434898 52882 435134
rect 53118 434898 58813 435134
rect 59049 434898 73952 435134
rect 74188 434898 79882 435134
rect 80118 434898 85813 435134
rect 86049 434898 100952 435134
rect 101188 434898 106882 435134
rect 107118 434898 112813 435134
rect 113049 434898 127952 435134
rect 128188 434898 133882 435134
rect 134118 434898 139813 435134
rect 140049 434898 154952 435134
rect 155188 434898 160882 435134
rect 161118 434898 166813 435134
rect 167049 434898 181952 435134
rect 182188 434898 187882 435134
rect 188118 434898 193813 435134
rect 194049 434898 208952 435134
rect 209188 434898 214882 435134
rect 215118 434898 220813 435134
rect 221049 434898 235952 435134
rect 236188 434898 241882 435134
rect 242118 434898 247813 435134
rect 248049 434898 262952 435134
rect 263188 434898 268882 435134
rect 269118 434898 274813 435134
rect 275049 434898 289952 435134
rect 290188 434898 295882 435134
rect 296118 434898 301813 435134
rect 302049 434898 316952 435134
rect 317188 434898 322882 435134
rect 323118 434898 328813 435134
rect 329049 434898 343952 435134
rect 344188 434898 349882 435134
rect 350118 434898 355813 435134
rect 356049 434898 370952 435134
rect 371188 434898 376882 435134
rect 377118 434898 382813 435134
rect 383049 434898 397952 435134
rect 398188 434898 403882 435134
rect 404118 434898 409813 435134
rect 410049 434898 424952 435134
rect 425188 434898 430882 435134
rect 431118 434898 436813 435134
rect 437049 434898 451952 435134
rect 452188 434898 457882 435134
rect 458118 434898 463813 435134
rect 464049 434898 478952 435134
rect 479188 434898 484882 435134
rect 485118 434898 490813 435134
rect 491049 434898 505952 435134
rect 506188 434898 511882 435134
rect 512118 434898 517813 435134
rect 518049 434898 532952 435134
rect 533188 434898 538882 435134
rect 539118 434898 544813 435134
rect 545049 434898 559826 435134
rect 560062 434898 560146 435134
rect 560382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -2966 426454 586890 426486
rect -2966 426218 -2934 426454
rect -2698 426218 -2614 426454
rect -2378 426218 10826 426454
rect 11062 426218 11146 426454
rect 11382 426218 22916 426454
rect 23152 426218 28847 426454
rect 29083 426218 49916 426454
rect 50152 426218 55847 426454
rect 56083 426218 76916 426454
rect 77152 426218 82847 426454
rect 83083 426218 103916 426454
rect 104152 426218 109847 426454
rect 110083 426218 130916 426454
rect 131152 426218 136847 426454
rect 137083 426218 157916 426454
rect 158152 426218 163847 426454
rect 164083 426218 184916 426454
rect 185152 426218 190847 426454
rect 191083 426218 211916 426454
rect 212152 426218 217847 426454
rect 218083 426218 238916 426454
rect 239152 426218 244847 426454
rect 245083 426218 265916 426454
rect 266152 426218 271847 426454
rect 272083 426218 292916 426454
rect 293152 426218 298847 426454
rect 299083 426218 319916 426454
rect 320152 426218 325847 426454
rect 326083 426218 346916 426454
rect 347152 426218 352847 426454
rect 353083 426218 373916 426454
rect 374152 426218 379847 426454
rect 380083 426218 400916 426454
rect 401152 426218 406847 426454
rect 407083 426218 427916 426454
rect 428152 426218 433847 426454
rect 434083 426218 454916 426454
rect 455152 426218 460847 426454
rect 461083 426218 481916 426454
rect 482152 426218 487847 426454
rect 488083 426218 508916 426454
rect 509152 426218 514847 426454
rect 515083 426218 535916 426454
rect 536152 426218 541847 426454
rect 542083 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 586302 426454
rect 586538 426218 586622 426454
rect 586858 426218 586890 426454
rect -2966 426134 586890 426218
rect -2966 425898 -2934 426134
rect -2698 425898 -2614 426134
rect -2378 425898 10826 426134
rect 11062 425898 11146 426134
rect 11382 425898 22916 426134
rect 23152 425898 28847 426134
rect 29083 425898 49916 426134
rect 50152 425898 55847 426134
rect 56083 425898 76916 426134
rect 77152 425898 82847 426134
rect 83083 425898 103916 426134
rect 104152 425898 109847 426134
rect 110083 425898 130916 426134
rect 131152 425898 136847 426134
rect 137083 425898 157916 426134
rect 158152 425898 163847 426134
rect 164083 425898 184916 426134
rect 185152 425898 190847 426134
rect 191083 425898 211916 426134
rect 212152 425898 217847 426134
rect 218083 425898 238916 426134
rect 239152 425898 244847 426134
rect 245083 425898 265916 426134
rect 266152 425898 271847 426134
rect 272083 425898 292916 426134
rect 293152 425898 298847 426134
rect 299083 425898 319916 426134
rect 320152 425898 325847 426134
rect 326083 425898 346916 426134
rect 347152 425898 352847 426134
rect 353083 425898 373916 426134
rect 374152 425898 379847 426134
rect 380083 425898 400916 426134
rect 401152 425898 406847 426134
rect 407083 425898 427916 426134
rect 428152 425898 433847 426134
rect 434083 425898 454916 426134
rect 455152 425898 460847 426134
rect 461083 425898 481916 426134
rect 482152 425898 487847 426134
rect 488083 425898 508916 426134
rect 509152 425898 514847 426134
rect 515083 425898 535916 426134
rect 536152 425898 541847 426134
rect 542083 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 586302 426134
rect 586538 425898 586622 426134
rect 586858 425898 586890 426134
rect -2966 425866 586890 425898
rect 28794 418394 551414 418426
rect 28794 418158 28826 418394
rect 29062 418158 29146 418394
rect 29382 418158 46826 418394
rect 47062 418158 47146 418394
rect 47382 418158 64826 418394
rect 65062 418158 65146 418394
rect 65382 418158 82826 418394
rect 83062 418158 83146 418394
rect 83382 418158 100826 418394
rect 101062 418158 101146 418394
rect 101382 418158 118826 418394
rect 119062 418158 119146 418394
rect 119382 418158 136826 418394
rect 137062 418158 137146 418394
rect 137382 418158 154826 418394
rect 155062 418158 155146 418394
rect 155382 418158 172826 418394
rect 173062 418158 173146 418394
rect 173382 418158 190826 418394
rect 191062 418158 191146 418394
rect 191382 418158 208826 418394
rect 209062 418158 209146 418394
rect 209382 418158 226826 418394
rect 227062 418158 227146 418394
rect 227382 418158 244826 418394
rect 245062 418158 245146 418394
rect 245382 418158 262826 418394
rect 263062 418158 263146 418394
rect 263382 418158 280826 418394
rect 281062 418158 281146 418394
rect 281382 418158 298826 418394
rect 299062 418158 299146 418394
rect 299382 418158 316826 418394
rect 317062 418158 317146 418394
rect 317382 418158 334826 418394
rect 335062 418158 335146 418394
rect 335382 418158 352826 418394
rect 353062 418158 353146 418394
rect 353382 418158 370826 418394
rect 371062 418158 371146 418394
rect 371382 418158 388826 418394
rect 389062 418158 389146 418394
rect 389382 418158 406826 418394
rect 407062 418158 407146 418394
rect 407382 418158 424826 418394
rect 425062 418158 425146 418394
rect 425382 418158 442826 418394
rect 443062 418158 443146 418394
rect 443382 418158 460826 418394
rect 461062 418158 461146 418394
rect 461382 418158 478826 418394
rect 479062 418158 479146 418394
rect 479382 418158 496826 418394
rect 497062 418158 497146 418394
rect 497382 418158 514826 418394
rect 515062 418158 515146 418394
rect 515382 418158 532826 418394
rect 533062 418158 533146 418394
rect 533382 418158 550826 418394
rect 551062 418158 551146 418394
rect 551382 418158 551414 418394
rect 28794 418074 551414 418158
rect 28794 417838 28826 418074
rect 29062 417838 29146 418074
rect 29382 417838 46826 418074
rect 47062 417838 47146 418074
rect 47382 417838 64826 418074
rect 65062 417838 65146 418074
rect 65382 417838 82826 418074
rect 83062 417838 83146 418074
rect 83382 417838 100826 418074
rect 101062 417838 101146 418074
rect 101382 417838 118826 418074
rect 119062 417838 119146 418074
rect 119382 417838 136826 418074
rect 137062 417838 137146 418074
rect 137382 417838 154826 418074
rect 155062 417838 155146 418074
rect 155382 417838 172826 418074
rect 173062 417838 173146 418074
rect 173382 417838 190826 418074
rect 191062 417838 191146 418074
rect 191382 417838 208826 418074
rect 209062 417838 209146 418074
rect 209382 417838 226826 418074
rect 227062 417838 227146 418074
rect 227382 417838 244826 418074
rect 245062 417838 245146 418074
rect 245382 417838 262826 418074
rect 263062 417838 263146 418074
rect 263382 417838 280826 418074
rect 281062 417838 281146 418074
rect 281382 417838 298826 418074
rect 299062 417838 299146 418074
rect 299382 417838 316826 418074
rect 317062 417838 317146 418074
rect 317382 417838 334826 418074
rect 335062 417838 335146 418074
rect 335382 417838 352826 418074
rect 353062 417838 353146 418074
rect 353382 417838 370826 418074
rect 371062 417838 371146 418074
rect 371382 417838 388826 418074
rect 389062 417838 389146 418074
rect 389382 417838 406826 418074
rect 407062 417838 407146 418074
rect 407382 417838 424826 418074
rect 425062 417838 425146 418074
rect 425382 417838 442826 418074
rect 443062 417838 443146 418074
rect 443382 417838 460826 418074
rect 461062 417838 461146 418074
rect 461382 417838 478826 418074
rect 479062 417838 479146 418074
rect 479382 417838 496826 418074
rect 497062 417838 497146 418074
rect 497382 417838 514826 418074
rect 515062 417838 515146 418074
rect 515382 417838 532826 418074
rect 533062 417838 533146 418074
rect 533382 417838 550826 418074
rect 551062 417838 551146 418074
rect 551382 417838 551414 418074
rect 28794 417806 551414 417838
rect -2966 417454 586890 417486
rect -2966 417218 -1974 417454
rect -1738 417218 -1654 417454
rect -1418 417218 1826 417454
rect 2062 417218 2146 417454
rect 2382 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 37826 417454
rect 38062 417218 38146 417454
rect 38382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 73826 417454
rect 74062 417218 74146 417454
rect 74382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 109826 417454
rect 110062 417218 110146 417454
rect 110382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 145826 417454
rect 146062 417218 146146 417454
rect 146382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 181826 417454
rect 182062 417218 182146 417454
rect 182382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 217826 417454
rect 218062 417218 218146 417454
rect 218382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 253826 417454
rect 254062 417218 254146 417454
rect 254382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 289826 417454
rect 290062 417218 290146 417454
rect 290382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 325826 417454
rect 326062 417218 326146 417454
rect 326382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 361826 417454
rect 362062 417218 362146 417454
rect 362382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 397826 417454
rect 398062 417218 398146 417454
rect 398382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 433826 417454
rect 434062 417218 434146 417454
rect 434382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 469826 417454
rect 470062 417218 470146 417454
rect 470382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 505826 417454
rect 506062 417218 506146 417454
rect 506382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 541826 417454
rect 542062 417218 542146 417454
rect 542382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 577826 417454
rect 578062 417218 578146 417454
rect 578382 417218 585342 417454
rect 585578 417218 585662 417454
rect 585898 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -1974 417134
rect -1738 416898 -1654 417134
rect -1418 416898 1826 417134
rect 2062 416898 2146 417134
rect 2382 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 37826 417134
rect 38062 416898 38146 417134
rect 38382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 73826 417134
rect 74062 416898 74146 417134
rect 74382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 109826 417134
rect 110062 416898 110146 417134
rect 110382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 145826 417134
rect 146062 416898 146146 417134
rect 146382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 181826 417134
rect 182062 416898 182146 417134
rect 182382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 217826 417134
rect 218062 416898 218146 417134
rect 218382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 253826 417134
rect 254062 416898 254146 417134
rect 254382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 289826 417134
rect 290062 416898 290146 417134
rect 290382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 325826 417134
rect 326062 416898 326146 417134
rect 326382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 361826 417134
rect 362062 416898 362146 417134
rect 362382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 397826 417134
rect 398062 416898 398146 417134
rect 398382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 433826 417134
rect 434062 416898 434146 417134
rect 434382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 469826 417134
rect 470062 416898 470146 417134
rect 470382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 505826 417134
rect 506062 416898 506146 417134
rect 506382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 541826 417134
rect 542062 416898 542146 417134
rect 542382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 577826 417134
rect 578062 416898 578146 417134
rect 578382 416898 585342 417134
rect 585578 416898 585662 417134
rect 585898 416898 586890 417134
rect -2966 416866 586890 416898
rect -2966 408454 586890 408486
rect -2966 408218 -2934 408454
rect -2698 408218 -2614 408454
rect -2378 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 22916 408454
rect 23152 408218 28847 408454
rect 29083 408218 49916 408454
rect 50152 408218 55847 408454
rect 56083 408218 76916 408454
rect 77152 408218 82847 408454
rect 83083 408218 103916 408454
rect 104152 408218 109847 408454
rect 110083 408218 130916 408454
rect 131152 408218 136847 408454
rect 137083 408218 157916 408454
rect 158152 408218 163847 408454
rect 164083 408218 184916 408454
rect 185152 408218 190847 408454
rect 191083 408218 211916 408454
rect 212152 408218 217847 408454
rect 218083 408218 238916 408454
rect 239152 408218 244847 408454
rect 245083 408218 265916 408454
rect 266152 408218 271847 408454
rect 272083 408218 292916 408454
rect 293152 408218 298847 408454
rect 299083 408218 319916 408454
rect 320152 408218 325847 408454
rect 326083 408218 346916 408454
rect 347152 408218 352847 408454
rect 353083 408218 373916 408454
rect 374152 408218 379847 408454
rect 380083 408218 400916 408454
rect 401152 408218 406847 408454
rect 407083 408218 427916 408454
rect 428152 408218 433847 408454
rect 434083 408218 454916 408454
rect 455152 408218 460847 408454
rect 461083 408218 481916 408454
rect 482152 408218 487847 408454
rect 488083 408218 508916 408454
rect 509152 408218 514847 408454
rect 515083 408218 535916 408454
rect 536152 408218 541847 408454
rect 542083 408218 568826 408454
rect 569062 408218 569146 408454
rect 569382 408218 586302 408454
rect 586538 408218 586622 408454
rect 586858 408218 586890 408454
rect -2966 408134 586890 408218
rect -2966 407898 -2934 408134
rect -2698 407898 -2614 408134
rect -2378 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 22916 408134
rect 23152 407898 28847 408134
rect 29083 407898 49916 408134
rect 50152 407898 55847 408134
rect 56083 407898 76916 408134
rect 77152 407898 82847 408134
rect 83083 407898 103916 408134
rect 104152 407898 109847 408134
rect 110083 407898 130916 408134
rect 131152 407898 136847 408134
rect 137083 407898 157916 408134
rect 158152 407898 163847 408134
rect 164083 407898 184916 408134
rect 185152 407898 190847 408134
rect 191083 407898 211916 408134
rect 212152 407898 217847 408134
rect 218083 407898 238916 408134
rect 239152 407898 244847 408134
rect 245083 407898 265916 408134
rect 266152 407898 271847 408134
rect 272083 407898 292916 408134
rect 293152 407898 298847 408134
rect 299083 407898 319916 408134
rect 320152 407898 325847 408134
rect 326083 407898 346916 408134
rect 347152 407898 352847 408134
rect 353083 407898 373916 408134
rect 374152 407898 379847 408134
rect 380083 407898 400916 408134
rect 401152 407898 406847 408134
rect 407083 407898 427916 408134
rect 428152 407898 433847 408134
rect 434083 407898 454916 408134
rect 455152 407898 460847 408134
rect 461083 407898 481916 408134
rect 482152 407898 487847 408134
rect 488083 407898 508916 408134
rect 509152 407898 514847 408134
rect 515083 407898 535916 408134
rect 536152 407898 541847 408134
rect 542083 407898 568826 408134
rect 569062 407898 569146 408134
rect 569382 407898 586302 408134
rect 586538 407898 586622 408134
rect 586858 407898 586890 408134
rect -2966 407866 586890 407898
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 19952 399454
rect 20188 399218 25882 399454
rect 26118 399218 31813 399454
rect 32049 399218 46952 399454
rect 47188 399218 52882 399454
rect 53118 399218 58813 399454
rect 59049 399218 73952 399454
rect 74188 399218 79882 399454
rect 80118 399218 85813 399454
rect 86049 399218 100952 399454
rect 101188 399218 106882 399454
rect 107118 399218 112813 399454
rect 113049 399218 127952 399454
rect 128188 399218 133882 399454
rect 134118 399218 139813 399454
rect 140049 399218 154952 399454
rect 155188 399218 160882 399454
rect 161118 399218 166813 399454
rect 167049 399218 181952 399454
rect 182188 399218 187882 399454
rect 188118 399218 193813 399454
rect 194049 399218 208952 399454
rect 209188 399218 214882 399454
rect 215118 399218 220813 399454
rect 221049 399218 235952 399454
rect 236188 399218 241882 399454
rect 242118 399218 247813 399454
rect 248049 399218 262952 399454
rect 263188 399218 268882 399454
rect 269118 399218 274813 399454
rect 275049 399218 289952 399454
rect 290188 399218 295882 399454
rect 296118 399218 301813 399454
rect 302049 399218 316952 399454
rect 317188 399218 322882 399454
rect 323118 399218 328813 399454
rect 329049 399218 343952 399454
rect 344188 399218 349882 399454
rect 350118 399218 355813 399454
rect 356049 399218 370952 399454
rect 371188 399218 376882 399454
rect 377118 399218 382813 399454
rect 383049 399218 397952 399454
rect 398188 399218 403882 399454
rect 404118 399218 409813 399454
rect 410049 399218 424952 399454
rect 425188 399218 430882 399454
rect 431118 399218 436813 399454
rect 437049 399218 451952 399454
rect 452188 399218 457882 399454
rect 458118 399218 463813 399454
rect 464049 399218 478952 399454
rect 479188 399218 484882 399454
rect 485118 399218 490813 399454
rect 491049 399218 505952 399454
rect 506188 399218 511882 399454
rect 512118 399218 517813 399454
rect 518049 399218 532952 399454
rect 533188 399218 538882 399454
rect 539118 399218 544813 399454
rect 545049 399218 559826 399454
rect 560062 399218 560146 399454
rect 560382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 19952 399134
rect 20188 398898 25882 399134
rect 26118 398898 31813 399134
rect 32049 398898 46952 399134
rect 47188 398898 52882 399134
rect 53118 398898 58813 399134
rect 59049 398898 73952 399134
rect 74188 398898 79882 399134
rect 80118 398898 85813 399134
rect 86049 398898 100952 399134
rect 101188 398898 106882 399134
rect 107118 398898 112813 399134
rect 113049 398898 127952 399134
rect 128188 398898 133882 399134
rect 134118 398898 139813 399134
rect 140049 398898 154952 399134
rect 155188 398898 160882 399134
rect 161118 398898 166813 399134
rect 167049 398898 181952 399134
rect 182188 398898 187882 399134
rect 188118 398898 193813 399134
rect 194049 398898 208952 399134
rect 209188 398898 214882 399134
rect 215118 398898 220813 399134
rect 221049 398898 235952 399134
rect 236188 398898 241882 399134
rect 242118 398898 247813 399134
rect 248049 398898 262952 399134
rect 263188 398898 268882 399134
rect 269118 398898 274813 399134
rect 275049 398898 289952 399134
rect 290188 398898 295882 399134
rect 296118 398898 301813 399134
rect 302049 398898 316952 399134
rect 317188 398898 322882 399134
rect 323118 398898 328813 399134
rect 329049 398898 343952 399134
rect 344188 398898 349882 399134
rect 350118 398898 355813 399134
rect 356049 398898 370952 399134
rect 371188 398898 376882 399134
rect 377118 398898 382813 399134
rect 383049 398898 397952 399134
rect 398188 398898 403882 399134
rect 404118 398898 409813 399134
rect 410049 398898 424952 399134
rect 425188 398898 430882 399134
rect 431118 398898 436813 399134
rect 437049 398898 451952 399134
rect 452188 398898 457882 399134
rect 458118 398898 463813 399134
rect 464049 398898 478952 399134
rect 479188 398898 484882 399134
rect 485118 398898 490813 399134
rect 491049 398898 505952 399134
rect 506188 398898 511882 399134
rect 512118 398898 517813 399134
rect 518049 398898 532952 399134
rect 533188 398898 538882 399134
rect 539118 398898 544813 399134
rect 545049 398898 559826 399134
rect 560062 398898 560146 399134
rect 560382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect 19794 391394 542414 391426
rect 19794 391158 19826 391394
rect 20062 391158 20146 391394
rect 20382 391158 37826 391394
rect 38062 391158 38146 391394
rect 38382 391158 55826 391394
rect 56062 391158 56146 391394
rect 56382 391158 73826 391394
rect 74062 391158 74146 391394
rect 74382 391158 91826 391394
rect 92062 391158 92146 391394
rect 92382 391158 109826 391394
rect 110062 391158 110146 391394
rect 110382 391158 127826 391394
rect 128062 391158 128146 391394
rect 128382 391158 145826 391394
rect 146062 391158 146146 391394
rect 146382 391158 163826 391394
rect 164062 391158 164146 391394
rect 164382 391158 181826 391394
rect 182062 391158 182146 391394
rect 182382 391158 199826 391394
rect 200062 391158 200146 391394
rect 200382 391158 217826 391394
rect 218062 391158 218146 391394
rect 218382 391158 235826 391394
rect 236062 391158 236146 391394
rect 236382 391158 253826 391394
rect 254062 391158 254146 391394
rect 254382 391158 271826 391394
rect 272062 391158 272146 391394
rect 272382 391158 289826 391394
rect 290062 391158 290146 391394
rect 290382 391158 307826 391394
rect 308062 391158 308146 391394
rect 308382 391158 325826 391394
rect 326062 391158 326146 391394
rect 326382 391158 343826 391394
rect 344062 391158 344146 391394
rect 344382 391158 361826 391394
rect 362062 391158 362146 391394
rect 362382 391158 379826 391394
rect 380062 391158 380146 391394
rect 380382 391158 397826 391394
rect 398062 391158 398146 391394
rect 398382 391158 415826 391394
rect 416062 391158 416146 391394
rect 416382 391158 433826 391394
rect 434062 391158 434146 391394
rect 434382 391158 451826 391394
rect 452062 391158 452146 391394
rect 452382 391158 469826 391394
rect 470062 391158 470146 391394
rect 470382 391158 487826 391394
rect 488062 391158 488146 391394
rect 488382 391158 505826 391394
rect 506062 391158 506146 391394
rect 506382 391158 523826 391394
rect 524062 391158 524146 391394
rect 524382 391158 541826 391394
rect 542062 391158 542146 391394
rect 542382 391158 542414 391394
rect 19794 391074 542414 391158
rect 19794 390838 19826 391074
rect 20062 390838 20146 391074
rect 20382 390838 37826 391074
rect 38062 390838 38146 391074
rect 38382 390838 55826 391074
rect 56062 390838 56146 391074
rect 56382 390838 73826 391074
rect 74062 390838 74146 391074
rect 74382 390838 91826 391074
rect 92062 390838 92146 391074
rect 92382 390838 109826 391074
rect 110062 390838 110146 391074
rect 110382 390838 127826 391074
rect 128062 390838 128146 391074
rect 128382 390838 145826 391074
rect 146062 390838 146146 391074
rect 146382 390838 163826 391074
rect 164062 390838 164146 391074
rect 164382 390838 181826 391074
rect 182062 390838 182146 391074
rect 182382 390838 199826 391074
rect 200062 390838 200146 391074
rect 200382 390838 217826 391074
rect 218062 390838 218146 391074
rect 218382 390838 235826 391074
rect 236062 390838 236146 391074
rect 236382 390838 253826 391074
rect 254062 390838 254146 391074
rect 254382 390838 271826 391074
rect 272062 390838 272146 391074
rect 272382 390838 289826 391074
rect 290062 390838 290146 391074
rect 290382 390838 307826 391074
rect 308062 390838 308146 391074
rect 308382 390838 325826 391074
rect 326062 390838 326146 391074
rect 326382 390838 343826 391074
rect 344062 390838 344146 391074
rect 344382 390838 361826 391074
rect 362062 390838 362146 391074
rect 362382 390838 379826 391074
rect 380062 390838 380146 391074
rect 380382 390838 397826 391074
rect 398062 390838 398146 391074
rect 398382 390838 415826 391074
rect 416062 390838 416146 391074
rect 416382 390838 433826 391074
rect 434062 390838 434146 391074
rect 434382 390838 451826 391074
rect 452062 390838 452146 391074
rect 452382 390838 469826 391074
rect 470062 390838 470146 391074
rect 470382 390838 487826 391074
rect 488062 390838 488146 391074
rect 488382 390838 505826 391074
rect 506062 390838 506146 391074
rect 506382 390838 523826 391074
rect 524062 390838 524146 391074
rect 524382 390838 541826 391074
rect 542062 390838 542146 391074
rect 542382 390838 542414 391074
rect 19794 390806 542414 390838
rect -2966 390454 586890 390486
rect -2966 390218 -2934 390454
rect -2698 390218 -2614 390454
rect -2378 390218 10826 390454
rect 11062 390218 11146 390454
rect 11382 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 46826 390454
rect 47062 390218 47146 390454
rect 47382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 82826 390454
rect 83062 390218 83146 390454
rect 83382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 118826 390454
rect 119062 390218 119146 390454
rect 119382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 154826 390454
rect 155062 390218 155146 390454
rect 155382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 190826 390454
rect 191062 390218 191146 390454
rect 191382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 226826 390454
rect 227062 390218 227146 390454
rect 227382 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 262826 390454
rect 263062 390218 263146 390454
rect 263382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 298826 390454
rect 299062 390218 299146 390454
rect 299382 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 334826 390454
rect 335062 390218 335146 390454
rect 335382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 370826 390454
rect 371062 390218 371146 390454
rect 371382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 406826 390454
rect 407062 390218 407146 390454
rect 407382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 442826 390454
rect 443062 390218 443146 390454
rect 443382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 478826 390454
rect 479062 390218 479146 390454
rect 479382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 514826 390454
rect 515062 390218 515146 390454
rect 515382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 550826 390454
rect 551062 390218 551146 390454
rect 551382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 586302 390454
rect 586538 390218 586622 390454
rect 586858 390218 586890 390454
rect -2966 390134 586890 390218
rect -2966 389898 -2934 390134
rect -2698 389898 -2614 390134
rect -2378 389898 10826 390134
rect 11062 389898 11146 390134
rect 11382 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 46826 390134
rect 47062 389898 47146 390134
rect 47382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 82826 390134
rect 83062 389898 83146 390134
rect 83382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 118826 390134
rect 119062 389898 119146 390134
rect 119382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 154826 390134
rect 155062 389898 155146 390134
rect 155382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 190826 390134
rect 191062 389898 191146 390134
rect 191382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 226826 390134
rect 227062 389898 227146 390134
rect 227382 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 262826 390134
rect 263062 389898 263146 390134
rect 263382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 298826 390134
rect 299062 389898 299146 390134
rect 299382 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 334826 390134
rect 335062 389898 335146 390134
rect 335382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 370826 390134
rect 371062 389898 371146 390134
rect 371382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 406826 390134
rect 407062 389898 407146 390134
rect 407382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 442826 390134
rect 443062 389898 443146 390134
rect 443382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 478826 390134
rect 479062 389898 479146 390134
rect 479382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 514826 390134
rect 515062 389898 515146 390134
rect 515382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 550826 390134
rect 551062 389898 551146 390134
rect 551382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 586302 390134
rect 586538 389898 586622 390134
rect 586858 389898 586890 390134
rect -2966 389866 586890 389898
rect -2966 381454 586890 381486
rect -2966 381218 -1974 381454
rect -1738 381218 -1654 381454
rect -1418 381218 1826 381454
rect 2062 381218 2146 381454
rect 2382 381218 19952 381454
rect 20188 381218 25882 381454
rect 26118 381218 31813 381454
rect 32049 381218 46952 381454
rect 47188 381218 52882 381454
rect 53118 381218 58813 381454
rect 59049 381218 73952 381454
rect 74188 381218 79882 381454
rect 80118 381218 85813 381454
rect 86049 381218 100952 381454
rect 101188 381218 106882 381454
rect 107118 381218 112813 381454
rect 113049 381218 127952 381454
rect 128188 381218 133882 381454
rect 134118 381218 139813 381454
rect 140049 381218 154952 381454
rect 155188 381218 160882 381454
rect 161118 381218 166813 381454
rect 167049 381218 181952 381454
rect 182188 381218 187882 381454
rect 188118 381218 193813 381454
rect 194049 381218 208952 381454
rect 209188 381218 214882 381454
rect 215118 381218 220813 381454
rect 221049 381218 235952 381454
rect 236188 381218 241882 381454
rect 242118 381218 247813 381454
rect 248049 381218 262952 381454
rect 263188 381218 268882 381454
rect 269118 381218 274813 381454
rect 275049 381218 289952 381454
rect 290188 381218 295882 381454
rect 296118 381218 301813 381454
rect 302049 381218 316952 381454
rect 317188 381218 322882 381454
rect 323118 381218 328813 381454
rect 329049 381218 343952 381454
rect 344188 381218 349882 381454
rect 350118 381218 355813 381454
rect 356049 381218 370952 381454
rect 371188 381218 376882 381454
rect 377118 381218 382813 381454
rect 383049 381218 397952 381454
rect 398188 381218 403882 381454
rect 404118 381218 409813 381454
rect 410049 381218 424952 381454
rect 425188 381218 430882 381454
rect 431118 381218 436813 381454
rect 437049 381218 451952 381454
rect 452188 381218 457882 381454
rect 458118 381218 463813 381454
rect 464049 381218 478952 381454
rect 479188 381218 484882 381454
rect 485118 381218 490813 381454
rect 491049 381218 505952 381454
rect 506188 381218 511882 381454
rect 512118 381218 517813 381454
rect 518049 381218 532952 381454
rect 533188 381218 538882 381454
rect 539118 381218 544813 381454
rect 545049 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 577826 381454
rect 578062 381218 578146 381454
rect 578382 381218 585342 381454
rect 585578 381218 585662 381454
rect 585898 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -1974 381134
rect -1738 380898 -1654 381134
rect -1418 380898 1826 381134
rect 2062 380898 2146 381134
rect 2382 380898 19952 381134
rect 20188 380898 25882 381134
rect 26118 380898 31813 381134
rect 32049 380898 46952 381134
rect 47188 380898 52882 381134
rect 53118 380898 58813 381134
rect 59049 380898 73952 381134
rect 74188 380898 79882 381134
rect 80118 380898 85813 381134
rect 86049 380898 100952 381134
rect 101188 380898 106882 381134
rect 107118 380898 112813 381134
rect 113049 380898 127952 381134
rect 128188 380898 133882 381134
rect 134118 380898 139813 381134
rect 140049 380898 154952 381134
rect 155188 380898 160882 381134
rect 161118 380898 166813 381134
rect 167049 380898 181952 381134
rect 182188 380898 187882 381134
rect 188118 380898 193813 381134
rect 194049 380898 208952 381134
rect 209188 380898 214882 381134
rect 215118 380898 220813 381134
rect 221049 380898 235952 381134
rect 236188 380898 241882 381134
rect 242118 380898 247813 381134
rect 248049 380898 262952 381134
rect 263188 380898 268882 381134
rect 269118 380898 274813 381134
rect 275049 380898 289952 381134
rect 290188 380898 295882 381134
rect 296118 380898 301813 381134
rect 302049 380898 316952 381134
rect 317188 380898 322882 381134
rect 323118 380898 328813 381134
rect 329049 380898 343952 381134
rect 344188 380898 349882 381134
rect 350118 380898 355813 381134
rect 356049 380898 370952 381134
rect 371188 380898 376882 381134
rect 377118 380898 382813 381134
rect 383049 380898 397952 381134
rect 398188 380898 403882 381134
rect 404118 380898 409813 381134
rect 410049 380898 424952 381134
rect 425188 380898 430882 381134
rect 431118 380898 436813 381134
rect 437049 380898 451952 381134
rect 452188 380898 457882 381134
rect 458118 380898 463813 381134
rect 464049 380898 478952 381134
rect 479188 380898 484882 381134
rect 485118 380898 490813 381134
rect 491049 380898 505952 381134
rect 506188 380898 511882 381134
rect 512118 380898 517813 381134
rect 518049 380898 532952 381134
rect 533188 380898 538882 381134
rect 539118 380898 544813 381134
rect 545049 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 577826 381134
rect 578062 380898 578146 381134
rect 578382 380898 585342 381134
rect 585578 380898 585662 381134
rect 585898 380898 586890 381134
rect -2966 380866 586890 380898
rect -2966 372454 586890 372486
rect -2966 372218 -2934 372454
rect -2698 372218 -2614 372454
rect -2378 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 22916 372454
rect 23152 372218 28847 372454
rect 29083 372218 49916 372454
rect 50152 372218 55847 372454
rect 56083 372218 76916 372454
rect 77152 372218 82847 372454
rect 83083 372218 103916 372454
rect 104152 372218 109847 372454
rect 110083 372218 130916 372454
rect 131152 372218 136847 372454
rect 137083 372218 157916 372454
rect 158152 372218 163847 372454
rect 164083 372218 184916 372454
rect 185152 372218 190847 372454
rect 191083 372218 211916 372454
rect 212152 372218 217847 372454
rect 218083 372218 238916 372454
rect 239152 372218 244847 372454
rect 245083 372218 265916 372454
rect 266152 372218 271847 372454
rect 272083 372218 292916 372454
rect 293152 372218 298847 372454
rect 299083 372218 319916 372454
rect 320152 372218 325847 372454
rect 326083 372218 346916 372454
rect 347152 372218 352847 372454
rect 353083 372218 373916 372454
rect 374152 372218 379847 372454
rect 380083 372218 400916 372454
rect 401152 372218 406847 372454
rect 407083 372218 427916 372454
rect 428152 372218 433847 372454
rect 434083 372218 454916 372454
rect 455152 372218 460847 372454
rect 461083 372218 481916 372454
rect 482152 372218 487847 372454
rect 488083 372218 508916 372454
rect 509152 372218 514847 372454
rect 515083 372218 535916 372454
rect 536152 372218 541847 372454
rect 542083 372218 568826 372454
rect 569062 372218 569146 372454
rect 569382 372218 586302 372454
rect 586538 372218 586622 372454
rect 586858 372218 586890 372454
rect -2966 372134 586890 372218
rect -2966 371898 -2934 372134
rect -2698 371898 -2614 372134
rect -2378 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 22916 372134
rect 23152 371898 28847 372134
rect 29083 371898 49916 372134
rect 50152 371898 55847 372134
rect 56083 371898 76916 372134
rect 77152 371898 82847 372134
rect 83083 371898 103916 372134
rect 104152 371898 109847 372134
rect 110083 371898 130916 372134
rect 131152 371898 136847 372134
rect 137083 371898 157916 372134
rect 158152 371898 163847 372134
rect 164083 371898 184916 372134
rect 185152 371898 190847 372134
rect 191083 371898 211916 372134
rect 212152 371898 217847 372134
rect 218083 371898 238916 372134
rect 239152 371898 244847 372134
rect 245083 371898 265916 372134
rect 266152 371898 271847 372134
rect 272083 371898 292916 372134
rect 293152 371898 298847 372134
rect 299083 371898 319916 372134
rect 320152 371898 325847 372134
rect 326083 371898 346916 372134
rect 347152 371898 352847 372134
rect 353083 371898 373916 372134
rect 374152 371898 379847 372134
rect 380083 371898 400916 372134
rect 401152 371898 406847 372134
rect 407083 371898 427916 372134
rect 428152 371898 433847 372134
rect 434083 371898 454916 372134
rect 455152 371898 460847 372134
rect 461083 371898 481916 372134
rect 482152 371898 487847 372134
rect 488083 371898 508916 372134
rect 509152 371898 514847 372134
rect 515083 371898 535916 372134
rect 536152 371898 541847 372134
rect 542083 371898 568826 372134
rect 569062 371898 569146 372134
rect 569382 371898 586302 372134
rect 586538 371898 586622 372134
rect 586858 371898 586890 372134
rect -2966 371866 586890 371898
rect 28794 364394 551414 364426
rect 28794 364158 28826 364394
rect 29062 364158 29146 364394
rect 29382 364158 46826 364394
rect 47062 364158 47146 364394
rect 47382 364158 64826 364394
rect 65062 364158 65146 364394
rect 65382 364158 82826 364394
rect 83062 364158 83146 364394
rect 83382 364158 100826 364394
rect 101062 364158 101146 364394
rect 101382 364158 118826 364394
rect 119062 364158 119146 364394
rect 119382 364158 136826 364394
rect 137062 364158 137146 364394
rect 137382 364158 154826 364394
rect 155062 364158 155146 364394
rect 155382 364158 172826 364394
rect 173062 364158 173146 364394
rect 173382 364158 190826 364394
rect 191062 364158 191146 364394
rect 191382 364158 208826 364394
rect 209062 364158 209146 364394
rect 209382 364158 226826 364394
rect 227062 364158 227146 364394
rect 227382 364158 244826 364394
rect 245062 364158 245146 364394
rect 245382 364158 262826 364394
rect 263062 364158 263146 364394
rect 263382 364158 280826 364394
rect 281062 364158 281146 364394
rect 281382 364158 298826 364394
rect 299062 364158 299146 364394
rect 299382 364158 316826 364394
rect 317062 364158 317146 364394
rect 317382 364158 334826 364394
rect 335062 364158 335146 364394
rect 335382 364158 352826 364394
rect 353062 364158 353146 364394
rect 353382 364158 370826 364394
rect 371062 364158 371146 364394
rect 371382 364158 388826 364394
rect 389062 364158 389146 364394
rect 389382 364158 406826 364394
rect 407062 364158 407146 364394
rect 407382 364158 424826 364394
rect 425062 364158 425146 364394
rect 425382 364158 442826 364394
rect 443062 364158 443146 364394
rect 443382 364158 460826 364394
rect 461062 364158 461146 364394
rect 461382 364158 478826 364394
rect 479062 364158 479146 364394
rect 479382 364158 496826 364394
rect 497062 364158 497146 364394
rect 497382 364158 514826 364394
rect 515062 364158 515146 364394
rect 515382 364158 532826 364394
rect 533062 364158 533146 364394
rect 533382 364158 550826 364394
rect 551062 364158 551146 364394
rect 551382 364158 551414 364394
rect 28794 364074 551414 364158
rect 28794 363838 28826 364074
rect 29062 363838 29146 364074
rect 29382 363838 46826 364074
rect 47062 363838 47146 364074
rect 47382 363838 64826 364074
rect 65062 363838 65146 364074
rect 65382 363838 82826 364074
rect 83062 363838 83146 364074
rect 83382 363838 100826 364074
rect 101062 363838 101146 364074
rect 101382 363838 118826 364074
rect 119062 363838 119146 364074
rect 119382 363838 136826 364074
rect 137062 363838 137146 364074
rect 137382 363838 154826 364074
rect 155062 363838 155146 364074
rect 155382 363838 172826 364074
rect 173062 363838 173146 364074
rect 173382 363838 190826 364074
rect 191062 363838 191146 364074
rect 191382 363838 208826 364074
rect 209062 363838 209146 364074
rect 209382 363838 226826 364074
rect 227062 363838 227146 364074
rect 227382 363838 244826 364074
rect 245062 363838 245146 364074
rect 245382 363838 262826 364074
rect 263062 363838 263146 364074
rect 263382 363838 280826 364074
rect 281062 363838 281146 364074
rect 281382 363838 298826 364074
rect 299062 363838 299146 364074
rect 299382 363838 316826 364074
rect 317062 363838 317146 364074
rect 317382 363838 334826 364074
rect 335062 363838 335146 364074
rect 335382 363838 352826 364074
rect 353062 363838 353146 364074
rect 353382 363838 370826 364074
rect 371062 363838 371146 364074
rect 371382 363838 388826 364074
rect 389062 363838 389146 364074
rect 389382 363838 406826 364074
rect 407062 363838 407146 364074
rect 407382 363838 424826 364074
rect 425062 363838 425146 364074
rect 425382 363838 442826 364074
rect 443062 363838 443146 364074
rect 443382 363838 460826 364074
rect 461062 363838 461146 364074
rect 461382 363838 478826 364074
rect 479062 363838 479146 364074
rect 479382 363838 496826 364074
rect 497062 363838 497146 364074
rect 497382 363838 514826 364074
rect 515062 363838 515146 364074
rect 515382 363838 532826 364074
rect 533062 363838 533146 364074
rect 533382 363838 550826 364074
rect 551062 363838 551146 364074
rect 551382 363838 551414 364074
rect 28794 363806 551414 363838
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 19826 363454
rect 20062 363218 20146 363454
rect 20382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 55826 363454
rect 56062 363218 56146 363454
rect 56382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 91826 363454
rect 92062 363218 92146 363454
rect 92382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 127826 363454
rect 128062 363218 128146 363454
rect 128382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 163826 363454
rect 164062 363218 164146 363454
rect 164382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 199826 363454
rect 200062 363218 200146 363454
rect 200382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 235826 363454
rect 236062 363218 236146 363454
rect 236382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 271826 363454
rect 272062 363218 272146 363454
rect 272382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 307826 363454
rect 308062 363218 308146 363454
rect 308382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 343826 363454
rect 344062 363218 344146 363454
rect 344382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 379826 363454
rect 380062 363218 380146 363454
rect 380382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 415826 363454
rect 416062 363218 416146 363454
rect 416382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 451826 363454
rect 452062 363218 452146 363454
rect 452382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 487826 363454
rect 488062 363218 488146 363454
rect 488382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 523826 363454
rect 524062 363218 524146 363454
rect 524382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 559826 363454
rect 560062 363218 560146 363454
rect 560382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 19826 363134
rect 20062 362898 20146 363134
rect 20382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 55826 363134
rect 56062 362898 56146 363134
rect 56382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 91826 363134
rect 92062 362898 92146 363134
rect 92382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 127826 363134
rect 128062 362898 128146 363134
rect 128382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 163826 363134
rect 164062 362898 164146 363134
rect 164382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 199826 363134
rect 200062 362898 200146 363134
rect 200382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 235826 363134
rect 236062 362898 236146 363134
rect 236382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 271826 363134
rect 272062 362898 272146 363134
rect 272382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 307826 363134
rect 308062 362898 308146 363134
rect 308382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 343826 363134
rect 344062 362898 344146 363134
rect 344382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 379826 363134
rect 380062 362898 380146 363134
rect 380382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 415826 363134
rect 416062 362898 416146 363134
rect 416382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 451826 363134
rect 452062 362898 452146 363134
rect 452382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 487826 363134
rect 488062 362898 488146 363134
rect 488382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 523826 363134
rect 524062 362898 524146 363134
rect 524382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 559826 363134
rect 560062 362898 560146 363134
rect 560382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -2966 354454 586890 354486
rect -2966 354218 -2934 354454
rect -2698 354218 -2614 354454
rect -2378 354218 10826 354454
rect 11062 354218 11146 354454
rect 11382 354218 22916 354454
rect 23152 354218 28847 354454
rect 29083 354218 49916 354454
rect 50152 354218 55847 354454
rect 56083 354218 76916 354454
rect 77152 354218 82847 354454
rect 83083 354218 103916 354454
rect 104152 354218 109847 354454
rect 110083 354218 130916 354454
rect 131152 354218 136847 354454
rect 137083 354218 157916 354454
rect 158152 354218 163847 354454
rect 164083 354218 184916 354454
rect 185152 354218 190847 354454
rect 191083 354218 211916 354454
rect 212152 354218 217847 354454
rect 218083 354218 238916 354454
rect 239152 354218 244847 354454
rect 245083 354218 265916 354454
rect 266152 354218 271847 354454
rect 272083 354218 292916 354454
rect 293152 354218 298847 354454
rect 299083 354218 319916 354454
rect 320152 354218 325847 354454
rect 326083 354218 346916 354454
rect 347152 354218 352847 354454
rect 353083 354218 373916 354454
rect 374152 354218 379847 354454
rect 380083 354218 400916 354454
rect 401152 354218 406847 354454
rect 407083 354218 427916 354454
rect 428152 354218 433847 354454
rect 434083 354218 454916 354454
rect 455152 354218 460847 354454
rect 461083 354218 481916 354454
rect 482152 354218 487847 354454
rect 488083 354218 508916 354454
rect 509152 354218 514847 354454
rect 515083 354218 535916 354454
rect 536152 354218 541847 354454
rect 542083 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 586302 354454
rect 586538 354218 586622 354454
rect 586858 354218 586890 354454
rect -2966 354134 586890 354218
rect -2966 353898 -2934 354134
rect -2698 353898 -2614 354134
rect -2378 353898 10826 354134
rect 11062 353898 11146 354134
rect 11382 353898 22916 354134
rect 23152 353898 28847 354134
rect 29083 353898 49916 354134
rect 50152 353898 55847 354134
rect 56083 353898 76916 354134
rect 77152 353898 82847 354134
rect 83083 353898 103916 354134
rect 104152 353898 109847 354134
rect 110083 353898 130916 354134
rect 131152 353898 136847 354134
rect 137083 353898 157916 354134
rect 158152 353898 163847 354134
rect 164083 353898 184916 354134
rect 185152 353898 190847 354134
rect 191083 353898 211916 354134
rect 212152 353898 217847 354134
rect 218083 353898 238916 354134
rect 239152 353898 244847 354134
rect 245083 353898 265916 354134
rect 266152 353898 271847 354134
rect 272083 353898 292916 354134
rect 293152 353898 298847 354134
rect 299083 353898 319916 354134
rect 320152 353898 325847 354134
rect 326083 353898 346916 354134
rect 347152 353898 352847 354134
rect 353083 353898 373916 354134
rect 374152 353898 379847 354134
rect 380083 353898 400916 354134
rect 401152 353898 406847 354134
rect 407083 353898 427916 354134
rect 428152 353898 433847 354134
rect 434083 353898 454916 354134
rect 455152 353898 460847 354134
rect 461083 353898 481916 354134
rect 482152 353898 487847 354134
rect 488083 353898 508916 354134
rect 509152 353898 514847 354134
rect 515083 353898 535916 354134
rect 536152 353898 541847 354134
rect 542083 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 586302 354134
rect 586538 353898 586622 354134
rect 586858 353898 586890 354134
rect -2966 353866 586890 353898
rect -2966 345454 586890 345486
rect -2966 345218 -1974 345454
rect -1738 345218 -1654 345454
rect -1418 345218 1826 345454
rect 2062 345218 2146 345454
rect 2382 345218 19952 345454
rect 20188 345218 25882 345454
rect 26118 345218 31813 345454
rect 32049 345218 46952 345454
rect 47188 345218 52882 345454
rect 53118 345218 58813 345454
rect 59049 345218 73952 345454
rect 74188 345218 79882 345454
rect 80118 345218 85813 345454
rect 86049 345218 100952 345454
rect 101188 345218 106882 345454
rect 107118 345218 112813 345454
rect 113049 345218 127952 345454
rect 128188 345218 133882 345454
rect 134118 345218 139813 345454
rect 140049 345218 154952 345454
rect 155188 345218 160882 345454
rect 161118 345218 166813 345454
rect 167049 345218 181952 345454
rect 182188 345218 187882 345454
rect 188118 345218 193813 345454
rect 194049 345218 208952 345454
rect 209188 345218 214882 345454
rect 215118 345218 220813 345454
rect 221049 345218 235952 345454
rect 236188 345218 241882 345454
rect 242118 345218 247813 345454
rect 248049 345218 262952 345454
rect 263188 345218 268882 345454
rect 269118 345218 274813 345454
rect 275049 345218 289952 345454
rect 290188 345218 295882 345454
rect 296118 345218 301813 345454
rect 302049 345218 316952 345454
rect 317188 345218 322882 345454
rect 323118 345218 328813 345454
rect 329049 345218 343952 345454
rect 344188 345218 349882 345454
rect 350118 345218 355813 345454
rect 356049 345218 370952 345454
rect 371188 345218 376882 345454
rect 377118 345218 382813 345454
rect 383049 345218 397952 345454
rect 398188 345218 403882 345454
rect 404118 345218 409813 345454
rect 410049 345218 424952 345454
rect 425188 345218 430882 345454
rect 431118 345218 436813 345454
rect 437049 345218 451952 345454
rect 452188 345218 457882 345454
rect 458118 345218 463813 345454
rect 464049 345218 478952 345454
rect 479188 345218 484882 345454
rect 485118 345218 490813 345454
rect 491049 345218 505952 345454
rect 506188 345218 511882 345454
rect 512118 345218 517813 345454
rect 518049 345218 532952 345454
rect 533188 345218 538882 345454
rect 539118 345218 544813 345454
rect 545049 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 577826 345454
rect 578062 345218 578146 345454
rect 578382 345218 585342 345454
rect 585578 345218 585662 345454
rect 585898 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -1974 345134
rect -1738 344898 -1654 345134
rect -1418 344898 1826 345134
rect 2062 344898 2146 345134
rect 2382 344898 19952 345134
rect 20188 344898 25882 345134
rect 26118 344898 31813 345134
rect 32049 344898 46952 345134
rect 47188 344898 52882 345134
rect 53118 344898 58813 345134
rect 59049 344898 73952 345134
rect 74188 344898 79882 345134
rect 80118 344898 85813 345134
rect 86049 344898 100952 345134
rect 101188 344898 106882 345134
rect 107118 344898 112813 345134
rect 113049 344898 127952 345134
rect 128188 344898 133882 345134
rect 134118 344898 139813 345134
rect 140049 344898 154952 345134
rect 155188 344898 160882 345134
rect 161118 344898 166813 345134
rect 167049 344898 181952 345134
rect 182188 344898 187882 345134
rect 188118 344898 193813 345134
rect 194049 344898 208952 345134
rect 209188 344898 214882 345134
rect 215118 344898 220813 345134
rect 221049 344898 235952 345134
rect 236188 344898 241882 345134
rect 242118 344898 247813 345134
rect 248049 344898 262952 345134
rect 263188 344898 268882 345134
rect 269118 344898 274813 345134
rect 275049 344898 289952 345134
rect 290188 344898 295882 345134
rect 296118 344898 301813 345134
rect 302049 344898 316952 345134
rect 317188 344898 322882 345134
rect 323118 344898 328813 345134
rect 329049 344898 343952 345134
rect 344188 344898 349882 345134
rect 350118 344898 355813 345134
rect 356049 344898 370952 345134
rect 371188 344898 376882 345134
rect 377118 344898 382813 345134
rect 383049 344898 397952 345134
rect 398188 344898 403882 345134
rect 404118 344898 409813 345134
rect 410049 344898 424952 345134
rect 425188 344898 430882 345134
rect 431118 344898 436813 345134
rect 437049 344898 451952 345134
rect 452188 344898 457882 345134
rect 458118 344898 463813 345134
rect 464049 344898 478952 345134
rect 479188 344898 484882 345134
rect 485118 344898 490813 345134
rect 491049 344898 505952 345134
rect 506188 344898 511882 345134
rect 512118 344898 517813 345134
rect 518049 344898 532952 345134
rect 533188 344898 538882 345134
rect 539118 344898 544813 345134
rect 545049 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 577826 345134
rect 578062 344898 578146 345134
rect 578382 344898 585342 345134
rect 585578 344898 585662 345134
rect 585898 344898 586890 345134
rect -2966 344866 586890 344898
rect 19794 337394 542414 337426
rect 19794 337158 19826 337394
rect 20062 337158 20146 337394
rect 20382 337158 37826 337394
rect 38062 337158 38146 337394
rect 38382 337158 55826 337394
rect 56062 337158 56146 337394
rect 56382 337158 73826 337394
rect 74062 337158 74146 337394
rect 74382 337158 91826 337394
rect 92062 337158 92146 337394
rect 92382 337158 109826 337394
rect 110062 337158 110146 337394
rect 110382 337158 127826 337394
rect 128062 337158 128146 337394
rect 128382 337158 145826 337394
rect 146062 337158 146146 337394
rect 146382 337158 163826 337394
rect 164062 337158 164146 337394
rect 164382 337158 181826 337394
rect 182062 337158 182146 337394
rect 182382 337158 199826 337394
rect 200062 337158 200146 337394
rect 200382 337158 217826 337394
rect 218062 337158 218146 337394
rect 218382 337158 235826 337394
rect 236062 337158 236146 337394
rect 236382 337158 253826 337394
rect 254062 337158 254146 337394
rect 254382 337158 271826 337394
rect 272062 337158 272146 337394
rect 272382 337158 289826 337394
rect 290062 337158 290146 337394
rect 290382 337158 307826 337394
rect 308062 337158 308146 337394
rect 308382 337158 325826 337394
rect 326062 337158 326146 337394
rect 326382 337158 343826 337394
rect 344062 337158 344146 337394
rect 344382 337158 361826 337394
rect 362062 337158 362146 337394
rect 362382 337158 379826 337394
rect 380062 337158 380146 337394
rect 380382 337158 397826 337394
rect 398062 337158 398146 337394
rect 398382 337158 415826 337394
rect 416062 337158 416146 337394
rect 416382 337158 433826 337394
rect 434062 337158 434146 337394
rect 434382 337158 451826 337394
rect 452062 337158 452146 337394
rect 452382 337158 469826 337394
rect 470062 337158 470146 337394
rect 470382 337158 487826 337394
rect 488062 337158 488146 337394
rect 488382 337158 505826 337394
rect 506062 337158 506146 337394
rect 506382 337158 523826 337394
rect 524062 337158 524146 337394
rect 524382 337158 541826 337394
rect 542062 337158 542146 337394
rect 542382 337158 542414 337394
rect 19794 337074 542414 337158
rect 19794 336838 19826 337074
rect 20062 336838 20146 337074
rect 20382 336838 37826 337074
rect 38062 336838 38146 337074
rect 38382 336838 55826 337074
rect 56062 336838 56146 337074
rect 56382 336838 73826 337074
rect 74062 336838 74146 337074
rect 74382 336838 91826 337074
rect 92062 336838 92146 337074
rect 92382 336838 109826 337074
rect 110062 336838 110146 337074
rect 110382 336838 127826 337074
rect 128062 336838 128146 337074
rect 128382 336838 145826 337074
rect 146062 336838 146146 337074
rect 146382 336838 163826 337074
rect 164062 336838 164146 337074
rect 164382 336838 181826 337074
rect 182062 336838 182146 337074
rect 182382 336838 199826 337074
rect 200062 336838 200146 337074
rect 200382 336838 217826 337074
rect 218062 336838 218146 337074
rect 218382 336838 235826 337074
rect 236062 336838 236146 337074
rect 236382 336838 253826 337074
rect 254062 336838 254146 337074
rect 254382 336838 271826 337074
rect 272062 336838 272146 337074
rect 272382 336838 289826 337074
rect 290062 336838 290146 337074
rect 290382 336838 307826 337074
rect 308062 336838 308146 337074
rect 308382 336838 325826 337074
rect 326062 336838 326146 337074
rect 326382 336838 343826 337074
rect 344062 336838 344146 337074
rect 344382 336838 361826 337074
rect 362062 336838 362146 337074
rect 362382 336838 379826 337074
rect 380062 336838 380146 337074
rect 380382 336838 397826 337074
rect 398062 336838 398146 337074
rect 398382 336838 415826 337074
rect 416062 336838 416146 337074
rect 416382 336838 433826 337074
rect 434062 336838 434146 337074
rect 434382 336838 451826 337074
rect 452062 336838 452146 337074
rect 452382 336838 469826 337074
rect 470062 336838 470146 337074
rect 470382 336838 487826 337074
rect 488062 336838 488146 337074
rect 488382 336838 505826 337074
rect 506062 336838 506146 337074
rect 506382 336838 523826 337074
rect 524062 336838 524146 337074
rect 524382 336838 541826 337074
rect 542062 336838 542146 337074
rect 542382 336838 542414 337074
rect 19794 336806 542414 336838
rect -2966 336454 586890 336486
rect -2966 336218 -2934 336454
rect -2698 336218 -2614 336454
rect -2378 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 28826 336454
rect 29062 336218 29146 336454
rect 29382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 64826 336454
rect 65062 336218 65146 336454
rect 65382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 100826 336454
rect 101062 336218 101146 336454
rect 101382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 136826 336454
rect 137062 336218 137146 336454
rect 137382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 172826 336454
rect 173062 336218 173146 336454
rect 173382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 208826 336454
rect 209062 336218 209146 336454
rect 209382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 244826 336454
rect 245062 336218 245146 336454
rect 245382 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 280826 336454
rect 281062 336218 281146 336454
rect 281382 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 316826 336454
rect 317062 336218 317146 336454
rect 317382 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 352826 336454
rect 353062 336218 353146 336454
rect 353382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 388826 336454
rect 389062 336218 389146 336454
rect 389382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 424826 336454
rect 425062 336218 425146 336454
rect 425382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 460826 336454
rect 461062 336218 461146 336454
rect 461382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 496826 336454
rect 497062 336218 497146 336454
rect 497382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 532826 336454
rect 533062 336218 533146 336454
rect 533382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 568826 336454
rect 569062 336218 569146 336454
rect 569382 336218 586302 336454
rect 586538 336218 586622 336454
rect 586858 336218 586890 336454
rect -2966 336134 586890 336218
rect -2966 335898 -2934 336134
rect -2698 335898 -2614 336134
rect -2378 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 28826 336134
rect 29062 335898 29146 336134
rect 29382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 64826 336134
rect 65062 335898 65146 336134
rect 65382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 100826 336134
rect 101062 335898 101146 336134
rect 101382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 136826 336134
rect 137062 335898 137146 336134
rect 137382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 172826 336134
rect 173062 335898 173146 336134
rect 173382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 208826 336134
rect 209062 335898 209146 336134
rect 209382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 244826 336134
rect 245062 335898 245146 336134
rect 245382 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 280826 336134
rect 281062 335898 281146 336134
rect 281382 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 316826 336134
rect 317062 335898 317146 336134
rect 317382 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 352826 336134
rect 353062 335898 353146 336134
rect 353382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 388826 336134
rect 389062 335898 389146 336134
rect 389382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 424826 336134
rect 425062 335898 425146 336134
rect 425382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 460826 336134
rect 461062 335898 461146 336134
rect 461382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 496826 336134
rect 497062 335898 497146 336134
rect 497382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 532826 336134
rect 533062 335898 533146 336134
rect 533382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 568826 336134
rect 569062 335898 569146 336134
rect 569382 335898 586302 336134
rect 586538 335898 586622 336134
rect 586858 335898 586890 336134
rect -2966 335866 586890 335898
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 19952 327454
rect 20188 327218 25882 327454
rect 26118 327218 31813 327454
rect 32049 327218 46952 327454
rect 47188 327218 52882 327454
rect 53118 327218 58813 327454
rect 59049 327218 73952 327454
rect 74188 327218 79882 327454
rect 80118 327218 85813 327454
rect 86049 327218 100952 327454
rect 101188 327218 106882 327454
rect 107118 327218 112813 327454
rect 113049 327218 127952 327454
rect 128188 327218 133882 327454
rect 134118 327218 139813 327454
rect 140049 327218 154952 327454
rect 155188 327218 160882 327454
rect 161118 327218 166813 327454
rect 167049 327218 181952 327454
rect 182188 327218 187882 327454
rect 188118 327218 193813 327454
rect 194049 327218 208952 327454
rect 209188 327218 214882 327454
rect 215118 327218 220813 327454
rect 221049 327218 235952 327454
rect 236188 327218 241882 327454
rect 242118 327218 247813 327454
rect 248049 327218 262952 327454
rect 263188 327218 268882 327454
rect 269118 327218 274813 327454
rect 275049 327218 289952 327454
rect 290188 327218 295882 327454
rect 296118 327218 301813 327454
rect 302049 327218 316952 327454
rect 317188 327218 322882 327454
rect 323118 327218 328813 327454
rect 329049 327218 343952 327454
rect 344188 327218 349882 327454
rect 350118 327218 355813 327454
rect 356049 327218 370952 327454
rect 371188 327218 376882 327454
rect 377118 327218 382813 327454
rect 383049 327218 397952 327454
rect 398188 327218 403882 327454
rect 404118 327218 409813 327454
rect 410049 327218 424952 327454
rect 425188 327218 430882 327454
rect 431118 327218 436813 327454
rect 437049 327218 451952 327454
rect 452188 327218 457882 327454
rect 458118 327218 463813 327454
rect 464049 327218 478952 327454
rect 479188 327218 484882 327454
rect 485118 327218 490813 327454
rect 491049 327218 505952 327454
rect 506188 327218 511882 327454
rect 512118 327218 517813 327454
rect 518049 327218 532952 327454
rect 533188 327218 538882 327454
rect 539118 327218 544813 327454
rect 545049 327218 559826 327454
rect 560062 327218 560146 327454
rect 560382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 19952 327134
rect 20188 326898 25882 327134
rect 26118 326898 31813 327134
rect 32049 326898 46952 327134
rect 47188 326898 52882 327134
rect 53118 326898 58813 327134
rect 59049 326898 73952 327134
rect 74188 326898 79882 327134
rect 80118 326898 85813 327134
rect 86049 326898 100952 327134
rect 101188 326898 106882 327134
rect 107118 326898 112813 327134
rect 113049 326898 127952 327134
rect 128188 326898 133882 327134
rect 134118 326898 139813 327134
rect 140049 326898 154952 327134
rect 155188 326898 160882 327134
rect 161118 326898 166813 327134
rect 167049 326898 181952 327134
rect 182188 326898 187882 327134
rect 188118 326898 193813 327134
rect 194049 326898 208952 327134
rect 209188 326898 214882 327134
rect 215118 326898 220813 327134
rect 221049 326898 235952 327134
rect 236188 326898 241882 327134
rect 242118 326898 247813 327134
rect 248049 326898 262952 327134
rect 263188 326898 268882 327134
rect 269118 326898 274813 327134
rect 275049 326898 289952 327134
rect 290188 326898 295882 327134
rect 296118 326898 301813 327134
rect 302049 326898 316952 327134
rect 317188 326898 322882 327134
rect 323118 326898 328813 327134
rect 329049 326898 343952 327134
rect 344188 326898 349882 327134
rect 350118 326898 355813 327134
rect 356049 326898 370952 327134
rect 371188 326898 376882 327134
rect 377118 326898 382813 327134
rect 383049 326898 397952 327134
rect 398188 326898 403882 327134
rect 404118 326898 409813 327134
rect 410049 326898 424952 327134
rect 425188 326898 430882 327134
rect 431118 326898 436813 327134
rect 437049 326898 451952 327134
rect 452188 326898 457882 327134
rect 458118 326898 463813 327134
rect 464049 326898 478952 327134
rect 479188 326898 484882 327134
rect 485118 326898 490813 327134
rect 491049 326898 505952 327134
rect 506188 326898 511882 327134
rect 512118 326898 517813 327134
rect 518049 326898 532952 327134
rect 533188 326898 538882 327134
rect 539118 326898 544813 327134
rect 545049 326898 559826 327134
rect 560062 326898 560146 327134
rect 560382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -2966 318454 586890 318486
rect -2966 318218 -2934 318454
rect -2698 318218 -2614 318454
rect -2378 318218 10826 318454
rect 11062 318218 11146 318454
rect 11382 318218 22916 318454
rect 23152 318218 28847 318454
rect 29083 318218 49916 318454
rect 50152 318218 55847 318454
rect 56083 318218 76916 318454
rect 77152 318218 82847 318454
rect 83083 318218 103916 318454
rect 104152 318218 109847 318454
rect 110083 318218 130916 318454
rect 131152 318218 136847 318454
rect 137083 318218 157916 318454
rect 158152 318218 163847 318454
rect 164083 318218 184916 318454
rect 185152 318218 190847 318454
rect 191083 318218 211916 318454
rect 212152 318218 217847 318454
rect 218083 318218 238916 318454
rect 239152 318218 244847 318454
rect 245083 318218 265916 318454
rect 266152 318218 271847 318454
rect 272083 318218 292916 318454
rect 293152 318218 298847 318454
rect 299083 318218 319916 318454
rect 320152 318218 325847 318454
rect 326083 318218 346916 318454
rect 347152 318218 352847 318454
rect 353083 318218 373916 318454
rect 374152 318218 379847 318454
rect 380083 318218 400916 318454
rect 401152 318218 406847 318454
rect 407083 318218 427916 318454
rect 428152 318218 433847 318454
rect 434083 318218 454916 318454
rect 455152 318218 460847 318454
rect 461083 318218 481916 318454
rect 482152 318218 487847 318454
rect 488083 318218 508916 318454
rect 509152 318218 514847 318454
rect 515083 318218 535916 318454
rect 536152 318218 541847 318454
rect 542083 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 586302 318454
rect 586538 318218 586622 318454
rect 586858 318218 586890 318454
rect -2966 318134 586890 318218
rect -2966 317898 -2934 318134
rect -2698 317898 -2614 318134
rect -2378 317898 10826 318134
rect 11062 317898 11146 318134
rect 11382 317898 22916 318134
rect 23152 317898 28847 318134
rect 29083 317898 49916 318134
rect 50152 317898 55847 318134
rect 56083 317898 76916 318134
rect 77152 317898 82847 318134
rect 83083 317898 103916 318134
rect 104152 317898 109847 318134
rect 110083 317898 130916 318134
rect 131152 317898 136847 318134
rect 137083 317898 157916 318134
rect 158152 317898 163847 318134
rect 164083 317898 184916 318134
rect 185152 317898 190847 318134
rect 191083 317898 211916 318134
rect 212152 317898 217847 318134
rect 218083 317898 238916 318134
rect 239152 317898 244847 318134
rect 245083 317898 265916 318134
rect 266152 317898 271847 318134
rect 272083 317898 292916 318134
rect 293152 317898 298847 318134
rect 299083 317898 319916 318134
rect 320152 317898 325847 318134
rect 326083 317898 346916 318134
rect 347152 317898 352847 318134
rect 353083 317898 373916 318134
rect 374152 317898 379847 318134
rect 380083 317898 400916 318134
rect 401152 317898 406847 318134
rect 407083 317898 427916 318134
rect 428152 317898 433847 318134
rect 434083 317898 454916 318134
rect 455152 317898 460847 318134
rect 461083 317898 481916 318134
rect 482152 317898 487847 318134
rect 488083 317898 508916 318134
rect 509152 317898 514847 318134
rect 515083 317898 535916 318134
rect 536152 317898 541847 318134
rect 542083 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 586302 318134
rect 586538 317898 586622 318134
rect 586858 317898 586890 318134
rect -2966 317866 586890 317898
rect 28794 310394 551414 310426
rect 28794 310158 28826 310394
rect 29062 310158 29146 310394
rect 29382 310158 46826 310394
rect 47062 310158 47146 310394
rect 47382 310158 64826 310394
rect 65062 310158 65146 310394
rect 65382 310158 82826 310394
rect 83062 310158 83146 310394
rect 83382 310158 100826 310394
rect 101062 310158 101146 310394
rect 101382 310158 118826 310394
rect 119062 310158 119146 310394
rect 119382 310158 136826 310394
rect 137062 310158 137146 310394
rect 137382 310158 154826 310394
rect 155062 310158 155146 310394
rect 155382 310158 172826 310394
rect 173062 310158 173146 310394
rect 173382 310158 190826 310394
rect 191062 310158 191146 310394
rect 191382 310158 208826 310394
rect 209062 310158 209146 310394
rect 209382 310158 226826 310394
rect 227062 310158 227146 310394
rect 227382 310158 244826 310394
rect 245062 310158 245146 310394
rect 245382 310158 262826 310394
rect 263062 310158 263146 310394
rect 263382 310158 280826 310394
rect 281062 310158 281146 310394
rect 281382 310158 298826 310394
rect 299062 310158 299146 310394
rect 299382 310158 316826 310394
rect 317062 310158 317146 310394
rect 317382 310158 334826 310394
rect 335062 310158 335146 310394
rect 335382 310158 352826 310394
rect 353062 310158 353146 310394
rect 353382 310158 370826 310394
rect 371062 310158 371146 310394
rect 371382 310158 388826 310394
rect 389062 310158 389146 310394
rect 389382 310158 406826 310394
rect 407062 310158 407146 310394
rect 407382 310158 424826 310394
rect 425062 310158 425146 310394
rect 425382 310158 442826 310394
rect 443062 310158 443146 310394
rect 443382 310158 460826 310394
rect 461062 310158 461146 310394
rect 461382 310158 478826 310394
rect 479062 310158 479146 310394
rect 479382 310158 496826 310394
rect 497062 310158 497146 310394
rect 497382 310158 514826 310394
rect 515062 310158 515146 310394
rect 515382 310158 532826 310394
rect 533062 310158 533146 310394
rect 533382 310158 550826 310394
rect 551062 310158 551146 310394
rect 551382 310158 551414 310394
rect 28794 310074 551414 310158
rect 28794 309838 28826 310074
rect 29062 309838 29146 310074
rect 29382 309838 46826 310074
rect 47062 309838 47146 310074
rect 47382 309838 64826 310074
rect 65062 309838 65146 310074
rect 65382 309838 82826 310074
rect 83062 309838 83146 310074
rect 83382 309838 100826 310074
rect 101062 309838 101146 310074
rect 101382 309838 118826 310074
rect 119062 309838 119146 310074
rect 119382 309838 136826 310074
rect 137062 309838 137146 310074
rect 137382 309838 154826 310074
rect 155062 309838 155146 310074
rect 155382 309838 172826 310074
rect 173062 309838 173146 310074
rect 173382 309838 190826 310074
rect 191062 309838 191146 310074
rect 191382 309838 208826 310074
rect 209062 309838 209146 310074
rect 209382 309838 226826 310074
rect 227062 309838 227146 310074
rect 227382 309838 244826 310074
rect 245062 309838 245146 310074
rect 245382 309838 262826 310074
rect 263062 309838 263146 310074
rect 263382 309838 280826 310074
rect 281062 309838 281146 310074
rect 281382 309838 298826 310074
rect 299062 309838 299146 310074
rect 299382 309838 316826 310074
rect 317062 309838 317146 310074
rect 317382 309838 334826 310074
rect 335062 309838 335146 310074
rect 335382 309838 352826 310074
rect 353062 309838 353146 310074
rect 353382 309838 370826 310074
rect 371062 309838 371146 310074
rect 371382 309838 388826 310074
rect 389062 309838 389146 310074
rect 389382 309838 406826 310074
rect 407062 309838 407146 310074
rect 407382 309838 424826 310074
rect 425062 309838 425146 310074
rect 425382 309838 442826 310074
rect 443062 309838 443146 310074
rect 443382 309838 460826 310074
rect 461062 309838 461146 310074
rect 461382 309838 478826 310074
rect 479062 309838 479146 310074
rect 479382 309838 496826 310074
rect 497062 309838 497146 310074
rect 497382 309838 514826 310074
rect 515062 309838 515146 310074
rect 515382 309838 532826 310074
rect 533062 309838 533146 310074
rect 533382 309838 550826 310074
rect 551062 309838 551146 310074
rect 551382 309838 551414 310074
rect 28794 309806 551414 309838
rect -2966 309454 586890 309486
rect -2966 309218 -1974 309454
rect -1738 309218 -1654 309454
rect -1418 309218 1826 309454
rect 2062 309218 2146 309454
rect 2382 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 37826 309454
rect 38062 309218 38146 309454
rect 38382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 73826 309454
rect 74062 309218 74146 309454
rect 74382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 109826 309454
rect 110062 309218 110146 309454
rect 110382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 145826 309454
rect 146062 309218 146146 309454
rect 146382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 181826 309454
rect 182062 309218 182146 309454
rect 182382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 217826 309454
rect 218062 309218 218146 309454
rect 218382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 253826 309454
rect 254062 309218 254146 309454
rect 254382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 289826 309454
rect 290062 309218 290146 309454
rect 290382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 325826 309454
rect 326062 309218 326146 309454
rect 326382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 361826 309454
rect 362062 309218 362146 309454
rect 362382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 397826 309454
rect 398062 309218 398146 309454
rect 398382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 433826 309454
rect 434062 309218 434146 309454
rect 434382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 469826 309454
rect 470062 309218 470146 309454
rect 470382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 505826 309454
rect 506062 309218 506146 309454
rect 506382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 541826 309454
rect 542062 309218 542146 309454
rect 542382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 577826 309454
rect 578062 309218 578146 309454
rect 578382 309218 585342 309454
rect 585578 309218 585662 309454
rect 585898 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -1974 309134
rect -1738 308898 -1654 309134
rect -1418 308898 1826 309134
rect 2062 308898 2146 309134
rect 2382 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 37826 309134
rect 38062 308898 38146 309134
rect 38382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 73826 309134
rect 74062 308898 74146 309134
rect 74382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 109826 309134
rect 110062 308898 110146 309134
rect 110382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 145826 309134
rect 146062 308898 146146 309134
rect 146382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 181826 309134
rect 182062 308898 182146 309134
rect 182382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 217826 309134
rect 218062 308898 218146 309134
rect 218382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 253826 309134
rect 254062 308898 254146 309134
rect 254382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 289826 309134
rect 290062 308898 290146 309134
rect 290382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 325826 309134
rect 326062 308898 326146 309134
rect 326382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 361826 309134
rect 362062 308898 362146 309134
rect 362382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 397826 309134
rect 398062 308898 398146 309134
rect 398382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 433826 309134
rect 434062 308898 434146 309134
rect 434382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 469826 309134
rect 470062 308898 470146 309134
rect 470382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 505826 309134
rect 506062 308898 506146 309134
rect 506382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 541826 309134
rect 542062 308898 542146 309134
rect 542382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 577826 309134
rect 578062 308898 578146 309134
rect 578382 308898 585342 309134
rect 585578 308898 585662 309134
rect 585898 308898 586890 309134
rect -2966 308866 586890 308898
rect -2966 300454 586890 300486
rect -2966 300218 -2934 300454
rect -2698 300218 -2614 300454
rect -2378 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 22916 300454
rect 23152 300218 28847 300454
rect 29083 300218 49916 300454
rect 50152 300218 55847 300454
rect 56083 300218 76916 300454
rect 77152 300218 82847 300454
rect 83083 300218 103916 300454
rect 104152 300218 109847 300454
rect 110083 300218 130916 300454
rect 131152 300218 136847 300454
rect 137083 300218 157916 300454
rect 158152 300218 163847 300454
rect 164083 300218 184916 300454
rect 185152 300218 190847 300454
rect 191083 300218 211916 300454
rect 212152 300218 217847 300454
rect 218083 300218 238916 300454
rect 239152 300218 244847 300454
rect 245083 300218 265916 300454
rect 266152 300218 271847 300454
rect 272083 300218 292916 300454
rect 293152 300218 298847 300454
rect 299083 300218 319916 300454
rect 320152 300218 325847 300454
rect 326083 300218 346916 300454
rect 347152 300218 352847 300454
rect 353083 300218 373916 300454
rect 374152 300218 379847 300454
rect 380083 300218 400916 300454
rect 401152 300218 406847 300454
rect 407083 300218 427916 300454
rect 428152 300218 433847 300454
rect 434083 300218 454916 300454
rect 455152 300218 460847 300454
rect 461083 300218 481916 300454
rect 482152 300218 487847 300454
rect 488083 300218 508916 300454
rect 509152 300218 514847 300454
rect 515083 300218 535916 300454
rect 536152 300218 541847 300454
rect 542083 300218 568826 300454
rect 569062 300218 569146 300454
rect 569382 300218 586302 300454
rect 586538 300218 586622 300454
rect 586858 300218 586890 300454
rect -2966 300134 586890 300218
rect -2966 299898 -2934 300134
rect -2698 299898 -2614 300134
rect -2378 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 22916 300134
rect 23152 299898 28847 300134
rect 29083 299898 49916 300134
rect 50152 299898 55847 300134
rect 56083 299898 76916 300134
rect 77152 299898 82847 300134
rect 83083 299898 103916 300134
rect 104152 299898 109847 300134
rect 110083 299898 130916 300134
rect 131152 299898 136847 300134
rect 137083 299898 157916 300134
rect 158152 299898 163847 300134
rect 164083 299898 184916 300134
rect 185152 299898 190847 300134
rect 191083 299898 211916 300134
rect 212152 299898 217847 300134
rect 218083 299898 238916 300134
rect 239152 299898 244847 300134
rect 245083 299898 265916 300134
rect 266152 299898 271847 300134
rect 272083 299898 292916 300134
rect 293152 299898 298847 300134
rect 299083 299898 319916 300134
rect 320152 299898 325847 300134
rect 326083 299898 346916 300134
rect 347152 299898 352847 300134
rect 353083 299898 373916 300134
rect 374152 299898 379847 300134
rect 380083 299898 400916 300134
rect 401152 299898 406847 300134
rect 407083 299898 427916 300134
rect 428152 299898 433847 300134
rect 434083 299898 454916 300134
rect 455152 299898 460847 300134
rect 461083 299898 481916 300134
rect 482152 299898 487847 300134
rect 488083 299898 508916 300134
rect 509152 299898 514847 300134
rect 515083 299898 535916 300134
rect 536152 299898 541847 300134
rect 542083 299898 568826 300134
rect 569062 299898 569146 300134
rect 569382 299898 586302 300134
rect 586538 299898 586622 300134
rect 586858 299898 586890 300134
rect -2966 299866 586890 299898
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 19952 291454
rect 20188 291218 25882 291454
rect 26118 291218 31813 291454
rect 32049 291218 46952 291454
rect 47188 291218 52882 291454
rect 53118 291218 58813 291454
rect 59049 291218 73952 291454
rect 74188 291218 79882 291454
rect 80118 291218 85813 291454
rect 86049 291218 100952 291454
rect 101188 291218 106882 291454
rect 107118 291218 112813 291454
rect 113049 291218 127952 291454
rect 128188 291218 133882 291454
rect 134118 291218 139813 291454
rect 140049 291218 154952 291454
rect 155188 291218 160882 291454
rect 161118 291218 166813 291454
rect 167049 291218 181952 291454
rect 182188 291218 187882 291454
rect 188118 291218 193813 291454
rect 194049 291218 208952 291454
rect 209188 291218 214882 291454
rect 215118 291218 220813 291454
rect 221049 291218 235952 291454
rect 236188 291218 241882 291454
rect 242118 291218 247813 291454
rect 248049 291218 262952 291454
rect 263188 291218 268882 291454
rect 269118 291218 274813 291454
rect 275049 291218 289952 291454
rect 290188 291218 295882 291454
rect 296118 291218 301813 291454
rect 302049 291218 316952 291454
rect 317188 291218 322882 291454
rect 323118 291218 328813 291454
rect 329049 291218 343952 291454
rect 344188 291218 349882 291454
rect 350118 291218 355813 291454
rect 356049 291218 370952 291454
rect 371188 291218 376882 291454
rect 377118 291218 382813 291454
rect 383049 291218 397952 291454
rect 398188 291218 403882 291454
rect 404118 291218 409813 291454
rect 410049 291218 424952 291454
rect 425188 291218 430882 291454
rect 431118 291218 436813 291454
rect 437049 291218 451952 291454
rect 452188 291218 457882 291454
rect 458118 291218 463813 291454
rect 464049 291218 478952 291454
rect 479188 291218 484882 291454
rect 485118 291218 490813 291454
rect 491049 291218 505952 291454
rect 506188 291218 511882 291454
rect 512118 291218 517813 291454
rect 518049 291218 532952 291454
rect 533188 291218 538882 291454
rect 539118 291218 544813 291454
rect 545049 291218 559826 291454
rect 560062 291218 560146 291454
rect 560382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 19952 291134
rect 20188 290898 25882 291134
rect 26118 290898 31813 291134
rect 32049 290898 46952 291134
rect 47188 290898 52882 291134
rect 53118 290898 58813 291134
rect 59049 290898 73952 291134
rect 74188 290898 79882 291134
rect 80118 290898 85813 291134
rect 86049 290898 100952 291134
rect 101188 290898 106882 291134
rect 107118 290898 112813 291134
rect 113049 290898 127952 291134
rect 128188 290898 133882 291134
rect 134118 290898 139813 291134
rect 140049 290898 154952 291134
rect 155188 290898 160882 291134
rect 161118 290898 166813 291134
rect 167049 290898 181952 291134
rect 182188 290898 187882 291134
rect 188118 290898 193813 291134
rect 194049 290898 208952 291134
rect 209188 290898 214882 291134
rect 215118 290898 220813 291134
rect 221049 290898 235952 291134
rect 236188 290898 241882 291134
rect 242118 290898 247813 291134
rect 248049 290898 262952 291134
rect 263188 290898 268882 291134
rect 269118 290898 274813 291134
rect 275049 290898 289952 291134
rect 290188 290898 295882 291134
rect 296118 290898 301813 291134
rect 302049 290898 316952 291134
rect 317188 290898 322882 291134
rect 323118 290898 328813 291134
rect 329049 290898 343952 291134
rect 344188 290898 349882 291134
rect 350118 290898 355813 291134
rect 356049 290898 370952 291134
rect 371188 290898 376882 291134
rect 377118 290898 382813 291134
rect 383049 290898 397952 291134
rect 398188 290898 403882 291134
rect 404118 290898 409813 291134
rect 410049 290898 424952 291134
rect 425188 290898 430882 291134
rect 431118 290898 436813 291134
rect 437049 290898 451952 291134
rect 452188 290898 457882 291134
rect 458118 290898 463813 291134
rect 464049 290898 478952 291134
rect 479188 290898 484882 291134
rect 485118 290898 490813 291134
rect 491049 290898 505952 291134
rect 506188 290898 511882 291134
rect 512118 290898 517813 291134
rect 518049 290898 532952 291134
rect 533188 290898 538882 291134
rect 539118 290898 544813 291134
rect 545049 290898 559826 291134
rect 560062 290898 560146 291134
rect 560382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect 19794 283394 542414 283426
rect 19794 283158 19826 283394
rect 20062 283158 20146 283394
rect 20382 283158 37826 283394
rect 38062 283158 38146 283394
rect 38382 283158 55826 283394
rect 56062 283158 56146 283394
rect 56382 283158 73826 283394
rect 74062 283158 74146 283394
rect 74382 283158 91826 283394
rect 92062 283158 92146 283394
rect 92382 283158 109826 283394
rect 110062 283158 110146 283394
rect 110382 283158 127826 283394
rect 128062 283158 128146 283394
rect 128382 283158 145826 283394
rect 146062 283158 146146 283394
rect 146382 283158 163826 283394
rect 164062 283158 164146 283394
rect 164382 283158 181826 283394
rect 182062 283158 182146 283394
rect 182382 283158 199826 283394
rect 200062 283158 200146 283394
rect 200382 283158 217826 283394
rect 218062 283158 218146 283394
rect 218382 283158 235826 283394
rect 236062 283158 236146 283394
rect 236382 283158 253826 283394
rect 254062 283158 254146 283394
rect 254382 283158 271826 283394
rect 272062 283158 272146 283394
rect 272382 283158 289826 283394
rect 290062 283158 290146 283394
rect 290382 283158 307826 283394
rect 308062 283158 308146 283394
rect 308382 283158 325826 283394
rect 326062 283158 326146 283394
rect 326382 283158 343826 283394
rect 344062 283158 344146 283394
rect 344382 283158 361826 283394
rect 362062 283158 362146 283394
rect 362382 283158 379826 283394
rect 380062 283158 380146 283394
rect 380382 283158 397826 283394
rect 398062 283158 398146 283394
rect 398382 283158 415826 283394
rect 416062 283158 416146 283394
rect 416382 283158 433826 283394
rect 434062 283158 434146 283394
rect 434382 283158 451826 283394
rect 452062 283158 452146 283394
rect 452382 283158 469826 283394
rect 470062 283158 470146 283394
rect 470382 283158 487826 283394
rect 488062 283158 488146 283394
rect 488382 283158 505826 283394
rect 506062 283158 506146 283394
rect 506382 283158 523826 283394
rect 524062 283158 524146 283394
rect 524382 283158 541826 283394
rect 542062 283158 542146 283394
rect 542382 283158 542414 283394
rect 19794 283074 542414 283158
rect 19794 282838 19826 283074
rect 20062 282838 20146 283074
rect 20382 282838 37826 283074
rect 38062 282838 38146 283074
rect 38382 282838 55826 283074
rect 56062 282838 56146 283074
rect 56382 282838 73826 283074
rect 74062 282838 74146 283074
rect 74382 282838 91826 283074
rect 92062 282838 92146 283074
rect 92382 282838 109826 283074
rect 110062 282838 110146 283074
rect 110382 282838 127826 283074
rect 128062 282838 128146 283074
rect 128382 282838 145826 283074
rect 146062 282838 146146 283074
rect 146382 282838 163826 283074
rect 164062 282838 164146 283074
rect 164382 282838 181826 283074
rect 182062 282838 182146 283074
rect 182382 282838 199826 283074
rect 200062 282838 200146 283074
rect 200382 282838 217826 283074
rect 218062 282838 218146 283074
rect 218382 282838 235826 283074
rect 236062 282838 236146 283074
rect 236382 282838 253826 283074
rect 254062 282838 254146 283074
rect 254382 282838 271826 283074
rect 272062 282838 272146 283074
rect 272382 282838 289826 283074
rect 290062 282838 290146 283074
rect 290382 282838 307826 283074
rect 308062 282838 308146 283074
rect 308382 282838 325826 283074
rect 326062 282838 326146 283074
rect 326382 282838 343826 283074
rect 344062 282838 344146 283074
rect 344382 282838 361826 283074
rect 362062 282838 362146 283074
rect 362382 282838 379826 283074
rect 380062 282838 380146 283074
rect 380382 282838 397826 283074
rect 398062 282838 398146 283074
rect 398382 282838 415826 283074
rect 416062 282838 416146 283074
rect 416382 282838 433826 283074
rect 434062 282838 434146 283074
rect 434382 282838 451826 283074
rect 452062 282838 452146 283074
rect 452382 282838 469826 283074
rect 470062 282838 470146 283074
rect 470382 282838 487826 283074
rect 488062 282838 488146 283074
rect 488382 282838 505826 283074
rect 506062 282838 506146 283074
rect 506382 282838 523826 283074
rect 524062 282838 524146 283074
rect 524382 282838 541826 283074
rect 542062 282838 542146 283074
rect 542382 282838 542414 283074
rect 19794 282806 542414 282838
rect -2966 282454 586890 282486
rect -2966 282218 -2934 282454
rect -2698 282218 -2614 282454
rect -2378 282218 10826 282454
rect 11062 282218 11146 282454
rect 11382 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 46826 282454
rect 47062 282218 47146 282454
rect 47382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 82826 282454
rect 83062 282218 83146 282454
rect 83382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 118826 282454
rect 119062 282218 119146 282454
rect 119382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 154826 282454
rect 155062 282218 155146 282454
rect 155382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 190826 282454
rect 191062 282218 191146 282454
rect 191382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 226826 282454
rect 227062 282218 227146 282454
rect 227382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 262826 282454
rect 263062 282218 263146 282454
rect 263382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 298826 282454
rect 299062 282218 299146 282454
rect 299382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 334826 282454
rect 335062 282218 335146 282454
rect 335382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 370826 282454
rect 371062 282218 371146 282454
rect 371382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 406826 282454
rect 407062 282218 407146 282454
rect 407382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 442826 282454
rect 443062 282218 443146 282454
rect 443382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 478826 282454
rect 479062 282218 479146 282454
rect 479382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 514826 282454
rect 515062 282218 515146 282454
rect 515382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 550826 282454
rect 551062 282218 551146 282454
rect 551382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 586302 282454
rect 586538 282218 586622 282454
rect 586858 282218 586890 282454
rect -2966 282134 586890 282218
rect -2966 281898 -2934 282134
rect -2698 281898 -2614 282134
rect -2378 281898 10826 282134
rect 11062 281898 11146 282134
rect 11382 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 46826 282134
rect 47062 281898 47146 282134
rect 47382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 82826 282134
rect 83062 281898 83146 282134
rect 83382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 118826 282134
rect 119062 281898 119146 282134
rect 119382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 154826 282134
rect 155062 281898 155146 282134
rect 155382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 190826 282134
rect 191062 281898 191146 282134
rect 191382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 226826 282134
rect 227062 281898 227146 282134
rect 227382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 262826 282134
rect 263062 281898 263146 282134
rect 263382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 298826 282134
rect 299062 281898 299146 282134
rect 299382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 334826 282134
rect 335062 281898 335146 282134
rect 335382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 370826 282134
rect 371062 281898 371146 282134
rect 371382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 406826 282134
rect 407062 281898 407146 282134
rect 407382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 442826 282134
rect 443062 281898 443146 282134
rect 443382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 478826 282134
rect 479062 281898 479146 282134
rect 479382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 514826 282134
rect 515062 281898 515146 282134
rect 515382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 550826 282134
rect 551062 281898 551146 282134
rect 551382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 586302 282134
rect 586538 281898 586622 282134
rect 586858 281898 586890 282134
rect -2966 281866 586890 281898
rect -2966 273454 586890 273486
rect -2966 273218 -1974 273454
rect -1738 273218 -1654 273454
rect -1418 273218 1826 273454
rect 2062 273218 2146 273454
rect 2382 273218 19952 273454
rect 20188 273218 25882 273454
rect 26118 273218 31813 273454
rect 32049 273218 46952 273454
rect 47188 273218 52882 273454
rect 53118 273218 58813 273454
rect 59049 273218 73952 273454
rect 74188 273218 79882 273454
rect 80118 273218 85813 273454
rect 86049 273218 100952 273454
rect 101188 273218 106882 273454
rect 107118 273218 112813 273454
rect 113049 273218 127952 273454
rect 128188 273218 133882 273454
rect 134118 273218 139813 273454
rect 140049 273218 154952 273454
rect 155188 273218 160882 273454
rect 161118 273218 166813 273454
rect 167049 273218 181952 273454
rect 182188 273218 187882 273454
rect 188118 273218 193813 273454
rect 194049 273218 208952 273454
rect 209188 273218 214882 273454
rect 215118 273218 220813 273454
rect 221049 273218 235952 273454
rect 236188 273218 241882 273454
rect 242118 273218 247813 273454
rect 248049 273218 262952 273454
rect 263188 273218 268882 273454
rect 269118 273218 274813 273454
rect 275049 273218 289952 273454
rect 290188 273218 295882 273454
rect 296118 273218 301813 273454
rect 302049 273218 316952 273454
rect 317188 273218 322882 273454
rect 323118 273218 328813 273454
rect 329049 273218 343952 273454
rect 344188 273218 349882 273454
rect 350118 273218 355813 273454
rect 356049 273218 370952 273454
rect 371188 273218 376882 273454
rect 377118 273218 382813 273454
rect 383049 273218 397952 273454
rect 398188 273218 403882 273454
rect 404118 273218 409813 273454
rect 410049 273218 424952 273454
rect 425188 273218 430882 273454
rect 431118 273218 436813 273454
rect 437049 273218 451952 273454
rect 452188 273218 457882 273454
rect 458118 273218 463813 273454
rect 464049 273218 478952 273454
rect 479188 273218 484882 273454
rect 485118 273218 490813 273454
rect 491049 273218 505952 273454
rect 506188 273218 511882 273454
rect 512118 273218 517813 273454
rect 518049 273218 532952 273454
rect 533188 273218 538882 273454
rect 539118 273218 544813 273454
rect 545049 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 577826 273454
rect 578062 273218 578146 273454
rect 578382 273218 585342 273454
rect 585578 273218 585662 273454
rect 585898 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -1974 273134
rect -1738 272898 -1654 273134
rect -1418 272898 1826 273134
rect 2062 272898 2146 273134
rect 2382 272898 19952 273134
rect 20188 272898 25882 273134
rect 26118 272898 31813 273134
rect 32049 272898 46952 273134
rect 47188 272898 52882 273134
rect 53118 272898 58813 273134
rect 59049 272898 73952 273134
rect 74188 272898 79882 273134
rect 80118 272898 85813 273134
rect 86049 272898 100952 273134
rect 101188 272898 106882 273134
rect 107118 272898 112813 273134
rect 113049 272898 127952 273134
rect 128188 272898 133882 273134
rect 134118 272898 139813 273134
rect 140049 272898 154952 273134
rect 155188 272898 160882 273134
rect 161118 272898 166813 273134
rect 167049 272898 181952 273134
rect 182188 272898 187882 273134
rect 188118 272898 193813 273134
rect 194049 272898 208952 273134
rect 209188 272898 214882 273134
rect 215118 272898 220813 273134
rect 221049 272898 235952 273134
rect 236188 272898 241882 273134
rect 242118 272898 247813 273134
rect 248049 272898 262952 273134
rect 263188 272898 268882 273134
rect 269118 272898 274813 273134
rect 275049 272898 289952 273134
rect 290188 272898 295882 273134
rect 296118 272898 301813 273134
rect 302049 272898 316952 273134
rect 317188 272898 322882 273134
rect 323118 272898 328813 273134
rect 329049 272898 343952 273134
rect 344188 272898 349882 273134
rect 350118 272898 355813 273134
rect 356049 272898 370952 273134
rect 371188 272898 376882 273134
rect 377118 272898 382813 273134
rect 383049 272898 397952 273134
rect 398188 272898 403882 273134
rect 404118 272898 409813 273134
rect 410049 272898 424952 273134
rect 425188 272898 430882 273134
rect 431118 272898 436813 273134
rect 437049 272898 451952 273134
rect 452188 272898 457882 273134
rect 458118 272898 463813 273134
rect 464049 272898 478952 273134
rect 479188 272898 484882 273134
rect 485118 272898 490813 273134
rect 491049 272898 505952 273134
rect 506188 272898 511882 273134
rect 512118 272898 517813 273134
rect 518049 272898 532952 273134
rect 533188 272898 538882 273134
rect 539118 272898 544813 273134
rect 545049 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 577826 273134
rect 578062 272898 578146 273134
rect 578382 272898 585342 273134
rect 585578 272898 585662 273134
rect 585898 272898 586890 273134
rect -2966 272866 586890 272898
rect -2966 264454 586890 264486
rect -2966 264218 -2934 264454
rect -2698 264218 -2614 264454
rect -2378 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 22916 264454
rect 23152 264218 28847 264454
rect 29083 264218 49916 264454
rect 50152 264218 55847 264454
rect 56083 264218 76916 264454
rect 77152 264218 82847 264454
rect 83083 264218 103916 264454
rect 104152 264218 109847 264454
rect 110083 264218 130916 264454
rect 131152 264218 136847 264454
rect 137083 264218 157916 264454
rect 158152 264218 163847 264454
rect 164083 264218 184916 264454
rect 185152 264218 190847 264454
rect 191083 264218 211916 264454
rect 212152 264218 217847 264454
rect 218083 264218 238916 264454
rect 239152 264218 244847 264454
rect 245083 264218 265916 264454
rect 266152 264218 271847 264454
rect 272083 264218 292916 264454
rect 293152 264218 298847 264454
rect 299083 264218 319916 264454
rect 320152 264218 325847 264454
rect 326083 264218 346916 264454
rect 347152 264218 352847 264454
rect 353083 264218 373916 264454
rect 374152 264218 379847 264454
rect 380083 264218 400916 264454
rect 401152 264218 406847 264454
rect 407083 264218 427916 264454
rect 428152 264218 433847 264454
rect 434083 264218 454916 264454
rect 455152 264218 460847 264454
rect 461083 264218 481916 264454
rect 482152 264218 487847 264454
rect 488083 264218 508916 264454
rect 509152 264218 514847 264454
rect 515083 264218 535916 264454
rect 536152 264218 541847 264454
rect 542083 264218 568826 264454
rect 569062 264218 569146 264454
rect 569382 264218 586302 264454
rect 586538 264218 586622 264454
rect 586858 264218 586890 264454
rect -2966 264134 586890 264218
rect -2966 263898 -2934 264134
rect -2698 263898 -2614 264134
rect -2378 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 22916 264134
rect 23152 263898 28847 264134
rect 29083 263898 49916 264134
rect 50152 263898 55847 264134
rect 56083 263898 76916 264134
rect 77152 263898 82847 264134
rect 83083 263898 103916 264134
rect 104152 263898 109847 264134
rect 110083 263898 130916 264134
rect 131152 263898 136847 264134
rect 137083 263898 157916 264134
rect 158152 263898 163847 264134
rect 164083 263898 184916 264134
rect 185152 263898 190847 264134
rect 191083 263898 211916 264134
rect 212152 263898 217847 264134
rect 218083 263898 238916 264134
rect 239152 263898 244847 264134
rect 245083 263898 265916 264134
rect 266152 263898 271847 264134
rect 272083 263898 292916 264134
rect 293152 263898 298847 264134
rect 299083 263898 319916 264134
rect 320152 263898 325847 264134
rect 326083 263898 346916 264134
rect 347152 263898 352847 264134
rect 353083 263898 373916 264134
rect 374152 263898 379847 264134
rect 380083 263898 400916 264134
rect 401152 263898 406847 264134
rect 407083 263898 427916 264134
rect 428152 263898 433847 264134
rect 434083 263898 454916 264134
rect 455152 263898 460847 264134
rect 461083 263898 481916 264134
rect 482152 263898 487847 264134
rect 488083 263898 508916 264134
rect 509152 263898 514847 264134
rect 515083 263898 535916 264134
rect 536152 263898 541847 264134
rect 542083 263898 568826 264134
rect 569062 263898 569146 264134
rect 569382 263898 586302 264134
rect 586538 263898 586622 264134
rect 586858 263898 586890 264134
rect -2966 263866 586890 263898
rect 28794 256394 551414 256426
rect 28794 256158 28826 256394
rect 29062 256158 29146 256394
rect 29382 256158 46826 256394
rect 47062 256158 47146 256394
rect 47382 256158 64826 256394
rect 65062 256158 65146 256394
rect 65382 256158 82826 256394
rect 83062 256158 83146 256394
rect 83382 256158 100826 256394
rect 101062 256158 101146 256394
rect 101382 256158 118826 256394
rect 119062 256158 119146 256394
rect 119382 256158 136826 256394
rect 137062 256158 137146 256394
rect 137382 256158 154826 256394
rect 155062 256158 155146 256394
rect 155382 256158 172826 256394
rect 173062 256158 173146 256394
rect 173382 256158 190826 256394
rect 191062 256158 191146 256394
rect 191382 256158 208826 256394
rect 209062 256158 209146 256394
rect 209382 256158 226826 256394
rect 227062 256158 227146 256394
rect 227382 256158 244826 256394
rect 245062 256158 245146 256394
rect 245382 256158 262826 256394
rect 263062 256158 263146 256394
rect 263382 256158 280826 256394
rect 281062 256158 281146 256394
rect 281382 256158 298826 256394
rect 299062 256158 299146 256394
rect 299382 256158 316826 256394
rect 317062 256158 317146 256394
rect 317382 256158 334826 256394
rect 335062 256158 335146 256394
rect 335382 256158 352826 256394
rect 353062 256158 353146 256394
rect 353382 256158 370826 256394
rect 371062 256158 371146 256394
rect 371382 256158 388826 256394
rect 389062 256158 389146 256394
rect 389382 256158 406826 256394
rect 407062 256158 407146 256394
rect 407382 256158 424826 256394
rect 425062 256158 425146 256394
rect 425382 256158 442826 256394
rect 443062 256158 443146 256394
rect 443382 256158 460826 256394
rect 461062 256158 461146 256394
rect 461382 256158 478826 256394
rect 479062 256158 479146 256394
rect 479382 256158 496826 256394
rect 497062 256158 497146 256394
rect 497382 256158 514826 256394
rect 515062 256158 515146 256394
rect 515382 256158 532826 256394
rect 533062 256158 533146 256394
rect 533382 256158 550826 256394
rect 551062 256158 551146 256394
rect 551382 256158 551414 256394
rect 28794 256074 551414 256158
rect 28794 255838 28826 256074
rect 29062 255838 29146 256074
rect 29382 255838 46826 256074
rect 47062 255838 47146 256074
rect 47382 255838 64826 256074
rect 65062 255838 65146 256074
rect 65382 255838 82826 256074
rect 83062 255838 83146 256074
rect 83382 255838 100826 256074
rect 101062 255838 101146 256074
rect 101382 255838 118826 256074
rect 119062 255838 119146 256074
rect 119382 255838 136826 256074
rect 137062 255838 137146 256074
rect 137382 255838 154826 256074
rect 155062 255838 155146 256074
rect 155382 255838 172826 256074
rect 173062 255838 173146 256074
rect 173382 255838 190826 256074
rect 191062 255838 191146 256074
rect 191382 255838 208826 256074
rect 209062 255838 209146 256074
rect 209382 255838 226826 256074
rect 227062 255838 227146 256074
rect 227382 255838 244826 256074
rect 245062 255838 245146 256074
rect 245382 255838 262826 256074
rect 263062 255838 263146 256074
rect 263382 255838 280826 256074
rect 281062 255838 281146 256074
rect 281382 255838 298826 256074
rect 299062 255838 299146 256074
rect 299382 255838 316826 256074
rect 317062 255838 317146 256074
rect 317382 255838 334826 256074
rect 335062 255838 335146 256074
rect 335382 255838 352826 256074
rect 353062 255838 353146 256074
rect 353382 255838 370826 256074
rect 371062 255838 371146 256074
rect 371382 255838 388826 256074
rect 389062 255838 389146 256074
rect 389382 255838 406826 256074
rect 407062 255838 407146 256074
rect 407382 255838 424826 256074
rect 425062 255838 425146 256074
rect 425382 255838 442826 256074
rect 443062 255838 443146 256074
rect 443382 255838 460826 256074
rect 461062 255838 461146 256074
rect 461382 255838 478826 256074
rect 479062 255838 479146 256074
rect 479382 255838 496826 256074
rect 497062 255838 497146 256074
rect 497382 255838 514826 256074
rect 515062 255838 515146 256074
rect 515382 255838 532826 256074
rect 533062 255838 533146 256074
rect 533382 255838 550826 256074
rect 551062 255838 551146 256074
rect 551382 255838 551414 256074
rect 28794 255806 551414 255838
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 19826 255454
rect 20062 255218 20146 255454
rect 20382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 55826 255454
rect 56062 255218 56146 255454
rect 56382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 91826 255454
rect 92062 255218 92146 255454
rect 92382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 127826 255454
rect 128062 255218 128146 255454
rect 128382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 163826 255454
rect 164062 255218 164146 255454
rect 164382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 199826 255454
rect 200062 255218 200146 255454
rect 200382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 235826 255454
rect 236062 255218 236146 255454
rect 236382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 271826 255454
rect 272062 255218 272146 255454
rect 272382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 307826 255454
rect 308062 255218 308146 255454
rect 308382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 343826 255454
rect 344062 255218 344146 255454
rect 344382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 379826 255454
rect 380062 255218 380146 255454
rect 380382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 415826 255454
rect 416062 255218 416146 255454
rect 416382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 451826 255454
rect 452062 255218 452146 255454
rect 452382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 487826 255454
rect 488062 255218 488146 255454
rect 488382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 523826 255454
rect 524062 255218 524146 255454
rect 524382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 559826 255454
rect 560062 255218 560146 255454
rect 560382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 19826 255134
rect 20062 254898 20146 255134
rect 20382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 55826 255134
rect 56062 254898 56146 255134
rect 56382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 91826 255134
rect 92062 254898 92146 255134
rect 92382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 127826 255134
rect 128062 254898 128146 255134
rect 128382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 163826 255134
rect 164062 254898 164146 255134
rect 164382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 199826 255134
rect 200062 254898 200146 255134
rect 200382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 235826 255134
rect 236062 254898 236146 255134
rect 236382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 271826 255134
rect 272062 254898 272146 255134
rect 272382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 307826 255134
rect 308062 254898 308146 255134
rect 308382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 343826 255134
rect 344062 254898 344146 255134
rect 344382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 379826 255134
rect 380062 254898 380146 255134
rect 380382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 415826 255134
rect 416062 254898 416146 255134
rect 416382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 451826 255134
rect 452062 254898 452146 255134
rect 452382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 487826 255134
rect 488062 254898 488146 255134
rect 488382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 523826 255134
rect 524062 254898 524146 255134
rect 524382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 559826 255134
rect 560062 254898 560146 255134
rect 560382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -2966 246454 586890 246486
rect -2966 246218 -2934 246454
rect -2698 246218 -2614 246454
rect -2378 246218 10826 246454
rect 11062 246218 11146 246454
rect 11382 246218 22916 246454
rect 23152 246218 28847 246454
rect 29083 246218 49916 246454
rect 50152 246218 55847 246454
rect 56083 246218 76916 246454
rect 77152 246218 82847 246454
rect 83083 246218 103916 246454
rect 104152 246218 109847 246454
rect 110083 246218 130916 246454
rect 131152 246218 136847 246454
rect 137083 246218 157916 246454
rect 158152 246218 163847 246454
rect 164083 246218 184916 246454
rect 185152 246218 190847 246454
rect 191083 246218 211916 246454
rect 212152 246218 217847 246454
rect 218083 246218 238916 246454
rect 239152 246218 244847 246454
rect 245083 246218 265916 246454
rect 266152 246218 271847 246454
rect 272083 246218 292916 246454
rect 293152 246218 298847 246454
rect 299083 246218 319916 246454
rect 320152 246218 325847 246454
rect 326083 246218 346916 246454
rect 347152 246218 352847 246454
rect 353083 246218 373916 246454
rect 374152 246218 379847 246454
rect 380083 246218 400916 246454
rect 401152 246218 406847 246454
rect 407083 246218 427916 246454
rect 428152 246218 433847 246454
rect 434083 246218 454916 246454
rect 455152 246218 460847 246454
rect 461083 246218 481916 246454
rect 482152 246218 487847 246454
rect 488083 246218 508916 246454
rect 509152 246218 514847 246454
rect 515083 246218 535916 246454
rect 536152 246218 541847 246454
rect 542083 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 586302 246454
rect 586538 246218 586622 246454
rect 586858 246218 586890 246454
rect -2966 246134 586890 246218
rect -2966 245898 -2934 246134
rect -2698 245898 -2614 246134
rect -2378 245898 10826 246134
rect 11062 245898 11146 246134
rect 11382 245898 22916 246134
rect 23152 245898 28847 246134
rect 29083 245898 49916 246134
rect 50152 245898 55847 246134
rect 56083 245898 76916 246134
rect 77152 245898 82847 246134
rect 83083 245898 103916 246134
rect 104152 245898 109847 246134
rect 110083 245898 130916 246134
rect 131152 245898 136847 246134
rect 137083 245898 157916 246134
rect 158152 245898 163847 246134
rect 164083 245898 184916 246134
rect 185152 245898 190847 246134
rect 191083 245898 211916 246134
rect 212152 245898 217847 246134
rect 218083 245898 238916 246134
rect 239152 245898 244847 246134
rect 245083 245898 265916 246134
rect 266152 245898 271847 246134
rect 272083 245898 292916 246134
rect 293152 245898 298847 246134
rect 299083 245898 319916 246134
rect 320152 245898 325847 246134
rect 326083 245898 346916 246134
rect 347152 245898 352847 246134
rect 353083 245898 373916 246134
rect 374152 245898 379847 246134
rect 380083 245898 400916 246134
rect 401152 245898 406847 246134
rect 407083 245898 427916 246134
rect 428152 245898 433847 246134
rect 434083 245898 454916 246134
rect 455152 245898 460847 246134
rect 461083 245898 481916 246134
rect 482152 245898 487847 246134
rect 488083 245898 508916 246134
rect 509152 245898 514847 246134
rect 515083 245898 535916 246134
rect 536152 245898 541847 246134
rect 542083 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 586302 246134
rect 586538 245898 586622 246134
rect 586858 245898 586890 246134
rect -2966 245866 586890 245898
rect -2966 237454 586890 237486
rect -2966 237218 -1974 237454
rect -1738 237218 -1654 237454
rect -1418 237218 1826 237454
rect 2062 237218 2146 237454
rect 2382 237218 19952 237454
rect 20188 237218 25882 237454
rect 26118 237218 31813 237454
rect 32049 237218 46952 237454
rect 47188 237218 52882 237454
rect 53118 237218 58813 237454
rect 59049 237218 73952 237454
rect 74188 237218 79882 237454
rect 80118 237218 85813 237454
rect 86049 237218 100952 237454
rect 101188 237218 106882 237454
rect 107118 237218 112813 237454
rect 113049 237218 127952 237454
rect 128188 237218 133882 237454
rect 134118 237218 139813 237454
rect 140049 237218 154952 237454
rect 155188 237218 160882 237454
rect 161118 237218 166813 237454
rect 167049 237218 181952 237454
rect 182188 237218 187882 237454
rect 188118 237218 193813 237454
rect 194049 237218 208952 237454
rect 209188 237218 214882 237454
rect 215118 237218 220813 237454
rect 221049 237218 235952 237454
rect 236188 237218 241882 237454
rect 242118 237218 247813 237454
rect 248049 237218 262952 237454
rect 263188 237218 268882 237454
rect 269118 237218 274813 237454
rect 275049 237218 289952 237454
rect 290188 237218 295882 237454
rect 296118 237218 301813 237454
rect 302049 237218 316952 237454
rect 317188 237218 322882 237454
rect 323118 237218 328813 237454
rect 329049 237218 343952 237454
rect 344188 237218 349882 237454
rect 350118 237218 355813 237454
rect 356049 237218 370952 237454
rect 371188 237218 376882 237454
rect 377118 237218 382813 237454
rect 383049 237218 397952 237454
rect 398188 237218 403882 237454
rect 404118 237218 409813 237454
rect 410049 237218 424952 237454
rect 425188 237218 430882 237454
rect 431118 237218 436813 237454
rect 437049 237218 451952 237454
rect 452188 237218 457882 237454
rect 458118 237218 463813 237454
rect 464049 237218 478952 237454
rect 479188 237218 484882 237454
rect 485118 237218 490813 237454
rect 491049 237218 505952 237454
rect 506188 237218 511882 237454
rect 512118 237218 517813 237454
rect 518049 237218 532952 237454
rect 533188 237218 538882 237454
rect 539118 237218 544813 237454
rect 545049 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 577826 237454
rect 578062 237218 578146 237454
rect 578382 237218 585342 237454
rect 585578 237218 585662 237454
rect 585898 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -1974 237134
rect -1738 236898 -1654 237134
rect -1418 236898 1826 237134
rect 2062 236898 2146 237134
rect 2382 236898 19952 237134
rect 20188 236898 25882 237134
rect 26118 236898 31813 237134
rect 32049 236898 46952 237134
rect 47188 236898 52882 237134
rect 53118 236898 58813 237134
rect 59049 236898 73952 237134
rect 74188 236898 79882 237134
rect 80118 236898 85813 237134
rect 86049 236898 100952 237134
rect 101188 236898 106882 237134
rect 107118 236898 112813 237134
rect 113049 236898 127952 237134
rect 128188 236898 133882 237134
rect 134118 236898 139813 237134
rect 140049 236898 154952 237134
rect 155188 236898 160882 237134
rect 161118 236898 166813 237134
rect 167049 236898 181952 237134
rect 182188 236898 187882 237134
rect 188118 236898 193813 237134
rect 194049 236898 208952 237134
rect 209188 236898 214882 237134
rect 215118 236898 220813 237134
rect 221049 236898 235952 237134
rect 236188 236898 241882 237134
rect 242118 236898 247813 237134
rect 248049 236898 262952 237134
rect 263188 236898 268882 237134
rect 269118 236898 274813 237134
rect 275049 236898 289952 237134
rect 290188 236898 295882 237134
rect 296118 236898 301813 237134
rect 302049 236898 316952 237134
rect 317188 236898 322882 237134
rect 323118 236898 328813 237134
rect 329049 236898 343952 237134
rect 344188 236898 349882 237134
rect 350118 236898 355813 237134
rect 356049 236898 370952 237134
rect 371188 236898 376882 237134
rect 377118 236898 382813 237134
rect 383049 236898 397952 237134
rect 398188 236898 403882 237134
rect 404118 236898 409813 237134
rect 410049 236898 424952 237134
rect 425188 236898 430882 237134
rect 431118 236898 436813 237134
rect 437049 236898 451952 237134
rect 452188 236898 457882 237134
rect 458118 236898 463813 237134
rect 464049 236898 478952 237134
rect 479188 236898 484882 237134
rect 485118 236898 490813 237134
rect 491049 236898 505952 237134
rect 506188 236898 511882 237134
rect 512118 236898 517813 237134
rect 518049 236898 532952 237134
rect 533188 236898 538882 237134
rect 539118 236898 544813 237134
rect 545049 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 577826 237134
rect 578062 236898 578146 237134
rect 578382 236898 585342 237134
rect 585578 236898 585662 237134
rect 585898 236898 586890 237134
rect -2966 236866 586890 236898
rect 19794 229394 542414 229426
rect 19794 229158 19826 229394
rect 20062 229158 20146 229394
rect 20382 229158 37826 229394
rect 38062 229158 38146 229394
rect 38382 229158 55826 229394
rect 56062 229158 56146 229394
rect 56382 229158 73826 229394
rect 74062 229158 74146 229394
rect 74382 229158 91826 229394
rect 92062 229158 92146 229394
rect 92382 229158 109826 229394
rect 110062 229158 110146 229394
rect 110382 229158 127826 229394
rect 128062 229158 128146 229394
rect 128382 229158 145826 229394
rect 146062 229158 146146 229394
rect 146382 229158 163826 229394
rect 164062 229158 164146 229394
rect 164382 229158 181826 229394
rect 182062 229158 182146 229394
rect 182382 229158 199826 229394
rect 200062 229158 200146 229394
rect 200382 229158 217826 229394
rect 218062 229158 218146 229394
rect 218382 229158 235826 229394
rect 236062 229158 236146 229394
rect 236382 229158 253826 229394
rect 254062 229158 254146 229394
rect 254382 229158 271826 229394
rect 272062 229158 272146 229394
rect 272382 229158 289826 229394
rect 290062 229158 290146 229394
rect 290382 229158 307826 229394
rect 308062 229158 308146 229394
rect 308382 229158 325826 229394
rect 326062 229158 326146 229394
rect 326382 229158 343826 229394
rect 344062 229158 344146 229394
rect 344382 229158 361826 229394
rect 362062 229158 362146 229394
rect 362382 229158 379826 229394
rect 380062 229158 380146 229394
rect 380382 229158 397826 229394
rect 398062 229158 398146 229394
rect 398382 229158 415826 229394
rect 416062 229158 416146 229394
rect 416382 229158 433826 229394
rect 434062 229158 434146 229394
rect 434382 229158 451826 229394
rect 452062 229158 452146 229394
rect 452382 229158 469826 229394
rect 470062 229158 470146 229394
rect 470382 229158 487826 229394
rect 488062 229158 488146 229394
rect 488382 229158 505826 229394
rect 506062 229158 506146 229394
rect 506382 229158 523826 229394
rect 524062 229158 524146 229394
rect 524382 229158 541826 229394
rect 542062 229158 542146 229394
rect 542382 229158 542414 229394
rect 19794 229074 542414 229158
rect 19794 228838 19826 229074
rect 20062 228838 20146 229074
rect 20382 228838 37826 229074
rect 38062 228838 38146 229074
rect 38382 228838 55826 229074
rect 56062 228838 56146 229074
rect 56382 228838 73826 229074
rect 74062 228838 74146 229074
rect 74382 228838 91826 229074
rect 92062 228838 92146 229074
rect 92382 228838 109826 229074
rect 110062 228838 110146 229074
rect 110382 228838 127826 229074
rect 128062 228838 128146 229074
rect 128382 228838 145826 229074
rect 146062 228838 146146 229074
rect 146382 228838 163826 229074
rect 164062 228838 164146 229074
rect 164382 228838 181826 229074
rect 182062 228838 182146 229074
rect 182382 228838 199826 229074
rect 200062 228838 200146 229074
rect 200382 228838 217826 229074
rect 218062 228838 218146 229074
rect 218382 228838 235826 229074
rect 236062 228838 236146 229074
rect 236382 228838 253826 229074
rect 254062 228838 254146 229074
rect 254382 228838 271826 229074
rect 272062 228838 272146 229074
rect 272382 228838 289826 229074
rect 290062 228838 290146 229074
rect 290382 228838 307826 229074
rect 308062 228838 308146 229074
rect 308382 228838 325826 229074
rect 326062 228838 326146 229074
rect 326382 228838 343826 229074
rect 344062 228838 344146 229074
rect 344382 228838 361826 229074
rect 362062 228838 362146 229074
rect 362382 228838 379826 229074
rect 380062 228838 380146 229074
rect 380382 228838 397826 229074
rect 398062 228838 398146 229074
rect 398382 228838 415826 229074
rect 416062 228838 416146 229074
rect 416382 228838 433826 229074
rect 434062 228838 434146 229074
rect 434382 228838 451826 229074
rect 452062 228838 452146 229074
rect 452382 228838 469826 229074
rect 470062 228838 470146 229074
rect 470382 228838 487826 229074
rect 488062 228838 488146 229074
rect 488382 228838 505826 229074
rect 506062 228838 506146 229074
rect 506382 228838 523826 229074
rect 524062 228838 524146 229074
rect 524382 228838 541826 229074
rect 542062 228838 542146 229074
rect 542382 228838 542414 229074
rect 19794 228806 542414 228838
rect -2966 228454 586890 228486
rect -2966 228218 -2934 228454
rect -2698 228218 -2614 228454
rect -2378 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 28826 228454
rect 29062 228218 29146 228454
rect 29382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 64826 228454
rect 65062 228218 65146 228454
rect 65382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 100826 228454
rect 101062 228218 101146 228454
rect 101382 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 136826 228454
rect 137062 228218 137146 228454
rect 137382 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 172826 228454
rect 173062 228218 173146 228454
rect 173382 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 208826 228454
rect 209062 228218 209146 228454
rect 209382 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 244826 228454
rect 245062 228218 245146 228454
rect 245382 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 280826 228454
rect 281062 228218 281146 228454
rect 281382 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 316826 228454
rect 317062 228218 317146 228454
rect 317382 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 352826 228454
rect 353062 228218 353146 228454
rect 353382 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 388826 228454
rect 389062 228218 389146 228454
rect 389382 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 424826 228454
rect 425062 228218 425146 228454
rect 425382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 460826 228454
rect 461062 228218 461146 228454
rect 461382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 496826 228454
rect 497062 228218 497146 228454
rect 497382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 532826 228454
rect 533062 228218 533146 228454
rect 533382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 568826 228454
rect 569062 228218 569146 228454
rect 569382 228218 586302 228454
rect 586538 228218 586622 228454
rect 586858 228218 586890 228454
rect -2966 228134 586890 228218
rect -2966 227898 -2934 228134
rect -2698 227898 -2614 228134
rect -2378 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 28826 228134
rect 29062 227898 29146 228134
rect 29382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 64826 228134
rect 65062 227898 65146 228134
rect 65382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 100826 228134
rect 101062 227898 101146 228134
rect 101382 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 136826 228134
rect 137062 227898 137146 228134
rect 137382 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 172826 228134
rect 173062 227898 173146 228134
rect 173382 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 208826 228134
rect 209062 227898 209146 228134
rect 209382 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 244826 228134
rect 245062 227898 245146 228134
rect 245382 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 280826 228134
rect 281062 227898 281146 228134
rect 281382 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 316826 228134
rect 317062 227898 317146 228134
rect 317382 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 352826 228134
rect 353062 227898 353146 228134
rect 353382 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 388826 228134
rect 389062 227898 389146 228134
rect 389382 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 424826 228134
rect 425062 227898 425146 228134
rect 425382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 460826 228134
rect 461062 227898 461146 228134
rect 461382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 496826 228134
rect 497062 227898 497146 228134
rect 497382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 532826 228134
rect 533062 227898 533146 228134
rect 533382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 568826 228134
rect 569062 227898 569146 228134
rect 569382 227898 586302 228134
rect 586538 227898 586622 228134
rect 586858 227898 586890 228134
rect -2966 227866 586890 227898
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 19952 219454
rect 20188 219218 25882 219454
rect 26118 219218 31813 219454
rect 32049 219218 46952 219454
rect 47188 219218 52882 219454
rect 53118 219218 58813 219454
rect 59049 219218 73952 219454
rect 74188 219218 79882 219454
rect 80118 219218 85813 219454
rect 86049 219218 100952 219454
rect 101188 219218 106882 219454
rect 107118 219218 112813 219454
rect 113049 219218 127952 219454
rect 128188 219218 133882 219454
rect 134118 219218 139813 219454
rect 140049 219218 154952 219454
rect 155188 219218 160882 219454
rect 161118 219218 166813 219454
rect 167049 219218 181952 219454
rect 182188 219218 187882 219454
rect 188118 219218 193813 219454
rect 194049 219218 208952 219454
rect 209188 219218 214882 219454
rect 215118 219218 220813 219454
rect 221049 219218 235952 219454
rect 236188 219218 241882 219454
rect 242118 219218 247813 219454
rect 248049 219218 262952 219454
rect 263188 219218 268882 219454
rect 269118 219218 274813 219454
rect 275049 219218 289952 219454
rect 290188 219218 295882 219454
rect 296118 219218 301813 219454
rect 302049 219218 316952 219454
rect 317188 219218 322882 219454
rect 323118 219218 328813 219454
rect 329049 219218 343952 219454
rect 344188 219218 349882 219454
rect 350118 219218 355813 219454
rect 356049 219218 370952 219454
rect 371188 219218 376882 219454
rect 377118 219218 382813 219454
rect 383049 219218 397952 219454
rect 398188 219218 403882 219454
rect 404118 219218 409813 219454
rect 410049 219218 424952 219454
rect 425188 219218 430882 219454
rect 431118 219218 436813 219454
rect 437049 219218 451952 219454
rect 452188 219218 457882 219454
rect 458118 219218 463813 219454
rect 464049 219218 478952 219454
rect 479188 219218 484882 219454
rect 485118 219218 490813 219454
rect 491049 219218 505952 219454
rect 506188 219218 511882 219454
rect 512118 219218 517813 219454
rect 518049 219218 532952 219454
rect 533188 219218 538882 219454
rect 539118 219218 544813 219454
rect 545049 219218 559826 219454
rect 560062 219218 560146 219454
rect 560382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 19952 219134
rect 20188 218898 25882 219134
rect 26118 218898 31813 219134
rect 32049 218898 46952 219134
rect 47188 218898 52882 219134
rect 53118 218898 58813 219134
rect 59049 218898 73952 219134
rect 74188 218898 79882 219134
rect 80118 218898 85813 219134
rect 86049 218898 100952 219134
rect 101188 218898 106882 219134
rect 107118 218898 112813 219134
rect 113049 218898 127952 219134
rect 128188 218898 133882 219134
rect 134118 218898 139813 219134
rect 140049 218898 154952 219134
rect 155188 218898 160882 219134
rect 161118 218898 166813 219134
rect 167049 218898 181952 219134
rect 182188 218898 187882 219134
rect 188118 218898 193813 219134
rect 194049 218898 208952 219134
rect 209188 218898 214882 219134
rect 215118 218898 220813 219134
rect 221049 218898 235952 219134
rect 236188 218898 241882 219134
rect 242118 218898 247813 219134
rect 248049 218898 262952 219134
rect 263188 218898 268882 219134
rect 269118 218898 274813 219134
rect 275049 218898 289952 219134
rect 290188 218898 295882 219134
rect 296118 218898 301813 219134
rect 302049 218898 316952 219134
rect 317188 218898 322882 219134
rect 323118 218898 328813 219134
rect 329049 218898 343952 219134
rect 344188 218898 349882 219134
rect 350118 218898 355813 219134
rect 356049 218898 370952 219134
rect 371188 218898 376882 219134
rect 377118 218898 382813 219134
rect 383049 218898 397952 219134
rect 398188 218898 403882 219134
rect 404118 218898 409813 219134
rect 410049 218898 424952 219134
rect 425188 218898 430882 219134
rect 431118 218898 436813 219134
rect 437049 218898 451952 219134
rect 452188 218898 457882 219134
rect 458118 218898 463813 219134
rect 464049 218898 478952 219134
rect 479188 218898 484882 219134
rect 485118 218898 490813 219134
rect 491049 218898 505952 219134
rect 506188 218898 511882 219134
rect 512118 218898 517813 219134
rect 518049 218898 532952 219134
rect 533188 218898 538882 219134
rect 539118 218898 544813 219134
rect 545049 218898 559826 219134
rect 560062 218898 560146 219134
rect 560382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -2966 210454 586890 210486
rect -2966 210218 -2934 210454
rect -2698 210218 -2614 210454
rect -2378 210218 10826 210454
rect 11062 210218 11146 210454
rect 11382 210218 22916 210454
rect 23152 210218 28847 210454
rect 29083 210218 49916 210454
rect 50152 210218 55847 210454
rect 56083 210218 76916 210454
rect 77152 210218 82847 210454
rect 83083 210218 103916 210454
rect 104152 210218 109847 210454
rect 110083 210218 130916 210454
rect 131152 210218 136847 210454
rect 137083 210218 157916 210454
rect 158152 210218 163847 210454
rect 164083 210218 184916 210454
rect 185152 210218 190847 210454
rect 191083 210218 211916 210454
rect 212152 210218 217847 210454
rect 218083 210218 238916 210454
rect 239152 210218 244847 210454
rect 245083 210218 265916 210454
rect 266152 210218 271847 210454
rect 272083 210218 292916 210454
rect 293152 210218 298847 210454
rect 299083 210218 319916 210454
rect 320152 210218 325847 210454
rect 326083 210218 346916 210454
rect 347152 210218 352847 210454
rect 353083 210218 373916 210454
rect 374152 210218 379847 210454
rect 380083 210218 400916 210454
rect 401152 210218 406847 210454
rect 407083 210218 427916 210454
rect 428152 210218 433847 210454
rect 434083 210218 454916 210454
rect 455152 210218 460847 210454
rect 461083 210218 481916 210454
rect 482152 210218 487847 210454
rect 488083 210218 508916 210454
rect 509152 210218 514847 210454
rect 515083 210218 535916 210454
rect 536152 210218 541847 210454
rect 542083 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 586302 210454
rect 586538 210218 586622 210454
rect 586858 210218 586890 210454
rect -2966 210134 586890 210218
rect -2966 209898 -2934 210134
rect -2698 209898 -2614 210134
rect -2378 209898 10826 210134
rect 11062 209898 11146 210134
rect 11382 209898 22916 210134
rect 23152 209898 28847 210134
rect 29083 209898 49916 210134
rect 50152 209898 55847 210134
rect 56083 209898 76916 210134
rect 77152 209898 82847 210134
rect 83083 209898 103916 210134
rect 104152 209898 109847 210134
rect 110083 209898 130916 210134
rect 131152 209898 136847 210134
rect 137083 209898 157916 210134
rect 158152 209898 163847 210134
rect 164083 209898 184916 210134
rect 185152 209898 190847 210134
rect 191083 209898 211916 210134
rect 212152 209898 217847 210134
rect 218083 209898 238916 210134
rect 239152 209898 244847 210134
rect 245083 209898 265916 210134
rect 266152 209898 271847 210134
rect 272083 209898 292916 210134
rect 293152 209898 298847 210134
rect 299083 209898 319916 210134
rect 320152 209898 325847 210134
rect 326083 209898 346916 210134
rect 347152 209898 352847 210134
rect 353083 209898 373916 210134
rect 374152 209898 379847 210134
rect 380083 209898 400916 210134
rect 401152 209898 406847 210134
rect 407083 209898 427916 210134
rect 428152 209898 433847 210134
rect 434083 209898 454916 210134
rect 455152 209898 460847 210134
rect 461083 209898 481916 210134
rect 482152 209898 487847 210134
rect 488083 209898 508916 210134
rect 509152 209898 514847 210134
rect 515083 209898 535916 210134
rect 536152 209898 541847 210134
rect 542083 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 586302 210134
rect 586538 209898 586622 210134
rect 586858 209898 586890 210134
rect -2966 209866 586890 209898
rect 28794 202394 551414 202426
rect 28794 202158 28826 202394
rect 29062 202158 29146 202394
rect 29382 202158 46826 202394
rect 47062 202158 47146 202394
rect 47382 202158 64826 202394
rect 65062 202158 65146 202394
rect 65382 202158 82826 202394
rect 83062 202158 83146 202394
rect 83382 202158 100826 202394
rect 101062 202158 101146 202394
rect 101382 202158 118826 202394
rect 119062 202158 119146 202394
rect 119382 202158 136826 202394
rect 137062 202158 137146 202394
rect 137382 202158 154826 202394
rect 155062 202158 155146 202394
rect 155382 202158 172826 202394
rect 173062 202158 173146 202394
rect 173382 202158 190826 202394
rect 191062 202158 191146 202394
rect 191382 202158 208826 202394
rect 209062 202158 209146 202394
rect 209382 202158 226826 202394
rect 227062 202158 227146 202394
rect 227382 202158 244826 202394
rect 245062 202158 245146 202394
rect 245382 202158 262826 202394
rect 263062 202158 263146 202394
rect 263382 202158 280826 202394
rect 281062 202158 281146 202394
rect 281382 202158 298826 202394
rect 299062 202158 299146 202394
rect 299382 202158 316826 202394
rect 317062 202158 317146 202394
rect 317382 202158 334826 202394
rect 335062 202158 335146 202394
rect 335382 202158 352826 202394
rect 353062 202158 353146 202394
rect 353382 202158 370826 202394
rect 371062 202158 371146 202394
rect 371382 202158 388826 202394
rect 389062 202158 389146 202394
rect 389382 202158 406826 202394
rect 407062 202158 407146 202394
rect 407382 202158 424826 202394
rect 425062 202158 425146 202394
rect 425382 202158 442826 202394
rect 443062 202158 443146 202394
rect 443382 202158 460826 202394
rect 461062 202158 461146 202394
rect 461382 202158 478826 202394
rect 479062 202158 479146 202394
rect 479382 202158 496826 202394
rect 497062 202158 497146 202394
rect 497382 202158 514826 202394
rect 515062 202158 515146 202394
rect 515382 202158 532826 202394
rect 533062 202158 533146 202394
rect 533382 202158 550826 202394
rect 551062 202158 551146 202394
rect 551382 202158 551414 202394
rect 28794 202074 551414 202158
rect 28794 201838 28826 202074
rect 29062 201838 29146 202074
rect 29382 201838 46826 202074
rect 47062 201838 47146 202074
rect 47382 201838 64826 202074
rect 65062 201838 65146 202074
rect 65382 201838 82826 202074
rect 83062 201838 83146 202074
rect 83382 201838 100826 202074
rect 101062 201838 101146 202074
rect 101382 201838 118826 202074
rect 119062 201838 119146 202074
rect 119382 201838 136826 202074
rect 137062 201838 137146 202074
rect 137382 201838 154826 202074
rect 155062 201838 155146 202074
rect 155382 201838 172826 202074
rect 173062 201838 173146 202074
rect 173382 201838 190826 202074
rect 191062 201838 191146 202074
rect 191382 201838 208826 202074
rect 209062 201838 209146 202074
rect 209382 201838 226826 202074
rect 227062 201838 227146 202074
rect 227382 201838 244826 202074
rect 245062 201838 245146 202074
rect 245382 201838 262826 202074
rect 263062 201838 263146 202074
rect 263382 201838 280826 202074
rect 281062 201838 281146 202074
rect 281382 201838 298826 202074
rect 299062 201838 299146 202074
rect 299382 201838 316826 202074
rect 317062 201838 317146 202074
rect 317382 201838 334826 202074
rect 335062 201838 335146 202074
rect 335382 201838 352826 202074
rect 353062 201838 353146 202074
rect 353382 201838 370826 202074
rect 371062 201838 371146 202074
rect 371382 201838 388826 202074
rect 389062 201838 389146 202074
rect 389382 201838 406826 202074
rect 407062 201838 407146 202074
rect 407382 201838 424826 202074
rect 425062 201838 425146 202074
rect 425382 201838 442826 202074
rect 443062 201838 443146 202074
rect 443382 201838 460826 202074
rect 461062 201838 461146 202074
rect 461382 201838 478826 202074
rect 479062 201838 479146 202074
rect 479382 201838 496826 202074
rect 497062 201838 497146 202074
rect 497382 201838 514826 202074
rect 515062 201838 515146 202074
rect 515382 201838 532826 202074
rect 533062 201838 533146 202074
rect 533382 201838 550826 202074
rect 551062 201838 551146 202074
rect 551382 201838 551414 202074
rect 28794 201806 551414 201838
rect -2966 201454 586890 201486
rect -2966 201218 -1974 201454
rect -1738 201218 -1654 201454
rect -1418 201218 1826 201454
rect 2062 201218 2146 201454
rect 2382 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 37826 201454
rect 38062 201218 38146 201454
rect 38382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 73826 201454
rect 74062 201218 74146 201454
rect 74382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 109826 201454
rect 110062 201218 110146 201454
rect 110382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 145826 201454
rect 146062 201218 146146 201454
rect 146382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 181826 201454
rect 182062 201218 182146 201454
rect 182382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 217826 201454
rect 218062 201218 218146 201454
rect 218382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 253826 201454
rect 254062 201218 254146 201454
rect 254382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 289826 201454
rect 290062 201218 290146 201454
rect 290382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 325826 201454
rect 326062 201218 326146 201454
rect 326382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 361826 201454
rect 362062 201218 362146 201454
rect 362382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 397826 201454
rect 398062 201218 398146 201454
rect 398382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 433826 201454
rect 434062 201218 434146 201454
rect 434382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 469826 201454
rect 470062 201218 470146 201454
rect 470382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 505826 201454
rect 506062 201218 506146 201454
rect 506382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 541826 201454
rect 542062 201218 542146 201454
rect 542382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 577826 201454
rect 578062 201218 578146 201454
rect 578382 201218 585342 201454
rect 585578 201218 585662 201454
rect 585898 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -1974 201134
rect -1738 200898 -1654 201134
rect -1418 200898 1826 201134
rect 2062 200898 2146 201134
rect 2382 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 37826 201134
rect 38062 200898 38146 201134
rect 38382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 73826 201134
rect 74062 200898 74146 201134
rect 74382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 109826 201134
rect 110062 200898 110146 201134
rect 110382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 145826 201134
rect 146062 200898 146146 201134
rect 146382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 181826 201134
rect 182062 200898 182146 201134
rect 182382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 217826 201134
rect 218062 200898 218146 201134
rect 218382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 253826 201134
rect 254062 200898 254146 201134
rect 254382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 289826 201134
rect 290062 200898 290146 201134
rect 290382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 325826 201134
rect 326062 200898 326146 201134
rect 326382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 361826 201134
rect 362062 200898 362146 201134
rect 362382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 397826 201134
rect 398062 200898 398146 201134
rect 398382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 433826 201134
rect 434062 200898 434146 201134
rect 434382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 469826 201134
rect 470062 200898 470146 201134
rect 470382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 505826 201134
rect 506062 200898 506146 201134
rect 506382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 541826 201134
rect 542062 200898 542146 201134
rect 542382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 577826 201134
rect 578062 200898 578146 201134
rect 578382 200898 585342 201134
rect 585578 200898 585662 201134
rect 585898 200898 586890 201134
rect -2966 200866 586890 200898
rect -2966 192454 586890 192486
rect -2966 192218 -2934 192454
rect -2698 192218 -2614 192454
rect -2378 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 22916 192454
rect 23152 192218 28847 192454
rect 29083 192218 49916 192454
rect 50152 192218 55847 192454
rect 56083 192218 76916 192454
rect 77152 192218 82847 192454
rect 83083 192218 103916 192454
rect 104152 192218 109847 192454
rect 110083 192218 130916 192454
rect 131152 192218 136847 192454
rect 137083 192218 157916 192454
rect 158152 192218 163847 192454
rect 164083 192218 184916 192454
rect 185152 192218 190847 192454
rect 191083 192218 211916 192454
rect 212152 192218 217847 192454
rect 218083 192218 238916 192454
rect 239152 192218 244847 192454
rect 245083 192218 265916 192454
rect 266152 192218 271847 192454
rect 272083 192218 292916 192454
rect 293152 192218 298847 192454
rect 299083 192218 319916 192454
rect 320152 192218 325847 192454
rect 326083 192218 346916 192454
rect 347152 192218 352847 192454
rect 353083 192218 373916 192454
rect 374152 192218 379847 192454
rect 380083 192218 400916 192454
rect 401152 192218 406847 192454
rect 407083 192218 427916 192454
rect 428152 192218 433847 192454
rect 434083 192218 454916 192454
rect 455152 192218 460847 192454
rect 461083 192218 481916 192454
rect 482152 192218 487847 192454
rect 488083 192218 508916 192454
rect 509152 192218 514847 192454
rect 515083 192218 535916 192454
rect 536152 192218 541847 192454
rect 542083 192218 568826 192454
rect 569062 192218 569146 192454
rect 569382 192218 586302 192454
rect 586538 192218 586622 192454
rect 586858 192218 586890 192454
rect -2966 192134 586890 192218
rect -2966 191898 -2934 192134
rect -2698 191898 -2614 192134
rect -2378 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 22916 192134
rect 23152 191898 28847 192134
rect 29083 191898 49916 192134
rect 50152 191898 55847 192134
rect 56083 191898 76916 192134
rect 77152 191898 82847 192134
rect 83083 191898 103916 192134
rect 104152 191898 109847 192134
rect 110083 191898 130916 192134
rect 131152 191898 136847 192134
rect 137083 191898 157916 192134
rect 158152 191898 163847 192134
rect 164083 191898 184916 192134
rect 185152 191898 190847 192134
rect 191083 191898 211916 192134
rect 212152 191898 217847 192134
rect 218083 191898 238916 192134
rect 239152 191898 244847 192134
rect 245083 191898 265916 192134
rect 266152 191898 271847 192134
rect 272083 191898 292916 192134
rect 293152 191898 298847 192134
rect 299083 191898 319916 192134
rect 320152 191898 325847 192134
rect 326083 191898 346916 192134
rect 347152 191898 352847 192134
rect 353083 191898 373916 192134
rect 374152 191898 379847 192134
rect 380083 191898 400916 192134
rect 401152 191898 406847 192134
rect 407083 191898 427916 192134
rect 428152 191898 433847 192134
rect 434083 191898 454916 192134
rect 455152 191898 460847 192134
rect 461083 191898 481916 192134
rect 482152 191898 487847 192134
rect 488083 191898 508916 192134
rect 509152 191898 514847 192134
rect 515083 191898 535916 192134
rect 536152 191898 541847 192134
rect 542083 191898 568826 192134
rect 569062 191898 569146 192134
rect 569382 191898 586302 192134
rect 586538 191898 586622 192134
rect 586858 191898 586890 192134
rect -2966 191866 586890 191898
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 19952 183454
rect 20188 183218 25882 183454
rect 26118 183218 31813 183454
rect 32049 183218 46952 183454
rect 47188 183218 52882 183454
rect 53118 183218 58813 183454
rect 59049 183218 73952 183454
rect 74188 183218 79882 183454
rect 80118 183218 85813 183454
rect 86049 183218 100952 183454
rect 101188 183218 106882 183454
rect 107118 183218 112813 183454
rect 113049 183218 127952 183454
rect 128188 183218 133882 183454
rect 134118 183218 139813 183454
rect 140049 183218 154952 183454
rect 155188 183218 160882 183454
rect 161118 183218 166813 183454
rect 167049 183218 181952 183454
rect 182188 183218 187882 183454
rect 188118 183218 193813 183454
rect 194049 183218 208952 183454
rect 209188 183218 214882 183454
rect 215118 183218 220813 183454
rect 221049 183218 235952 183454
rect 236188 183218 241882 183454
rect 242118 183218 247813 183454
rect 248049 183218 262952 183454
rect 263188 183218 268882 183454
rect 269118 183218 274813 183454
rect 275049 183218 289952 183454
rect 290188 183218 295882 183454
rect 296118 183218 301813 183454
rect 302049 183218 316952 183454
rect 317188 183218 322882 183454
rect 323118 183218 328813 183454
rect 329049 183218 343952 183454
rect 344188 183218 349882 183454
rect 350118 183218 355813 183454
rect 356049 183218 370952 183454
rect 371188 183218 376882 183454
rect 377118 183218 382813 183454
rect 383049 183218 397952 183454
rect 398188 183218 403882 183454
rect 404118 183218 409813 183454
rect 410049 183218 424952 183454
rect 425188 183218 430882 183454
rect 431118 183218 436813 183454
rect 437049 183218 451952 183454
rect 452188 183218 457882 183454
rect 458118 183218 463813 183454
rect 464049 183218 478952 183454
rect 479188 183218 484882 183454
rect 485118 183218 490813 183454
rect 491049 183218 505952 183454
rect 506188 183218 511882 183454
rect 512118 183218 517813 183454
rect 518049 183218 532952 183454
rect 533188 183218 538882 183454
rect 539118 183218 544813 183454
rect 545049 183218 559826 183454
rect 560062 183218 560146 183454
rect 560382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 19952 183134
rect 20188 182898 25882 183134
rect 26118 182898 31813 183134
rect 32049 182898 46952 183134
rect 47188 182898 52882 183134
rect 53118 182898 58813 183134
rect 59049 182898 73952 183134
rect 74188 182898 79882 183134
rect 80118 182898 85813 183134
rect 86049 182898 100952 183134
rect 101188 182898 106882 183134
rect 107118 182898 112813 183134
rect 113049 182898 127952 183134
rect 128188 182898 133882 183134
rect 134118 182898 139813 183134
rect 140049 182898 154952 183134
rect 155188 182898 160882 183134
rect 161118 182898 166813 183134
rect 167049 182898 181952 183134
rect 182188 182898 187882 183134
rect 188118 182898 193813 183134
rect 194049 182898 208952 183134
rect 209188 182898 214882 183134
rect 215118 182898 220813 183134
rect 221049 182898 235952 183134
rect 236188 182898 241882 183134
rect 242118 182898 247813 183134
rect 248049 182898 262952 183134
rect 263188 182898 268882 183134
rect 269118 182898 274813 183134
rect 275049 182898 289952 183134
rect 290188 182898 295882 183134
rect 296118 182898 301813 183134
rect 302049 182898 316952 183134
rect 317188 182898 322882 183134
rect 323118 182898 328813 183134
rect 329049 182898 343952 183134
rect 344188 182898 349882 183134
rect 350118 182898 355813 183134
rect 356049 182898 370952 183134
rect 371188 182898 376882 183134
rect 377118 182898 382813 183134
rect 383049 182898 397952 183134
rect 398188 182898 403882 183134
rect 404118 182898 409813 183134
rect 410049 182898 424952 183134
rect 425188 182898 430882 183134
rect 431118 182898 436813 183134
rect 437049 182898 451952 183134
rect 452188 182898 457882 183134
rect 458118 182898 463813 183134
rect 464049 182898 478952 183134
rect 479188 182898 484882 183134
rect 485118 182898 490813 183134
rect 491049 182898 505952 183134
rect 506188 182898 511882 183134
rect 512118 182898 517813 183134
rect 518049 182898 532952 183134
rect 533188 182898 538882 183134
rect 539118 182898 544813 183134
rect 545049 182898 559826 183134
rect 560062 182898 560146 183134
rect 560382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect 19794 175394 542414 175426
rect 19794 175158 19826 175394
rect 20062 175158 20146 175394
rect 20382 175158 37826 175394
rect 38062 175158 38146 175394
rect 38382 175158 55826 175394
rect 56062 175158 56146 175394
rect 56382 175158 73826 175394
rect 74062 175158 74146 175394
rect 74382 175158 91826 175394
rect 92062 175158 92146 175394
rect 92382 175158 109826 175394
rect 110062 175158 110146 175394
rect 110382 175158 127826 175394
rect 128062 175158 128146 175394
rect 128382 175158 145826 175394
rect 146062 175158 146146 175394
rect 146382 175158 163826 175394
rect 164062 175158 164146 175394
rect 164382 175158 181826 175394
rect 182062 175158 182146 175394
rect 182382 175158 199826 175394
rect 200062 175158 200146 175394
rect 200382 175158 217826 175394
rect 218062 175158 218146 175394
rect 218382 175158 235826 175394
rect 236062 175158 236146 175394
rect 236382 175158 253826 175394
rect 254062 175158 254146 175394
rect 254382 175158 271826 175394
rect 272062 175158 272146 175394
rect 272382 175158 289826 175394
rect 290062 175158 290146 175394
rect 290382 175158 307826 175394
rect 308062 175158 308146 175394
rect 308382 175158 325826 175394
rect 326062 175158 326146 175394
rect 326382 175158 343826 175394
rect 344062 175158 344146 175394
rect 344382 175158 361826 175394
rect 362062 175158 362146 175394
rect 362382 175158 379826 175394
rect 380062 175158 380146 175394
rect 380382 175158 397826 175394
rect 398062 175158 398146 175394
rect 398382 175158 415826 175394
rect 416062 175158 416146 175394
rect 416382 175158 433826 175394
rect 434062 175158 434146 175394
rect 434382 175158 451826 175394
rect 452062 175158 452146 175394
rect 452382 175158 469826 175394
rect 470062 175158 470146 175394
rect 470382 175158 487826 175394
rect 488062 175158 488146 175394
rect 488382 175158 505826 175394
rect 506062 175158 506146 175394
rect 506382 175158 523826 175394
rect 524062 175158 524146 175394
rect 524382 175158 541826 175394
rect 542062 175158 542146 175394
rect 542382 175158 542414 175394
rect 19794 175074 542414 175158
rect 19794 174838 19826 175074
rect 20062 174838 20146 175074
rect 20382 174838 37826 175074
rect 38062 174838 38146 175074
rect 38382 174838 55826 175074
rect 56062 174838 56146 175074
rect 56382 174838 73826 175074
rect 74062 174838 74146 175074
rect 74382 174838 91826 175074
rect 92062 174838 92146 175074
rect 92382 174838 109826 175074
rect 110062 174838 110146 175074
rect 110382 174838 127826 175074
rect 128062 174838 128146 175074
rect 128382 174838 145826 175074
rect 146062 174838 146146 175074
rect 146382 174838 163826 175074
rect 164062 174838 164146 175074
rect 164382 174838 181826 175074
rect 182062 174838 182146 175074
rect 182382 174838 199826 175074
rect 200062 174838 200146 175074
rect 200382 174838 217826 175074
rect 218062 174838 218146 175074
rect 218382 174838 235826 175074
rect 236062 174838 236146 175074
rect 236382 174838 253826 175074
rect 254062 174838 254146 175074
rect 254382 174838 271826 175074
rect 272062 174838 272146 175074
rect 272382 174838 289826 175074
rect 290062 174838 290146 175074
rect 290382 174838 307826 175074
rect 308062 174838 308146 175074
rect 308382 174838 325826 175074
rect 326062 174838 326146 175074
rect 326382 174838 343826 175074
rect 344062 174838 344146 175074
rect 344382 174838 361826 175074
rect 362062 174838 362146 175074
rect 362382 174838 379826 175074
rect 380062 174838 380146 175074
rect 380382 174838 397826 175074
rect 398062 174838 398146 175074
rect 398382 174838 415826 175074
rect 416062 174838 416146 175074
rect 416382 174838 433826 175074
rect 434062 174838 434146 175074
rect 434382 174838 451826 175074
rect 452062 174838 452146 175074
rect 452382 174838 469826 175074
rect 470062 174838 470146 175074
rect 470382 174838 487826 175074
rect 488062 174838 488146 175074
rect 488382 174838 505826 175074
rect 506062 174838 506146 175074
rect 506382 174838 523826 175074
rect 524062 174838 524146 175074
rect 524382 174838 541826 175074
rect 542062 174838 542146 175074
rect 542382 174838 542414 175074
rect 19794 174806 542414 174838
rect -2966 174454 586890 174486
rect -2966 174218 -2934 174454
rect -2698 174218 -2614 174454
rect -2378 174218 10826 174454
rect 11062 174218 11146 174454
rect 11382 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 46826 174454
rect 47062 174218 47146 174454
rect 47382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 82826 174454
rect 83062 174218 83146 174454
rect 83382 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 118826 174454
rect 119062 174218 119146 174454
rect 119382 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 154826 174454
rect 155062 174218 155146 174454
rect 155382 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 190826 174454
rect 191062 174218 191146 174454
rect 191382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 226826 174454
rect 227062 174218 227146 174454
rect 227382 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 262826 174454
rect 263062 174218 263146 174454
rect 263382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 298826 174454
rect 299062 174218 299146 174454
rect 299382 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 334826 174454
rect 335062 174218 335146 174454
rect 335382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 370826 174454
rect 371062 174218 371146 174454
rect 371382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 406826 174454
rect 407062 174218 407146 174454
rect 407382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 442826 174454
rect 443062 174218 443146 174454
rect 443382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 478826 174454
rect 479062 174218 479146 174454
rect 479382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 514826 174454
rect 515062 174218 515146 174454
rect 515382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 550826 174454
rect 551062 174218 551146 174454
rect 551382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 586302 174454
rect 586538 174218 586622 174454
rect 586858 174218 586890 174454
rect -2966 174134 586890 174218
rect -2966 173898 -2934 174134
rect -2698 173898 -2614 174134
rect -2378 173898 10826 174134
rect 11062 173898 11146 174134
rect 11382 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 46826 174134
rect 47062 173898 47146 174134
rect 47382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 82826 174134
rect 83062 173898 83146 174134
rect 83382 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 118826 174134
rect 119062 173898 119146 174134
rect 119382 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 154826 174134
rect 155062 173898 155146 174134
rect 155382 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 190826 174134
rect 191062 173898 191146 174134
rect 191382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 226826 174134
rect 227062 173898 227146 174134
rect 227382 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 262826 174134
rect 263062 173898 263146 174134
rect 263382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 298826 174134
rect 299062 173898 299146 174134
rect 299382 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 334826 174134
rect 335062 173898 335146 174134
rect 335382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 370826 174134
rect 371062 173898 371146 174134
rect 371382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 406826 174134
rect 407062 173898 407146 174134
rect 407382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 442826 174134
rect 443062 173898 443146 174134
rect 443382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 478826 174134
rect 479062 173898 479146 174134
rect 479382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 514826 174134
rect 515062 173898 515146 174134
rect 515382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 550826 174134
rect 551062 173898 551146 174134
rect 551382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 586302 174134
rect 586538 173898 586622 174134
rect 586858 173898 586890 174134
rect -2966 173866 586890 173898
rect -2966 165454 586890 165486
rect -2966 165218 -1974 165454
rect -1738 165218 -1654 165454
rect -1418 165218 1826 165454
rect 2062 165218 2146 165454
rect 2382 165218 19952 165454
rect 20188 165218 25882 165454
rect 26118 165218 31813 165454
rect 32049 165218 46952 165454
rect 47188 165218 52882 165454
rect 53118 165218 58813 165454
rect 59049 165218 73952 165454
rect 74188 165218 79882 165454
rect 80118 165218 85813 165454
rect 86049 165218 100952 165454
rect 101188 165218 106882 165454
rect 107118 165218 112813 165454
rect 113049 165218 127952 165454
rect 128188 165218 133882 165454
rect 134118 165218 139813 165454
rect 140049 165218 154952 165454
rect 155188 165218 160882 165454
rect 161118 165218 166813 165454
rect 167049 165218 181952 165454
rect 182188 165218 187882 165454
rect 188118 165218 193813 165454
rect 194049 165218 208952 165454
rect 209188 165218 214882 165454
rect 215118 165218 220813 165454
rect 221049 165218 235952 165454
rect 236188 165218 241882 165454
rect 242118 165218 247813 165454
rect 248049 165218 262952 165454
rect 263188 165218 268882 165454
rect 269118 165218 274813 165454
rect 275049 165218 289952 165454
rect 290188 165218 295882 165454
rect 296118 165218 301813 165454
rect 302049 165218 316952 165454
rect 317188 165218 322882 165454
rect 323118 165218 328813 165454
rect 329049 165218 343952 165454
rect 344188 165218 349882 165454
rect 350118 165218 355813 165454
rect 356049 165218 370952 165454
rect 371188 165218 376882 165454
rect 377118 165218 382813 165454
rect 383049 165218 397952 165454
rect 398188 165218 403882 165454
rect 404118 165218 409813 165454
rect 410049 165218 424952 165454
rect 425188 165218 430882 165454
rect 431118 165218 436813 165454
rect 437049 165218 451952 165454
rect 452188 165218 457882 165454
rect 458118 165218 463813 165454
rect 464049 165218 478952 165454
rect 479188 165218 484882 165454
rect 485118 165218 490813 165454
rect 491049 165218 505952 165454
rect 506188 165218 511882 165454
rect 512118 165218 517813 165454
rect 518049 165218 532952 165454
rect 533188 165218 538882 165454
rect 539118 165218 544813 165454
rect 545049 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 577826 165454
rect 578062 165218 578146 165454
rect 578382 165218 585342 165454
rect 585578 165218 585662 165454
rect 585898 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -1974 165134
rect -1738 164898 -1654 165134
rect -1418 164898 1826 165134
rect 2062 164898 2146 165134
rect 2382 164898 19952 165134
rect 20188 164898 25882 165134
rect 26118 164898 31813 165134
rect 32049 164898 46952 165134
rect 47188 164898 52882 165134
rect 53118 164898 58813 165134
rect 59049 164898 73952 165134
rect 74188 164898 79882 165134
rect 80118 164898 85813 165134
rect 86049 164898 100952 165134
rect 101188 164898 106882 165134
rect 107118 164898 112813 165134
rect 113049 164898 127952 165134
rect 128188 164898 133882 165134
rect 134118 164898 139813 165134
rect 140049 164898 154952 165134
rect 155188 164898 160882 165134
rect 161118 164898 166813 165134
rect 167049 164898 181952 165134
rect 182188 164898 187882 165134
rect 188118 164898 193813 165134
rect 194049 164898 208952 165134
rect 209188 164898 214882 165134
rect 215118 164898 220813 165134
rect 221049 164898 235952 165134
rect 236188 164898 241882 165134
rect 242118 164898 247813 165134
rect 248049 164898 262952 165134
rect 263188 164898 268882 165134
rect 269118 164898 274813 165134
rect 275049 164898 289952 165134
rect 290188 164898 295882 165134
rect 296118 164898 301813 165134
rect 302049 164898 316952 165134
rect 317188 164898 322882 165134
rect 323118 164898 328813 165134
rect 329049 164898 343952 165134
rect 344188 164898 349882 165134
rect 350118 164898 355813 165134
rect 356049 164898 370952 165134
rect 371188 164898 376882 165134
rect 377118 164898 382813 165134
rect 383049 164898 397952 165134
rect 398188 164898 403882 165134
rect 404118 164898 409813 165134
rect 410049 164898 424952 165134
rect 425188 164898 430882 165134
rect 431118 164898 436813 165134
rect 437049 164898 451952 165134
rect 452188 164898 457882 165134
rect 458118 164898 463813 165134
rect 464049 164898 478952 165134
rect 479188 164898 484882 165134
rect 485118 164898 490813 165134
rect 491049 164898 505952 165134
rect 506188 164898 511882 165134
rect 512118 164898 517813 165134
rect 518049 164898 532952 165134
rect 533188 164898 538882 165134
rect 539118 164898 544813 165134
rect 545049 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 577826 165134
rect 578062 164898 578146 165134
rect 578382 164898 585342 165134
rect 585578 164898 585662 165134
rect 585898 164898 586890 165134
rect -2966 164866 586890 164898
rect -2966 156454 586890 156486
rect -2966 156218 -2934 156454
rect -2698 156218 -2614 156454
rect -2378 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 22916 156454
rect 23152 156218 28847 156454
rect 29083 156218 49916 156454
rect 50152 156218 55847 156454
rect 56083 156218 76916 156454
rect 77152 156218 82847 156454
rect 83083 156218 103916 156454
rect 104152 156218 109847 156454
rect 110083 156218 130916 156454
rect 131152 156218 136847 156454
rect 137083 156218 157916 156454
rect 158152 156218 163847 156454
rect 164083 156218 184916 156454
rect 185152 156218 190847 156454
rect 191083 156218 211916 156454
rect 212152 156218 217847 156454
rect 218083 156218 238916 156454
rect 239152 156218 244847 156454
rect 245083 156218 265916 156454
rect 266152 156218 271847 156454
rect 272083 156218 292916 156454
rect 293152 156218 298847 156454
rect 299083 156218 319916 156454
rect 320152 156218 325847 156454
rect 326083 156218 346916 156454
rect 347152 156218 352847 156454
rect 353083 156218 373916 156454
rect 374152 156218 379847 156454
rect 380083 156218 400916 156454
rect 401152 156218 406847 156454
rect 407083 156218 427916 156454
rect 428152 156218 433847 156454
rect 434083 156218 454916 156454
rect 455152 156218 460847 156454
rect 461083 156218 481916 156454
rect 482152 156218 487847 156454
rect 488083 156218 508916 156454
rect 509152 156218 514847 156454
rect 515083 156218 535916 156454
rect 536152 156218 541847 156454
rect 542083 156218 568826 156454
rect 569062 156218 569146 156454
rect 569382 156218 586302 156454
rect 586538 156218 586622 156454
rect 586858 156218 586890 156454
rect -2966 156134 586890 156218
rect -2966 155898 -2934 156134
rect -2698 155898 -2614 156134
rect -2378 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 22916 156134
rect 23152 155898 28847 156134
rect 29083 155898 49916 156134
rect 50152 155898 55847 156134
rect 56083 155898 76916 156134
rect 77152 155898 82847 156134
rect 83083 155898 103916 156134
rect 104152 155898 109847 156134
rect 110083 155898 130916 156134
rect 131152 155898 136847 156134
rect 137083 155898 157916 156134
rect 158152 155898 163847 156134
rect 164083 155898 184916 156134
rect 185152 155898 190847 156134
rect 191083 155898 211916 156134
rect 212152 155898 217847 156134
rect 218083 155898 238916 156134
rect 239152 155898 244847 156134
rect 245083 155898 265916 156134
rect 266152 155898 271847 156134
rect 272083 155898 292916 156134
rect 293152 155898 298847 156134
rect 299083 155898 319916 156134
rect 320152 155898 325847 156134
rect 326083 155898 346916 156134
rect 347152 155898 352847 156134
rect 353083 155898 373916 156134
rect 374152 155898 379847 156134
rect 380083 155898 400916 156134
rect 401152 155898 406847 156134
rect 407083 155898 427916 156134
rect 428152 155898 433847 156134
rect 434083 155898 454916 156134
rect 455152 155898 460847 156134
rect 461083 155898 481916 156134
rect 482152 155898 487847 156134
rect 488083 155898 508916 156134
rect 509152 155898 514847 156134
rect 515083 155898 535916 156134
rect 536152 155898 541847 156134
rect 542083 155898 568826 156134
rect 569062 155898 569146 156134
rect 569382 155898 586302 156134
rect 586538 155898 586622 156134
rect 586858 155898 586890 156134
rect -2966 155866 586890 155898
rect 28794 148394 551414 148426
rect 28794 148158 28826 148394
rect 29062 148158 29146 148394
rect 29382 148158 46826 148394
rect 47062 148158 47146 148394
rect 47382 148158 64826 148394
rect 65062 148158 65146 148394
rect 65382 148158 82826 148394
rect 83062 148158 83146 148394
rect 83382 148158 100826 148394
rect 101062 148158 101146 148394
rect 101382 148158 118826 148394
rect 119062 148158 119146 148394
rect 119382 148158 136826 148394
rect 137062 148158 137146 148394
rect 137382 148158 154826 148394
rect 155062 148158 155146 148394
rect 155382 148158 172826 148394
rect 173062 148158 173146 148394
rect 173382 148158 190826 148394
rect 191062 148158 191146 148394
rect 191382 148158 208826 148394
rect 209062 148158 209146 148394
rect 209382 148158 226826 148394
rect 227062 148158 227146 148394
rect 227382 148158 244826 148394
rect 245062 148158 245146 148394
rect 245382 148158 262826 148394
rect 263062 148158 263146 148394
rect 263382 148158 280826 148394
rect 281062 148158 281146 148394
rect 281382 148158 298826 148394
rect 299062 148158 299146 148394
rect 299382 148158 316826 148394
rect 317062 148158 317146 148394
rect 317382 148158 334826 148394
rect 335062 148158 335146 148394
rect 335382 148158 352826 148394
rect 353062 148158 353146 148394
rect 353382 148158 370826 148394
rect 371062 148158 371146 148394
rect 371382 148158 388826 148394
rect 389062 148158 389146 148394
rect 389382 148158 406826 148394
rect 407062 148158 407146 148394
rect 407382 148158 424826 148394
rect 425062 148158 425146 148394
rect 425382 148158 442826 148394
rect 443062 148158 443146 148394
rect 443382 148158 460826 148394
rect 461062 148158 461146 148394
rect 461382 148158 478826 148394
rect 479062 148158 479146 148394
rect 479382 148158 496826 148394
rect 497062 148158 497146 148394
rect 497382 148158 514826 148394
rect 515062 148158 515146 148394
rect 515382 148158 532826 148394
rect 533062 148158 533146 148394
rect 533382 148158 550826 148394
rect 551062 148158 551146 148394
rect 551382 148158 551414 148394
rect 28794 148074 551414 148158
rect 28794 147838 28826 148074
rect 29062 147838 29146 148074
rect 29382 147838 46826 148074
rect 47062 147838 47146 148074
rect 47382 147838 64826 148074
rect 65062 147838 65146 148074
rect 65382 147838 82826 148074
rect 83062 147838 83146 148074
rect 83382 147838 100826 148074
rect 101062 147838 101146 148074
rect 101382 147838 118826 148074
rect 119062 147838 119146 148074
rect 119382 147838 136826 148074
rect 137062 147838 137146 148074
rect 137382 147838 154826 148074
rect 155062 147838 155146 148074
rect 155382 147838 172826 148074
rect 173062 147838 173146 148074
rect 173382 147838 190826 148074
rect 191062 147838 191146 148074
rect 191382 147838 208826 148074
rect 209062 147838 209146 148074
rect 209382 147838 226826 148074
rect 227062 147838 227146 148074
rect 227382 147838 244826 148074
rect 245062 147838 245146 148074
rect 245382 147838 262826 148074
rect 263062 147838 263146 148074
rect 263382 147838 280826 148074
rect 281062 147838 281146 148074
rect 281382 147838 298826 148074
rect 299062 147838 299146 148074
rect 299382 147838 316826 148074
rect 317062 147838 317146 148074
rect 317382 147838 334826 148074
rect 335062 147838 335146 148074
rect 335382 147838 352826 148074
rect 353062 147838 353146 148074
rect 353382 147838 370826 148074
rect 371062 147838 371146 148074
rect 371382 147838 388826 148074
rect 389062 147838 389146 148074
rect 389382 147838 406826 148074
rect 407062 147838 407146 148074
rect 407382 147838 424826 148074
rect 425062 147838 425146 148074
rect 425382 147838 442826 148074
rect 443062 147838 443146 148074
rect 443382 147838 460826 148074
rect 461062 147838 461146 148074
rect 461382 147838 478826 148074
rect 479062 147838 479146 148074
rect 479382 147838 496826 148074
rect 497062 147838 497146 148074
rect 497382 147838 514826 148074
rect 515062 147838 515146 148074
rect 515382 147838 532826 148074
rect 533062 147838 533146 148074
rect 533382 147838 550826 148074
rect 551062 147838 551146 148074
rect 551382 147838 551414 148074
rect 28794 147806 551414 147838
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 19826 147454
rect 20062 147218 20146 147454
rect 20382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 55826 147454
rect 56062 147218 56146 147454
rect 56382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 91826 147454
rect 92062 147218 92146 147454
rect 92382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 127826 147454
rect 128062 147218 128146 147454
rect 128382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 163826 147454
rect 164062 147218 164146 147454
rect 164382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 199826 147454
rect 200062 147218 200146 147454
rect 200382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 235826 147454
rect 236062 147218 236146 147454
rect 236382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 271826 147454
rect 272062 147218 272146 147454
rect 272382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 307826 147454
rect 308062 147218 308146 147454
rect 308382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 343826 147454
rect 344062 147218 344146 147454
rect 344382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 379826 147454
rect 380062 147218 380146 147454
rect 380382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 415826 147454
rect 416062 147218 416146 147454
rect 416382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 451826 147454
rect 452062 147218 452146 147454
rect 452382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 487826 147454
rect 488062 147218 488146 147454
rect 488382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 523826 147454
rect 524062 147218 524146 147454
rect 524382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 559826 147454
rect 560062 147218 560146 147454
rect 560382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 19826 147134
rect 20062 146898 20146 147134
rect 20382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 55826 147134
rect 56062 146898 56146 147134
rect 56382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 91826 147134
rect 92062 146898 92146 147134
rect 92382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 127826 147134
rect 128062 146898 128146 147134
rect 128382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 163826 147134
rect 164062 146898 164146 147134
rect 164382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 199826 147134
rect 200062 146898 200146 147134
rect 200382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 235826 147134
rect 236062 146898 236146 147134
rect 236382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 271826 147134
rect 272062 146898 272146 147134
rect 272382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 307826 147134
rect 308062 146898 308146 147134
rect 308382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 343826 147134
rect 344062 146898 344146 147134
rect 344382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 379826 147134
rect 380062 146898 380146 147134
rect 380382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 415826 147134
rect 416062 146898 416146 147134
rect 416382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 451826 147134
rect 452062 146898 452146 147134
rect 452382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 487826 147134
rect 488062 146898 488146 147134
rect 488382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 523826 147134
rect 524062 146898 524146 147134
rect 524382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 559826 147134
rect 560062 146898 560146 147134
rect 560382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -2966 138454 586890 138486
rect -2966 138218 -2934 138454
rect -2698 138218 -2614 138454
rect -2378 138218 10826 138454
rect 11062 138218 11146 138454
rect 11382 138218 22916 138454
rect 23152 138218 28847 138454
rect 29083 138218 49916 138454
rect 50152 138218 55847 138454
rect 56083 138218 76916 138454
rect 77152 138218 82847 138454
rect 83083 138218 103916 138454
rect 104152 138218 109847 138454
rect 110083 138218 130916 138454
rect 131152 138218 136847 138454
rect 137083 138218 157916 138454
rect 158152 138218 163847 138454
rect 164083 138218 184916 138454
rect 185152 138218 190847 138454
rect 191083 138218 211916 138454
rect 212152 138218 217847 138454
rect 218083 138218 238916 138454
rect 239152 138218 244847 138454
rect 245083 138218 265916 138454
rect 266152 138218 271847 138454
rect 272083 138218 292916 138454
rect 293152 138218 298847 138454
rect 299083 138218 319916 138454
rect 320152 138218 325847 138454
rect 326083 138218 346916 138454
rect 347152 138218 352847 138454
rect 353083 138218 373916 138454
rect 374152 138218 379847 138454
rect 380083 138218 400916 138454
rect 401152 138218 406847 138454
rect 407083 138218 427916 138454
rect 428152 138218 433847 138454
rect 434083 138218 454916 138454
rect 455152 138218 460847 138454
rect 461083 138218 481916 138454
rect 482152 138218 487847 138454
rect 488083 138218 508916 138454
rect 509152 138218 514847 138454
rect 515083 138218 535916 138454
rect 536152 138218 541847 138454
rect 542083 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 586302 138454
rect 586538 138218 586622 138454
rect 586858 138218 586890 138454
rect -2966 138134 586890 138218
rect -2966 137898 -2934 138134
rect -2698 137898 -2614 138134
rect -2378 137898 10826 138134
rect 11062 137898 11146 138134
rect 11382 137898 22916 138134
rect 23152 137898 28847 138134
rect 29083 137898 49916 138134
rect 50152 137898 55847 138134
rect 56083 137898 76916 138134
rect 77152 137898 82847 138134
rect 83083 137898 103916 138134
rect 104152 137898 109847 138134
rect 110083 137898 130916 138134
rect 131152 137898 136847 138134
rect 137083 137898 157916 138134
rect 158152 137898 163847 138134
rect 164083 137898 184916 138134
rect 185152 137898 190847 138134
rect 191083 137898 211916 138134
rect 212152 137898 217847 138134
rect 218083 137898 238916 138134
rect 239152 137898 244847 138134
rect 245083 137898 265916 138134
rect 266152 137898 271847 138134
rect 272083 137898 292916 138134
rect 293152 137898 298847 138134
rect 299083 137898 319916 138134
rect 320152 137898 325847 138134
rect 326083 137898 346916 138134
rect 347152 137898 352847 138134
rect 353083 137898 373916 138134
rect 374152 137898 379847 138134
rect 380083 137898 400916 138134
rect 401152 137898 406847 138134
rect 407083 137898 427916 138134
rect 428152 137898 433847 138134
rect 434083 137898 454916 138134
rect 455152 137898 460847 138134
rect 461083 137898 481916 138134
rect 482152 137898 487847 138134
rect 488083 137898 508916 138134
rect 509152 137898 514847 138134
rect 515083 137898 535916 138134
rect 536152 137898 541847 138134
rect 542083 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 586302 138134
rect 586538 137898 586622 138134
rect 586858 137898 586890 138134
rect -2966 137866 586890 137898
rect -2966 129454 586890 129486
rect -2966 129218 -1974 129454
rect -1738 129218 -1654 129454
rect -1418 129218 1826 129454
rect 2062 129218 2146 129454
rect 2382 129218 19952 129454
rect 20188 129218 25882 129454
rect 26118 129218 31813 129454
rect 32049 129218 46952 129454
rect 47188 129218 52882 129454
rect 53118 129218 58813 129454
rect 59049 129218 73952 129454
rect 74188 129218 79882 129454
rect 80118 129218 85813 129454
rect 86049 129218 100952 129454
rect 101188 129218 106882 129454
rect 107118 129218 112813 129454
rect 113049 129218 127952 129454
rect 128188 129218 133882 129454
rect 134118 129218 139813 129454
rect 140049 129218 154952 129454
rect 155188 129218 160882 129454
rect 161118 129218 166813 129454
rect 167049 129218 181952 129454
rect 182188 129218 187882 129454
rect 188118 129218 193813 129454
rect 194049 129218 208952 129454
rect 209188 129218 214882 129454
rect 215118 129218 220813 129454
rect 221049 129218 235952 129454
rect 236188 129218 241882 129454
rect 242118 129218 247813 129454
rect 248049 129218 262952 129454
rect 263188 129218 268882 129454
rect 269118 129218 274813 129454
rect 275049 129218 289952 129454
rect 290188 129218 295882 129454
rect 296118 129218 301813 129454
rect 302049 129218 316952 129454
rect 317188 129218 322882 129454
rect 323118 129218 328813 129454
rect 329049 129218 343952 129454
rect 344188 129218 349882 129454
rect 350118 129218 355813 129454
rect 356049 129218 370952 129454
rect 371188 129218 376882 129454
rect 377118 129218 382813 129454
rect 383049 129218 397952 129454
rect 398188 129218 403882 129454
rect 404118 129218 409813 129454
rect 410049 129218 424952 129454
rect 425188 129218 430882 129454
rect 431118 129218 436813 129454
rect 437049 129218 451952 129454
rect 452188 129218 457882 129454
rect 458118 129218 463813 129454
rect 464049 129218 478952 129454
rect 479188 129218 484882 129454
rect 485118 129218 490813 129454
rect 491049 129218 505952 129454
rect 506188 129218 511882 129454
rect 512118 129218 517813 129454
rect 518049 129218 532952 129454
rect 533188 129218 538882 129454
rect 539118 129218 544813 129454
rect 545049 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 577826 129454
rect 578062 129218 578146 129454
rect 578382 129218 585342 129454
rect 585578 129218 585662 129454
rect 585898 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -1974 129134
rect -1738 128898 -1654 129134
rect -1418 128898 1826 129134
rect 2062 128898 2146 129134
rect 2382 128898 19952 129134
rect 20188 128898 25882 129134
rect 26118 128898 31813 129134
rect 32049 128898 46952 129134
rect 47188 128898 52882 129134
rect 53118 128898 58813 129134
rect 59049 128898 73952 129134
rect 74188 128898 79882 129134
rect 80118 128898 85813 129134
rect 86049 128898 100952 129134
rect 101188 128898 106882 129134
rect 107118 128898 112813 129134
rect 113049 128898 127952 129134
rect 128188 128898 133882 129134
rect 134118 128898 139813 129134
rect 140049 128898 154952 129134
rect 155188 128898 160882 129134
rect 161118 128898 166813 129134
rect 167049 128898 181952 129134
rect 182188 128898 187882 129134
rect 188118 128898 193813 129134
rect 194049 128898 208952 129134
rect 209188 128898 214882 129134
rect 215118 128898 220813 129134
rect 221049 128898 235952 129134
rect 236188 128898 241882 129134
rect 242118 128898 247813 129134
rect 248049 128898 262952 129134
rect 263188 128898 268882 129134
rect 269118 128898 274813 129134
rect 275049 128898 289952 129134
rect 290188 128898 295882 129134
rect 296118 128898 301813 129134
rect 302049 128898 316952 129134
rect 317188 128898 322882 129134
rect 323118 128898 328813 129134
rect 329049 128898 343952 129134
rect 344188 128898 349882 129134
rect 350118 128898 355813 129134
rect 356049 128898 370952 129134
rect 371188 128898 376882 129134
rect 377118 128898 382813 129134
rect 383049 128898 397952 129134
rect 398188 128898 403882 129134
rect 404118 128898 409813 129134
rect 410049 128898 424952 129134
rect 425188 128898 430882 129134
rect 431118 128898 436813 129134
rect 437049 128898 451952 129134
rect 452188 128898 457882 129134
rect 458118 128898 463813 129134
rect 464049 128898 478952 129134
rect 479188 128898 484882 129134
rect 485118 128898 490813 129134
rect 491049 128898 505952 129134
rect 506188 128898 511882 129134
rect 512118 128898 517813 129134
rect 518049 128898 532952 129134
rect 533188 128898 538882 129134
rect 539118 128898 544813 129134
rect 545049 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 577826 129134
rect 578062 128898 578146 129134
rect 578382 128898 585342 129134
rect 585578 128898 585662 129134
rect 585898 128898 586890 129134
rect -2966 128866 586890 128898
rect 19794 121394 542414 121426
rect 19794 121158 19826 121394
rect 20062 121158 20146 121394
rect 20382 121158 37826 121394
rect 38062 121158 38146 121394
rect 38382 121158 55826 121394
rect 56062 121158 56146 121394
rect 56382 121158 73826 121394
rect 74062 121158 74146 121394
rect 74382 121158 91826 121394
rect 92062 121158 92146 121394
rect 92382 121158 109826 121394
rect 110062 121158 110146 121394
rect 110382 121158 127826 121394
rect 128062 121158 128146 121394
rect 128382 121158 145826 121394
rect 146062 121158 146146 121394
rect 146382 121158 163826 121394
rect 164062 121158 164146 121394
rect 164382 121158 181826 121394
rect 182062 121158 182146 121394
rect 182382 121158 199826 121394
rect 200062 121158 200146 121394
rect 200382 121158 217826 121394
rect 218062 121158 218146 121394
rect 218382 121158 235826 121394
rect 236062 121158 236146 121394
rect 236382 121158 253826 121394
rect 254062 121158 254146 121394
rect 254382 121158 271826 121394
rect 272062 121158 272146 121394
rect 272382 121158 289826 121394
rect 290062 121158 290146 121394
rect 290382 121158 307826 121394
rect 308062 121158 308146 121394
rect 308382 121158 325826 121394
rect 326062 121158 326146 121394
rect 326382 121158 343826 121394
rect 344062 121158 344146 121394
rect 344382 121158 361826 121394
rect 362062 121158 362146 121394
rect 362382 121158 379826 121394
rect 380062 121158 380146 121394
rect 380382 121158 397826 121394
rect 398062 121158 398146 121394
rect 398382 121158 415826 121394
rect 416062 121158 416146 121394
rect 416382 121158 433826 121394
rect 434062 121158 434146 121394
rect 434382 121158 451826 121394
rect 452062 121158 452146 121394
rect 452382 121158 469826 121394
rect 470062 121158 470146 121394
rect 470382 121158 487826 121394
rect 488062 121158 488146 121394
rect 488382 121158 505826 121394
rect 506062 121158 506146 121394
rect 506382 121158 523826 121394
rect 524062 121158 524146 121394
rect 524382 121158 541826 121394
rect 542062 121158 542146 121394
rect 542382 121158 542414 121394
rect 19794 121074 542414 121158
rect 19794 120838 19826 121074
rect 20062 120838 20146 121074
rect 20382 120838 37826 121074
rect 38062 120838 38146 121074
rect 38382 120838 55826 121074
rect 56062 120838 56146 121074
rect 56382 120838 73826 121074
rect 74062 120838 74146 121074
rect 74382 120838 91826 121074
rect 92062 120838 92146 121074
rect 92382 120838 109826 121074
rect 110062 120838 110146 121074
rect 110382 120838 127826 121074
rect 128062 120838 128146 121074
rect 128382 120838 145826 121074
rect 146062 120838 146146 121074
rect 146382 120838 163826 121074
rect 164062 120838 164146 121074
rect 164382 120838 181826 121074
rect 182062 120838 182146 121074
rect 182382 120838 199826 121074
rect 200062 120838 200146 121074
rect 200382 120838 217826 121074
rect 218062 120838 218146 121074
rect 218382 120838 235826 121074
rect 236062 120838 236146 121074
rect 236382 120838 253826 121074
rect 254062 120838 254146 121074
rect 254382 120838 271826 121074
rect 272062 120838 272146 121074
rect 272382 120838 289826 121074
rect 290062 120838 290146 121074
rect 290382 120838 307826 121074
rect 308062 120838 308146 121074
rect 308382 120838 325826 121074
rect 326062 120838 326146 121074
rect 326382 120838 343826 121074
rect 344062 120838 344146 121074
rect 344382 120838 361826 121074
rect 362062 120838 362146 121074
rect 362382 120838 379826 121074
rect 380062 120838 380146 121074
rect 380382 120838 397826 121074
rect 398062 120838 398146 121074
rect 398382 120838 415826 121074
rect 416062 120838 416146 121074
rect 416382 120838 433826 121074
rect 434062 120838 434146 121074
rect 434382 120838 451826 121074
rect 452062 120838 452146 121074
rect 452382 120838 469826 121074
rect 470062 120838 470146 121074
rect 470382 120838 487826 121074
rect 488062 120838 488146 121074
rect 488382 120838 505826 121074
rect 506062 120838 506146 121074
rect 506382 120838 523826 121074
rect 524062 120838 524146 121074
rect 524382 120838 541826 121074
rect 542062 120838 542146 121074
rect 542382 120838 542414 121074
rect 19794 120806 542414 120838
rect -2966 120454 586890 120486
rect -2966 120218 -2934 120454
rect -2698 120218 -2614 120454
rect -2378 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 28826 120454
rect 29062 120218 29146 120454
rect 29382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 64826 120454
rect 65062 120218 65146 120454
rect 65382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 100826 120454
rect 101062 120218 101146 120454
rect 101382 120218 118826 120454
rect 119062 120218 119146 120454
rect 119382 120218 136826 120454
rect 137062 120218 137146 120454
rect 137382 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 172826 120454
rect 173062 120218 173146 120454
rect 173382 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 208826 120454
rect 209062 120218 209146 120454
rect 209382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 244826 120454
rect 245062 120218 245146 120454
rect 245382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 280826 120454
rect 281062 120218 281146 120454
rect 281382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 316826 120454
rect 317062 120218 317146 120454
rect 317382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 352826 120454
rect 353062 120218 353146 120454
rect 353382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 388826 120454
rect 389062 120218 389146 120454
rect 389382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 424826 120454
rect 425062 120218 425146 120454
rect 425382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 460826 120454
rect 461062 120218 461146 120454
rect 461382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 496826 120454
rect 497062 120218 497146 120454
rect 497382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 532826 120454
rect 533062 120218 533146 120454
rect 533382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 568826 120454
rect 569062 120218 569146 120454
rect 569382 120218 586302 120454
rect 586538 120218 586622 120454
rect 586858 120218 586890 120454
rect -2966 120134 586890 120218
rect -2966 119898 -2934 120134
rect -2698 119898 -2614 120134
rect -2378 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 28826 120134
rect 29062 119898 29146 120134
rect 29382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 64826 120134
rect 65062 119898 65146 120134
rect 65382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 100826 120134
rect 101062 119898 101146 120134
rect 101382 119898 118826 120134
rect 119062 119898 119146 120134
rect 119382 119898 136826 120134
rect 137062 119898 137146 120134
rect 137382 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 172826 120134
rect 173062 119898 173146 120134
rect 173382 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 208826 120134
rect 209062 119898 209146 120134
rect 209382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 244826 120134
rect 245062 119898 245146 120134
rect 245382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 280826 120134
rect 281062 119898 281146 120134
rect 281382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 316826 120134
rect 317062 119898 317146 120134
rect 317382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 352826 120134
rect 353062 119898 353146 120134
rect 353382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 388826 120134
rect 389062 119898 389146 120134
rect 389382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 424826 120134
rect 425062 119898 425146 120134
rect 425382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 460826 120134
rect 461062 119898 461146 120134
rect 461382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 496826 120134
rect 497062 119898 497146 120134
rect 497382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 532826 120134
rect 533062 119898 533146 120134
rect 533382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 568826 120134
rect 569062 119898 569146 120134
rect 569382 119898 586302 120134
rect 586538 119898 586622 120134
rect 586858 119898 586890 120134
rect -2966 119866 586890 119898
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 19952 111454
rect 20188 111218 25882 111454
rect 26118 111218 31813 111454
rect 32049 111218 46952 111454
rect 47188 111218 52882 111454
rect 53118 111218 58813 111454
rect 59049 111218 73952 111454
rect 74188 111218 79882 111454
rect 80118 111218 85813 111454
rect 86049 111218 100952 111454
rect 101188 111218 106882 111454
rect 107118 111218 112813 111454
rect 113049 111218 127952 111454
rect 128188 111218 133882 111454
rect 134118 111218 139813 111454
rect 140049 111218 154952 111454
rect 155188 111218 160882 111454
rect 161118 111218 166813 111454
rect 167049 111218 181952 111454
rect 182188 111218 187882 111454
rect 188118 111218 193813 111454
rect 194049 111218 208952 111454
rect 209188 111218 214882 111454
rect 215118 111218 220813 111454
rect 221049 111218 235952 111454
rect 236188 111218 241882 111454
rect 242118 111218 247813 111454
rect 248049 111218 262952 111454
rect 263188 111218 268882 111454
rect 269118 111218 274813 111454
rect 275049 111218 289952 111454
rect 290188 111218 295882 111454
rect 296118 111218 301813 111454
rect 302049 111218 316952 111454
rect 317188 111218 322882 111454
rect 323118 111218 328813 111454
rect 329049 111218 343952 111454
rect 344188 111218 349882 111454
rect 350118 111218 355813 111454
rect 356049 111218 370952 111454
rect 371188 111218 376882 111454
rect 377118 111218 382813 111454
rect 383049 111218 397952 111454
rect 398188 111218 403882 111454
rect 404118 111218 409813 111454
rect 410049 111218 424952 111454
rect 425188 111218 430882 111454
rect 431118 111218 436813 111454
rect 437049 111218 451952 111454
rect 452188 111218 457882 111454
rect 458118 111218 463813 111454
rect 464049 111218 478952 111454
rect 479188 111218 484882 111454
rect 485118 111218 490813 111454
rect 491049 111218 505952 111454
rect 506188 111218 511882 111454
rect 512118 111218 517813 111454
rect 518049 111218 532952 111454
rect 533188 111218 538882 111454
rect 539118 111218 544813 111454
rect 545049 111218 559826 111454
rect 560062 111218 560146 111454
rect 560382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 19952 111134
rect 20188 110898 25882 111134
rect 26118 110898 31813 111134
rect 32049 110898 46952 111134
rect 47188 110898 52882 111134
rect 53118 110898 58813 111134
rect 59049 110898 73952 111134
rect 74188 110898 79882 111134
rect 80118 110898 85813 111134
rect 86049 110898 100952 111134
rect 101188 110898 106882 111134
rect 107118 110898 112813 111134
rect 113049 110898 127952 111134
rect 128188 110898 133882 111134
rect 134118 110898 139813 111134
rect 140049 110898 154952 111134
rect 155188 110898 160882 111134
rect 161118 110898 166813 111134
rect 167049 110898 181952 111134
rect 182188 110898 187882 111134
rect 188118 110898 193813 111134
rect 194049 110898 208952 111134
rect 209188 110898 214882 111134
rect 215118 110898 220813 111134
rect 221049 110898 235952 111134
rect 236188 110898 241882 111134
rect 242118 110898 247813 111134
rect 248049 110898 262952 111134
rect 263188 110898 268882 111134
rect 269118 110898 274813 111134
rect 275049 110898 289952 111134
rect 290188 110898 295882 111134
rect 296118 110898 301813 111134
rect 302049 110898 316952 111134
rect 317188 110898 322882 111134
rect 323118 110898 328813 111134
rect 329049 110898 343952 111134
rect 344188 110898 349882 111134
rect 350118 110898 355813 111134
rect 356049 110898 370952 111134
rect 371188 110898 376882 111134
rect 377118 110898 382813 111134
rect 383049 110898 397952 111134
rect 398188 110898 403882 111134
rect 404118 110898 409813 111134
rect 410049 110898 424952 111134
rect 425188 110898 430882 111134
rect 431118 110898 436813 111134
rect 437049 110898 451952 111134
rect 452188 110898 457882 111134
rect 458118 110898 463813 111134
rect 464049 110898 478952 111134
rect 479188 110898 484882 111134
rect 485118 110898 490813 111134
rect 491049 110898 505952 111134
rect 506188 110898 511882 111134
rect 512118 110898 517813 111134
rect 518049 110898 532952 111134
rect 533188 110898 538882 111134
rect 539118 110898 544813 111134
rect 545049 110898 559826 111134
rect 560062 110898 560146 111134
rect 560382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -2966 102454 586890 102486
rect -2966 102218 -2934 102454
rect -2698 102218 -2614 102454
rect -2378 102218 10826 102454
rect 11062 102218 11146 102454
rect 11382 102218 22916 102454
rect 23152 102218 28847 102454
rect 29083 102218 49916 102454
rect 50152 102218 55847 102454
rect 56083 102218 76916 102454
rect 77152 102218 82847 102454
rect 83083 102218 103916 102454
rect 104152 102218 109847 102454
rect 110083 102218 130916 102454
rect 131152 102218 136847 102454
rect 137083 102218 157916 102454
rect 158152 102218 163847 102454
rect 164083 102218 184916 102454
rect 185152 102218 190847 102454
rect 191083 102218 211916 102454
rect 212152 102218 217847 102454
rect 218083 102218 238916 102454
rect 239152 102218 244847 102454
rect 245083 102218 265916 102454
rect 266152 102218 271847 102454
rect 272083 102218 292916 102454
rect 293152 102218 298847 102454
rect 299083 102218 319916 102454
rect 320152 102218 325847 102454
rect 326083 102218 346916 102454
rect 347152 102218 352847 102454
rect 353083 102218 373916 102454
rect 374152 102218 379847 102454
rect 380083 102218 400916 102454
rect 401152 102218 406847 102454
rect 407083 102218 427916 102454
rect 428152 102218 433847 102454
rect 434083 102218 454916 102454
rect 455152 102218 460847 102454
rect 461083 102218 481916 102454
rect 482152 102218 487847 102454
rect 488083 102218 508916 102454
rect 509152 102218 514847 102454
rect 515083 102218 535916 102454
rect 536152 102218 541847 102454
rect 542083 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 586302 102454
rect 586538 102218 586622 102454
rect 586858 102218 586890 102454
rect -2966 102134 586890 102218
rect -2966 101898 -2934 102134
rect -2698 101898 -2614 102134
rect -2378 101898 10826 102134
rect 11062 101898 11146 102134
rect 11382 101898 22916 102134
rect 23152 101898 28847 102134
rect 29083 101898 49916 102134
rect 50152 101898 55847 102134
rect 56083 101898 76916 102134
rect 77152 101898 82847 102134
rect 83083 101898 103916 102134
rect 104152 101898 109847 102134
rect 110083 101898 130916 102134
rect 131152 101898 136847 102134
rect 137083 101898 157916 102134
rect 158152 101898 163847 102134
rect 164083 101898 184916 102134
rect 185152 101898 190847 102134
rect 191083 101898 211916 102134
rect 212152 101898 217847 102134
rect 218083 101898 238916 102134
rect 239152 101898 244847 102134
rect 245083 101898 265916 102134
rect 266152 101898 271847 102134
rect 272083 101898 292916 102134
rect 293152 101898 298847 102134
rect 299083 101898 319916 102134
rect 320152 101898 325847 102134
rect 326083 101898 346916 102134
rect 347152 101898 352847 102134
rect 353083 101898 373916 102134
rect 374152 101898 379847 102134
rect 380083 101898 400916 102134
rect 401152 101898 406847 102134
rect 407083 101898 427916 102134
rect 428152 101898 433847 102134
rect 434083 101898 454916 102134
rect 455152 101898 460847 102134
rect 461083 101898 481916 102134
rect 482152 101898 487847 102134
rect 488083 101898 508916 102134
rect 509152 101898 514847 102134
rect 515083 101898 535916 102134
rect 536152 101898 541847 102134
rect 542083 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 586302 102134
rect 586538 101898 586622 102134
rect 586858 101898 586890 102134
rect -2966 101866 586890 101898
rect 28794 94394 551414 94426
rect 28794 94158 28826 94394
rect 29062 94158 29146 94394
rect 29382 94158 46826 94394
rect 47062 94158 47146 94394
rect 47382 94158 64826 94394
rect 65062 94158 65146 94394
rect 65382 94158 82826 94394
rect 83062 94158 83146 94394
rect 83382 94158 100826 94394
rect 101062 94158 101146 94394
rect 101382 94158 118826 94394
rect 119062 94158 119146 94394
rect 119382 94158 136826 94394
rect 137062 94158 137146 94394
rect 137382 94158 154826 94394
rect 155062 94158 155146 94394
rect 155382 94158 172826 94394
rect 173062 94158 173146 94394
rect 173382 94158 190826 94394
rect 191062 94158 191146 94394
rect 191382 94158 208826 94394
rect 209062 94158 209146 94394
rect 209382 94158 226826 94394
rect 227062 94158 227146 94394
rect 227382 94158 244826 94394
rect 245062 94158 245146 94394
rect 245382 94158 262826 94394
rect 263062 94158 263146 94394
rect 263382 94158 280826 94394
rect 281062 94158 281146 94394
rect 281382 94158 298826 94394
rect 299062 94158 299146 94394
rect 299382 94158 316826 94394
rect 317062 94158 317146 94394
rect 317382 94158 334826 94394
rect 335062 94158 335146 94394
rect 335382 94158 352826 94394
rect 353062 94158 353146 94394
rect 353382 94158 370826 94394
rect 371062 94158 371146 94394
rect 371382 94158 388826 94394
rect 389062 94158 389146 94394
rect 389382 94158 406826 94394
rect 407062 94158 407146 94394
rect 407382 94158 424826 94394
rect 425062 94158 425146 94394
rect 425382 94158 442826 94394
rect 443062 94158 443146 94394
rect 443382 94158 460826 94394
rect 461062 94158 461146 94394
rect 461382 94158 478826 94394
rect 479062 94158 479146 94394
rect 479382 94158 496826 94394
rect 497062 94158 497146 94394
rect 497382 94158 514826 94394
rect 515062 94158 515146 94394
rect 515382 94158 532826 94394
rect 533062 94158 533146 94394
rect 533382 94158 550826 94394
rect 551062 94158 551146 94394
rect 551382 94158 551414 94394
rect 28794 94074 551414 94158
rect 28794 93838 28826 94074
rect 29062 93838 29146 94074
rect 29382 93838 46826 94074
rect 47062 93838 47146 94074
rect 47382 93838 64826 94074
rect 65062 93838 65146 94074
rect 65382 93838 82826 94074
rect 83062 93838 83146 94074
rect 83382 93838 100826 94074
rect 101062 93838 101146 94074
rect 101382 93838 118826 94074
rect 119062 93838 119146 94074
rect 119382 93838 136826 94074
rect 137062 93838 137146 94074
rect 137382 93838 154826 94074
rect 155062 93838 155146 94074
rect 155382 93838 172826 94074
rect 173062 93838 173146 94074
rect 173382 93838 190826 94074
rect 191062 93838 191146 94074
rect 191382 93838 208826 94074
rect 209062 93838 209146 94074
rect 209382 93838 226826 94074
rect 227062 93838 227146 94074
rect 227382 93838 244826 94074
rect 245062 93838 245146 94074
rect 245382 93838 262826 94074
rect 263062 93838 263146 94074
rect 263382 93838 280826 94074
rect 281062 93838 281146 94074
rect 281382 93838 298826 94074
rect 299062 93838 299146 94074
rect 299382 93838 316826 94074
rect 317062 93838 317146 94074
rect 317382 93838 334826 94074
rect 335062 93838 335146 94074
rect 335382 93838 352826 94074
rect 353062 93838 353146 94074
rect 353382 93838 370826 94074
rect 371062 93838 371146 94074
rect 371382 93838 388826 94074
rect 389062 93838 389146 94074
rect 389382 93838 406826 94074
rect 407062 93838 407146 94074
rect 407382 93838 424826 94074
rect 425062 93838 425146 94074
rect 425382 93838 442826 94074
rect 443062 93838 443146 94074
rect 443382 93838 460826 94074
rect 461062 93838 461146 94074
rect 461382 93838 478826 94074
rect 479062 93838 479146 94074
rect 479382 93838 496826 94074
rect 497062 93838 497146 94074
rect 497382 93838 514826 94074
rect 515062 93838 515146 94074
rect 515382 93838 532826 94074
rect 533062 93838 533146 94074
rect 533382 93838 550826 94074
rect 551062 93838 551146 94074
rect 551382 93838 551414 94074
rect 28794 93806 551414 93838
rect -2966 93454 586890 93486
rect -2966 93218 -1974 93454
rect -1738 93218 -1654 93454
rect -1418 93218 1826 93454
rect 2062 93218 2146 93454
rect 2382 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 37826 93454
rect 38062 93218 38146 93454
rect 38382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 73826 93454
rect 74062 93218 74146 93454
rect 74382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 109826 93454
rect 110062 93218 110146 93454
rect 110382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 145826 93454
rect 146062 93218 146146 93454
rect 146382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 181826 93454
rect 182062 93218 182146 93454
rect 182382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 217826 93454
rect 218062 93218 218146 93454
rect 218382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 253826 93454
rect 254062 93218 254146 93454
rect 254382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 289826 93454
rect 290062 93218 290146 93454
rect 290382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 325826 93454
rect 326062 93218 326146 93454
rect 326382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 361826 93454
rect 362062 93218 362146 93454
rect 362382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 397826 93454
rect 398062 93218 398146 93454
rect 398382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 433826 93454
rect 434062 93218 434146 93454
rect 434382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 469826 93454
rect 470062 93218 470146 93454
rect 470382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 505826 93454
rect 506062 93218 506146 93454
rect 506382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 541826 93454
rect 542062 93218 542146 93454
rect 542382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 577826 93454
rect 578062 93218 578146 93454
rect 578382 93218 585342 93454
rect 585578 93218 585662 93454
rect 585898 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -1974 93134
rect -1738 92898 -1654 93134
rect -1418 92898 1826 93134
rect 2062 92898 2146 93134
rect 2382 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 37826 93134
rect 38062 92898 38146 93134
rect 38382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 73826 93134
rect 74062 92898 74146 93134
rect 74382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 109826 93134
rect 110062 92898 110146 93134
rect 110382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 145826 93134
rect 146062 92898 146146 93134
rect 146382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 181826 93134
rect 182062 92898 182146 93134
rect 182382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 217826 93134
rect 218062 92898 218146 93134
rect 218382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 253826 93134
rect 254062 92898 254146 93134
rect 254382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 289826 93134
rect 290062 92898 290146 93134
rect 290382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 325826 93134
rect 326062 92898 326146 93134
rect 326382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 361826 93134
rect 362062 92898 362146 93134
rect 362382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 397826 93134
rect 398062 92898 398146 93134
rect 398382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 433826 93134
rect 434062 92898 434146 93134
rect 434382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 469826 93134
rect 470062 92898 470146 93134
rect 470382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 505826 93134
rect 506062 92898 506146 93134
rect 506382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 541826 93134
rect 542062 92898 542146 93134
rect 542382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 577826 93134
rect 578062 92898 578146 93134
rect 578382 92898 585342 93134
rect 585578 92898 585662 93134
rect 585898 92898 586890 93134
rect -2966 92866 586890 92898
rect -2966 84454 586890 84486
rect -2966 84218 -2934 84454
rect -2698 84218 -2614 84454
rect -2378 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 22916 84454
rect 23152 84218 28847 84454
rect 29083 84218 49916 84454
rect 50152 84218 55847 84454
rect 56083 84218 76916 84454
rect 77152 84218 82847 84454
rect 83083 84218 103916 84454
rect 104152 84218 109847 84454
rect 110083 84218 130916 84454
rect 131152 84218 136847 84454
rect 137083 84218 157916 84454
rect 158152 84218 163847 84454
rect 164083 84218 184916 84454
rect 185152 84218 190847 84454
rect 191083 84218 211916 84454
rect 212152 84218 217847 84454
rect 218083 84218 238916 84454
rect 239152 84218 244847 84454
rect 245083 84218 265916 84454
rect 266152 84218 271847 84454
rect 272083 84218 292916 84454
rect 293152 84218 298847 84454
rect 299083 84218 319916 84454
rect 320152 84218 325847 84454
rect 326083 84218 346916 84454
rect 347152 84218 352847 84454
rect 353083 84218 373916 84454
rect 374152 84218 379847 84454
rect 380083 84218 400916 84454
rect 401152 84218 406847 84454
rect 407083 84218 427916 84454
rect 428152 84218 433847 84454
rect 434083 84218 454916 84454
rect 455152 84218 460847 84454
rect 461083 84218 481916 84454
rect 482152 84218 487847 84454
rect 488083 84218 508916 84454
rect 509152 84218 514847 84454
rect 515083 84218 535916 84454
rect 536152 84218 541847 84454
rect 542083 84218 568826 84454
rect 569062 84218 569146 84454
rect 569382 84218 586302 84454
rect 586538 84218 586622 84454
rect 586858 84218 586890 84454
rect -2966 84134 586890 84218
rect -2966 83898 -2934 84134
rect -2698 83898 -2614 84134
rect -2378 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 22916 84134
rect 23152 83898 28847 84134
rect 29083 83898 49916 84134
rect 50152 83898 55847 84134
rect 56083 83898 76916 84134
rect 77152 83898 82847 84134
rect 83083 83898 103916 84134
rect 104152 83898 109847 84134
rect 110083 83898 130916 84134
rect 131152 83898 136847 84134
rect 137083 83898 157916 84134
rect 158152 83898 163847 84134
rect 164083 83898 184916 84134
rect 185152 83898 190847 84134
rect 191083 83898 211916 84134
rect 212152 83898 217847 84134
rect 218083 83898 238916 84134
rect 239152 83898 244847 84134
rect 245083 83898 265916 84134
rect 266152 83898 271847 84134
rect 272083 83898 292916 84134
rect 293152 83898 298847 84134
rect 299083 83898 319916 84134
rect 320152 83898 325847 84134
rect 326083 83898 346916 84134
rect 347152 83898 352847 84134
rect 353083 83898 373916 84134
rect 374152 83898 379847 84134
rect 380083 83898 400916 84134
rect 401152 83898 406847 84134
rect 407083 83898 427916 84134
rect 428152 83898 433847 84134
rect 434083 83898 454916 84134
rect 455152 83898 460847 84134
rect 461083 83898 481916 84134
rect 482152 83898 487847 84134
rect 488083 83898 508916 84134
rect 509152 83898 514847 84134
rect 515083 83898 535916 84134
rect 536152 83898 541847 84134
rect 542083 83898 568826 84134
rect 569062 83898 569146 84134
rect 569382 83898 586302 84134
rect 586538 83898 586622 84134
rect 586858 83898 586890 84134
rect -2966 83866 586890 83898
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 19952 75454
rect 20188 75218 25882 75454
rect 26118 75218 31813 75454
rect 32049 75218 46952 75454
rect 47188 75218 52882 75454
rect 53118 75218 58813 75454
rect 59049 75218 73952 75454
rect 74188 75218 79882 75454
rect 80118 75218 85813 75454
rect 86049 75218 100952 75454
rect 101188 75218 106882 75454
rect 107118 75218 112813 75454
rect 113049 75218 127952 75454
rect 128188 75218 133882 75454
rect 134118 75218 139813 75454
rect 140049 75218 154952 75454
rect 155188 75218 160882 75454
rect 161118 75218 166813 75454
rect 167049 75218 181952 75454
rect 182188 75218 187882 75454
rect 188118 75218 193813 75454
rect 194049 75218 208952 75454
rect 209188 75218 214882 75454
rect 215118 75218 220813 75454
rect 221049 75218 235952 75454
rect 236188 75218 241882 75454
rect 242118 75218 247813 75454
rect 248049 75218 262952 75454
rect 263188 75218 268882 75454
rect 269118 75218 274813 75454
rect 275049 75218 289952 75454
rect 290188 75218 295882 75454
rect 296118 75218 301813 75454
rect 302049 75218 316952 75454
rect 317188 75218 322882 75454
rect 323118 75218 328813 75454
rect 329049 75218 343952 75454
rect 344188 75218 349882 75454
rect 350118 75218 355813 75454
rect 356049 75218 370952 75454
rect 371188 75218 376882 75454
rect 377118 75218 382813 75454
rect 383049 75218 397952 75454
rect 398188 75218 403882 75454
rect 404118 75218 409813 75454
rect 410049 75218 424952 75454
rect 425188 75218 430882 75454
rect 431118 75218 436813 75454
rect 437049 75218 451952 75454
rect 452188 75218 457882 75454
rect 458118 75218 463813 75454
rect 464049 75218 478952 75454
rect 479188 75218 484882 75454
rect 485118 75218 490813 75454
rect 491049 75218 505952 75454
rect 506188 75218 511882 75454
rect 512118 75218 517813 75454
rect 518049 75218 532952 75454
rect 533188 75218 538882 75454
rect 539118 75218 544813 75454
rect 545049 75218 559826 75454
rect 560062 75218 560146 75454
rect 560382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 19952 75134
rect 20188 74898 25882 75134
rect 26118 74898 31813 75134
rect 32049 74898 46952 75134
rect 47188 74898 52882 75134
rect 53118 74898 58813 75134
rect 59049 74898 73952 75134
rect 74188 74898 79882 75134
rect 80118 74898 85813 75134
rect 86049 74898 100952 75134
rect 101188 74898 106882 75134
rect 107118 74898 112813 75134
rect 113049 74898 127952 75134
rect 128188 74898 133882 75134
rect 134118 74898 139813 75134
rect 140049 74898 154952 75134
rect 155188 74898 160882 75134
rect 161118 74898 166813 75134
rect 167049 74898 181952 75134
rect 182188 74898 187882 75134
rect 188118 74898 193813 75134
rect 194049 74898 208952 75134
rect 209188 74898 214882 75134
rect 215118 74898 220813 75134
rect 221049 74898 235952 75134
rect 236188 74898 241882 75134
rect 242118 74898 247813 75134
rect 248049 74898 262952 75134
rect 263188 74898 268882 75134
rect 269118 74898 274813 75134
rect 275049 74898 289952 75134
rect 290188 74898 295882 75134
rect 296118 74898 301813 75134
rect 302049 74898 316952 75134
rect 317188 74898 322882 75134
rect 323118 74898 328813 75134
rect 329049 74898 343952 75134
rect 344188 74898 349882 75134
rect 350118 74898 355813 75134
rect 356049 74898 370952 75134
rect 371188 74898 376882 75134
rect 377118 74898 382813 75134
rect 383049 74898 397952 75134
rect 398188 74898 403882 75134
rect 404118 74898 409813 75134
rect 410049 74898 424952 75134
rect 425188 74898 430882 75134
rect 431118 74898 436813 75134
rect 437049 74898 451952 75134
rect 452188 74898 457882 75134
rect 458118 74898 463813 75134
rect 464049 74898 478952 75134
rect 479188 74898 484882 75134
rect 485118 74898 490813 75134
rect 491049 74898 505952 75134
rect 506188 74898 511882 75134
rect 512118 74898 517813 75134
rect 518049 74898 532952 75134
rect 533188 74898 538882 75134
rect 539118 74898 544813 75134
rect 545049 74898 559826 75134
rect 560062 74898 560146 75134
rect 560382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect 19794 67394 542414 67426
rect 19794 67158 19826 67394
rect 20062 67158 20146 67394
rect 20382 67158 37826 67394
rect 38062 67158 38146 67394
rect 38382 67158 55826 67394
rect 56062 67158 56146 67394
rect 56382 67158 73826 67394
rect 74062 67158 74146 67394
rect 74382 67158 91826 67394
rect 92062 67158 92146 67394
rect 92382 67158 109826 67394
rect 110062 67158 110146 67394
rect 110382 67158 127826 67394
rect 128062 67158 128146 67394
rect 128382 67158 145826 67394
rect 146062 67158 146146 67394
rect 146382 67158 163826 67394
rect 164062 67158 164146 67394
rect 164382 67158 181826 67394
rect 182062 67158 182146 67394
rect 182382 67158 199826 67394
rect 200062 67158 200146 67394
rect 200382 67158 217826 67394
rect 218062 67158 218146 67394
rect 218382 67158 235826 67394
rect 236062 67158 236146 67394
rect 236382 67158 253826 67394
rect 254062 67158 254146 67394
rect 254382 67158 271826 67394
rect 272062 67158 272146 67394
rect 272382 67158 289826 67394
rect 290062 67158 290146 67394
rect 290382 67158 307826 67394
rect 308062 67158 308146 67394
rect 308382 67158 325826 67394
rect 326062 67158 326146 67394
rect 326382 67158 343826 67394
rect 344062 67158 344146 67394
rect 344382 67158 361826 67394
rect 362062 67158 362146 67394
rect 362382 67158 379826 67394
rect 380062 67158 380146 67394
rect 380382 67158 397826 67394
rect 398062 67158 398146 67394
rect 398382 67158 415826 67394
rect 416062 67158 416146 67394
rect 416382 67158 433826 67394
rect 434062 67158 434146 67394
rect 434382 67158 451826 67394
rect 452062 67158 452146 67394
rect 452382 67158 469826 67394
rect 470062 67158 470146 67394
rect 470382 67158 487826 67394
rect 488062 67158 488146 67394
rect 488382 67158 505826 67394
rect 506062 67158 506146 67394
rect 506382 67158 523826 67394
rect 524062 67158 524146 67394
rect 524382 67158 541826 67394
rect 542062 67158 542146 67394
rect 542382 67158 542414 67394
rect 19794 67074 542414 67158
rect 19794 66838 19826 67074
rect 20062 66838 20146 67074
rect 20382 66838 37826 67074
rect 38062 66838 38146 67074
rect 38382 66838 55826 67074
rect 56062 66838 56146 67074
rect 56382 66838 73826 67074
rect 74062 66838 74146 67074
rect 74382 66838 91826 67074
rect 92062 66838 92146 67074
rect 92382 66838 109826 67074
rect 110062 66838 110146 67074
rect 110382 66838 127826 67074
rect 128062 66838 128146 67074
rect 128382 66838 145826 67074
rect 146062 66838 146146 67074
rect 146382 66838 163826 67074
rect 164062 66838 164146 67074
rect 164382 66838 181826 67074
rect 182062 66838 182146 67074
rect 182382 66838 199826 67074
rect 200062 66838 200146 67074
rect 200382 66838 217826 67074
rect 218062 66838 218146 67074
rect 218382 66838 235826 67074
rect 236062 66838 236146 67074
rect 236382 66838 253826 67074
rect 254062 66838 254146 67074
rect 254382 66838 271826 67074
rect 272062 66838 272146 67074
rect 272382 66838 289826 67074
rect 290062 66838 290146 67074
rect 290382 66838 307826 67074
rect 308062 66838 308146 67074
rect 308382 66838 325826 67074
rect 326062 66838 326146 67074
rect 326382 66838 343826 67074
rect 344062 66838 344146 67074
rect 344382 66838 361826 67074
rect 362062 66838 362146 67074
rect 362382 66838 379826 67074
rect 380062 66838 380146 67074
rect 380382 66838 397826 67074
rect 398062 66838 398146 67074
rect 398382 66838 415826 67074
rect 416062 66838 416146 67074
rect 416382 66838 433826 67074
rect 434062 66838 434146 67074
rect 434382 66838 451826 67074
rect 452062 66838 452146 67074
rect 452382 66838 469826 67074
rect 470062 66838 470146 67074
rect 470382 66838 487826 67074
rect 488062 66838 488146 67074
rect 488382 66838 505826 67074
rect 506062 66838 506146 67074
rect 506382 66838 523826 67074
rect 524062 66838 524146 67074
rect 524382 66838 541826 67074
rect 542062 66838 542146 67074
rect 542382 66838 542414 67074
rect 19794 66806 542414 66838
rect -2966 66454 586890 66486
rect -2966 66218 -2934 66454
rect -2698 66218 -2614 66454
rect -2378 66218 10826 66454
rect 11062 66218 11146 66454
rect 11382 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 46826 66454
rect 47062 66218 47146 66454
rect 47382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 82826 66454
rect 83062 66218 83146 66454
rect 83382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 118826 66454
rect 119062 66218 119146 66454
rect 119382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 154826 66454
rect 155062 66218 155146 66454
rect 155382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 190826 66454
rect 191062 66218 191146 66454
rect 191382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 226826 66454
rect 227062 66218 227146 66454
rect 227382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 262826 66454
rect 263062 66218 263146 66454
rect 263382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 298826 66454
rect 299062 66218 299146 66454
rect 299382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 334826 66454
rect 335062 66218 335146 66454
rect 335382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 370826 66454
rect 371062 66218 371146 66454
rect 371382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 406826 66454
rect 407062 66218 407146 66454
rect 407382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 442826 66454
rect 443062 66218 443146 66454
rect 443382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 478826 66454
rect 479062 66218 479146 66454
rect 479382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 514826 66454
rect 515062 66218 515146 66454
rect 515382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 550826 66454
rect 551062 66218 551146 66454
rect 551382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 586302 66454
rect 586538 66218 586622 66454
rect 586858 66218 586890 66454
rect -2966 66134 586890 66218
rect -2966 65898 -2934 66134
rect -2698 65898 -2614 66134
rect -2378 65898 10826 66134
rect 11062 65898 11146 66134
rect 11382 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 46826 66134
rect 47062 65898 47146 66134
rect 47382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 82826 66134
rect 83062 65898 83146 66134
rect 83382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 118826 66134
rect 119062 65898 119146 66134
rect 119382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 154826 66134
rect 155062 65898 155146 66134
rect 155382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 190826 66134
rect 191062 65898 191146 66134
rect 191382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 226826 66134
rect 227062 65898 227146 66134
rect 227382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 262826 66134
rect 263062 65898 263146 66134
rect 263382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 298826 66134
rect 299062 65898 299146 66134
rect 299382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 334826 66134
rect 335062 65898 335146 66134
rect 335382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 370826 66134
rect 371062 65898 371146 66134
rect 371382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 406826 66134
rect 407062 65898 407146 66134
rect 407382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 442826 66134
rect 443062 65898 443146 66134
rect 443382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 478826 66134
rect 479062 65898 479146 66134
rect 479382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 514826 66134
rect 515062 65898 515146 66134
rect 515382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 550826 66134
rect 551062 65898 551146 66134
rect 551382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 586302 66134
rect 586538 65898 586622 66134
rect 586858 65898 586890 66134
rect -2966 65866 586890 65898
rect -2966 57454 586890 57486
rect -2966 57218 -1974 57454
rect -1738 57218 -1654 57454
rect -1418 57218 1826 57454
rect 2062 57218 2146 57454
rect 2382 57218 19952 57454
rect 20188 57218 25882 57454
rect 26118 57218 31813 57454
rect 32049 57218 46952 57454
rect 47188 57218 52882 57454
rect 53118 57218 58813 57454
rect 59049 57218 73952 57454
rect 74188 57218 79882 57454
rect 80118 57218 85813 57454
rect 86049 57218 100952 57454
rect 101188 57218 106882 57454
rect 107118 57218 112813 57454
rect 113049 57218 127952 57454
rect 128188 57218 133882 57454
rect 134118 57218 139813 57454
rect 140049 57218 154952 57454
rect 155188 57218 160882 57454
rect 161118 57218 166813 57454
rect 167049 57218 181952 57454
rect 182188 57218 187882 57454
rect 188118 57218 193813 57454
rect 194049 57218 208952 57454
rect 209188 57218 214882 57454
rect 215118 57218 220813 57454
rect 221049 57218 235952 57454
rect 236188 57218 241882 57454
rect 242118 57218 247813 57454
rect 248049 57218 262952 57454
rect 263188 57218 268882 57454
rect 269118 57218 274813 57454
rect 275049 57218 289952 57454
rect 290188 57218 295882 57454
rect 296118 57218 301813 57454
rect 302049 57218 316952 57454
rect 317188 57218 322882 57454
rect 323118 57218 328813 57454
rect 329049 57218 343952 57454
rect 344188 57218 349882 57454
rect 350118 57218 355813 57454
rect 356049 57218 370952 57454
rect 371188 57218 376882 57454
rect 377118 57218 382813 57454
rect 383049 57218 397952 57454
rect 398188 57218 403882 57454
rect 404118 57218 409813 57454
rect 410049 57218 424952 57454
rect 425188 57218 430882 57454
rect 431118 57218 436813 57454
rect 437049 57218 451952 57454
rect 452188 57218 457882 57454
rect 458118 57218 463813 57454
rect 464049 57218 478952 57454
rect 479188 57218 484882 57454
rect 485118 57218 490813 57454
rect 491049 57218 505952 57454
rect 506188 57218 511882 57454
rect 512118 57218 517813 57454
rect 518049 57218 532952 57454
rect 533188 57218 538882 57454
rect 539118 57218 544813 57454
rect 545049 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 577826 57454
rect 578062 57218 578146 57454
rect 578382 57218 585342 57454
rect 585578 57218 585662 57454
rect 585898 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -1974 57134
rect -1738 56898 -1654 57134
rect -1418 56898 1826 57134
rect 2062 56898 2146 57134
rect 2382 56898 19952 57134
rect 20188 56898 25882 57134
rect 26118 56898 31813 57134
rect 32049 56898 46952 57134
rect 47188 56898 52882 57134
rect 53118 56898 58813 57134
rect 59049 56898 73952 57134
rect 74188 56898 79882 57134
rect 80118 56898 85813 57134
rect 86049 56898 100952 57134
rect 101188 56898 106882 57134
rect 107118 56898 112813 57134
rect 113049 56898 127952 57134
rect 128188 56898 133882 57134
rect 134118 56898 139813 57134
rect 140049 56898 154952 57134
rect 155188 56898 160882 57134
rect 161118 56898 166813 57134
rect 167049 56898 181952 57134
rect 182188 56898 187882 57134
rect 188118 56898 193813 57134
rect 194049 56898 208952 57134
rect 209188 56898 214882 57134
rect 215118 56898 220813 57134
rect 221049 56898 235952 57134
rect 236188 56898 241882 57134
rect 242118 56898 247813 57134
rect 248049 56898 262952 57134
rect 263188 56898 268882 57134
rect 269118 56898 274813 57134
rect 275049 56898 289952 57134
rect 290188 56898 295882 57134
rect 296118 56898 301813 57134
rect 302049 56898 316952 57134
rect 317188 56898 322882 57134
rect 323118 56898 328813 57134
rect 329049 56898 343952 57134
rect 344188 56898 349882 57134
rect 350118 56898 355813 57134
rect 356049 56898 370952 57134
rect 371188 56898 376882 57134
rect 377118 56898 382813 57134
rect 383049 56898 397952 57134
rect 398188 56898 403882 57134
rect 404118 56898 409813 57134
rect 410049 56898 424952 57134
rect 425188 56898 430882 57134
rect 431118 56898 436813 57134
rect 437049 56898 451952 57134
rect 452188 56898 457882 57134
rect 458118 56898 463813 57134
rect 464049 56898 478952 57134
rect 479188 56898 484882 57134
rect 485118 56898 490813 57134
rect 491049 56898 505952 57134
rect 506188 56898 511882 57134
rect 512118 56898 517813 57134
rect 518049 56898 532952 57134
rect 533188 56898 538882 57134
rect 539118 56898 544813 57134
rect 545049 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 577826 57134
rect 578062 56898 578146 57134
rect 578382 56898 585342 57134
rect 585578 56898 585662 57134
rect 585898 56898 586890 57134
rect -2966 56866 586890 56898
rect -2966 48454 586890 48486
rect -2966 48218 -2934 48454
rect -2698 48218 -2614 48454
rect -2378 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 22916 48454
rect 23152 48218 28847 48454
rect 29083 48218 49916 48454
rect 50152 48218 55847 48454
rect 56083 48218 76916 48454
rect 77152 48218 82847 48454
rect 83083 48218 103916 48454
rect 104152 48218 109847 48454
rect 110083 48218 130916 48454
rect 131152 48218 136847 48454
rect 137083 48218 157916 48454
rect 158152 48218 163847 48454
rect 164083 48218 184916 48454
rect 185152 48218 190847 48454
rect 191083 48218 211916 48454
rect 212152 48218 217847 48454
rect 218083 48218 238916 48454
rect 239152 48218 244847 48454
rect 245083 48218 265916 48454
rect 266152 48218 271847 48454
rect 272083 48218 292916 48454
rect 293152 48218 298847 48454
rect 299083 48218 319916 48454
rect 320152 48218 325847 48454
rect 326083 48218 346916 48454
rect 347152 48218 352847 48454
rect 353083 48218 373916 48454
rect 374152 48218 379847 48454
rect 380083 48218 400916 48454
rect 401152 48218 406847 48454
rect 407083 48218 427916 48454
rect 428152 48218 433847 48454
rect 434083 48218 454916 48454
rect 455152 48218 460847 48454
rect 461083 48218 481916 48454
rect 482152 48218 487847 48454
rect 488083 48218 508916 48454
rect 509152 48218 514847 48454
rect 515083 48218 535916 48454
rect 536152 48218 541847 48454
rect 542083 48218 568826 48454
rect 569062 48218 569146 48454
rect 569382 48218 586302 48454
rect 586538 48218 586622 48454
rect 586858 48218 586890 48454
rect -2966 48134 586890 48218
rect -2966 47898 -2934 48134
rect -2698 47898 -2614 48134
rect -2378 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 22916 48134
rect 23152 47898 28847 48134
rect 29083 47898 49916 48134
rect 50152 47898 55847 48134
rect 56083 47898 76916 48134
rect 77152 47898 82847 48134
rect 83083 47898 103916 48134
rect 104152 47898 109847 48134
rect 110083 47898 130916 48134
rect 131152 47898 136847 48134
rect 137083 47898 157916 48134
rect 158152 47898 163847 48134
rect 164083 47898 184916 48134
rect 185152 47898 190847 48134
rect 191083 47898 211916 48134
rect 212152 47898 217847 48134
rect 218083 47898 238916 48134
rect 239152 47898 244847 48134
rect 245083 47898 265916 48134
rect 266152 47898 271847 48134
rect 272083 47898 292916 48134
rect 293152 47898 298847 48134
rect 299083 47898 319916 48134
rect 320152 47898 325847 48134
rect 326083 47898 346916 48134
rect 347152 47898 352847 48134
rect 353083 47898 373916 48134
rect 374152 47898 379847 48134
rect 380083 47898 400916 48134
rect 401152 47898 406847 48134
rect 407083 47898 427916 48134
rect 428152 47898 433847 48134
rect 434083 47898 454916 48134
rect 455152 47898 460847 48134
rect 461083 47898 481916 48134
rect 482152 47898 487847 48134
rect 488083 47898 508916 48134
rect 509152 47898 514847 48134
rect 515083 47898 535916 48134
rect 536152 47898 541847 48134
rect 542083 47898 568826 48134
rect 569062 47898 569146 48134
rect 569382 47898 586302 48134
rect 586538 47898 586622 48134
rect 586858 47898 586890 48134
rect -2966 47866 586890 47898
rect 28794 40394 551414 40426
rect 28794 40158 28826 40394
rect 29062 40158 29146 40394
rect 29382 40158 46826 40394
rect 47062 40158 47146 40394
rect 47382 40158 64826 40394
rect 65062 40158 65146 40394
rect 65382 40158 82826 40394
rect 83062 40158 83146 40394
rect 83382 40158 100826 40394
rect 101062 40158 101146 40394
rect 101382 40158 118826 40394
rect 119062 40158 119146 40394
rect 119382 40158 136826 40394
rect 137062 40158 137146 40394
rect 137382 40158 154826 40394
rect 155062 40158 155146 40394
rect 155382 40158 172826 40394
rect 173062 40158 173146 40394
rect 173382 40158 190826 40394
rect 191062 40158 191146 40394
rect 191382 40158 208826 40394
rect 209062 40158 209146 40394
rect 209382 40158 226826 40394
rect 227062 40158 227146 40394
rect 227382 40158 244826 40394
rect 245062 40158 245146 40394
rect 245382 40158 262826 40394
rect 263062 40158 263146 40394
rect 263382 40158 280826 40394
rect 281062 40158 281146 40394
rect 281382 40158 298826 40394
rect 299062 40158 299146 40394
rect 299382 40158 316826 40394
rect 317062 40158 317146 40394
rect 317382 40158 334826 40394
rect 335062 40158 335146 40394
rect 335382 40158 352826 40394
rect 353062 40158 353146 40394
rect 353382 40158 370826 40394
rect 371062 40158 371146 40394
rect 371382 40158 388826 40394
rect 389062 40158 389146 40394
rect 389382 40158 406826 40394
rect 407062 40158 407146 40394
rect 407382 40158 424826 40394
rect 425062 40158 425146 40394
rect 425382 40158 442826 40394
rect 443062 40158 443146 40394
rect 443382 40158 460826 40394
rect 461062 40158 461146 40394
rect 461382 40158 478826 40394
rect 479062 40158 479146 40394
rect 479382 40158 496826 40394
rect 497062 40158 497146 40394
rect 497382 40158 514826 40394
rect 515062 40158 515146 40394
rect 515382 40158 532826 40394
rect 533062 40158 533146 40394
rect 533382 40158 550826 40394
rect 551062 40158 551146 40394
rect 551382 40158 551414 40394
rect 28794 40074 551414 40158
rect 28794 39838 28826 40074
rect 29062 39838 29146 40074
rect 29382 39838 46826 40074
rect 47062 39838 47146 40074
rect 47382 39838 64826 40074
rect 65062 39838 65146 40074
rect 65382 39838 82826 40074
rect 83062 39838 83146 40074
rect 83382 39838 100826 40074
rect 101062 39838 101146 40074
rect 101382 39838 118826 40074
rect 119062 39838 119146 40074
rect 119382 39838 136826 40074
rect 137062 39838 137146 40074
rect 137382 39838 154826 40074
rect 155062 39838 155146 40074
rect 155382 39838 172826 40074
rect 173062 39838 173146 40074
rect 173382 39838 190826 40074
rect 191062 39838 191146 40074
rect 191382 39838 208826 40074
rect 209062 39838 209146 40074
rect 209382 39838 226826 40074
rect 227062 39838 227146 40074
rect 227382 39838 244826 40074
rect 245062 39838 245146 40074
rect 245382 39838 262826 40074
rect 263062 39838 263146 40074
rect 263382 39838 280826 40074
rect 281062 39838 281146 40074
rect 281382 39838 298826 40074
rect 299062 39838 299146 40074
rect 299382 39838 316826 40074
rect 317062 39838 317146 40074
rect 317382 39838 334826 40074
rect 335062 39838 335146 40074
rect 335382 39838 352826 40074
rect 353062 39838 353146 40074
rect 353382 39838 370826 40074
rect 371062 39838 371146 40074
rect 371382 39838 388826 40074
rect 389062 39838 389146 40074
rect 389382 39838 406826 40074
rect 407062 39838 407146 40074
rect 407382 39838 424826 40074
rect 425062 39838 425146 40074
rect 425382 39838 442826 40074
rect 443062 39838 443146 40074
rect 443382 39838 460826 40074
rect 461062 39838 461146 40074
rect 461382 39838 478826 40074
rect 479062 39838 479146 40074
rect 479382 39838 496826 40074
rect 497062 39838 497146 40074
rect 497382 39838 514826 40074
rect 515062 39838 515146 40074
rect 515382 39838 532826 40074
rect 533062 39838 533146 40074
rect 533382 39838 550826 40074
rect 551062 39838 551146 40074
rect 551382 39838 551414 40074
rect 28794 39806 551414 39838
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 19826 39454
rect 20062 39218 20146 39454
rect 20382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 55826 39454
rect 56062 39218 56146 39454
rect 56382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 91826 39454
rect 92062 39218 92146 39454
rect 92382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 127826 39454
rect 128062 39218 128146 39454
rect 128382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 163826 39454
rect 164062 39218 164146 39454
rect 164382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 199826 39454
rect 200062 39218 200146 39454
rect 200382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 235826 39454
rect 236062 39218 236146 39454
rect 236382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 271826 39454
rect 272062 39218 272146 39454
rect 272382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 307826 39454
rect 308062 39218 308146 39454
rect 308382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 343826 39454
rect 344062 39218 344146 39454
rect 344382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 379826 39454
rect 380062 39218 380146 39454
rect 380382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 415826 39454
rect 416062 39218 416146 39454
rect 416382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 451826 39454
rect 452062 39218 452146 39454
rect 452382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 487826 39454
rect 488062 39218 488146 39454
rect 488382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 523826 39454
rect 524062 39218 524146 39454
rect 524382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 559826 39454
rect 560062 39218 560146 39454
rect 560382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 19826 39134
rect 20062 38898 20146 39134
rect 20382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 55826 39134
rect 56062 38898 56146 39134
rect 56382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 91826 39134
rect 92062 38898 92146 39134
rect 92382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 127826 39134
rect 128062 38898 128146 39134
rect 128382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 163826 39134
rect 164062 38898 164146 39134
rect 164382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 199826 39134
rect 200062 38898 200146 39134
rect 200382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 235826 39134
rect 236062 38898 236146 39134
rect 236382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 271826 39134
rect 272062 38898 272146 39134
rect 272382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 307826 39134
rect 308062 38898 308146 39134
rect 308382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 343826 39134
rect 344062 38898 344146 39134
rect 344382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 379826 39134
rect 380062 38898 380146 39134
rect 380382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 415826 39134
rect 416062 38898 416146 39134
rect 416382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 451826 39134
rect 452062 38898 452146 39134
rect 452382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 487826 39134
rect 488062 38898 488146 39134
rect 488382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 523826 39134
rect 524062 38898 524146 39134
rect 524382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 559826 39134
rect 560062 38898 560146 39134
rect 560382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -2966 30454 586890 30486
rect -2966 30218 -2934 30454
rect -2698 30218 -2614 30454
rect -2378 30218 10826 30454
rect 11062 30218 11146 30454
rect 11382 30218 22916 30454
rect 23152 30218 28847 30454
rect 29083 30218 49916 30454
rect 50152 30218 55847 30454
rect 56083 30218 76916 30454
rect 77152 30218 82847 30454
rect 83083 30218 103916 30454
rect 104152 30218 109847 30454
rect 110083 30218 130916 30454
rect 131152 30218 136847 30454
rect 137083 30218 157916 30454
rect 158152 30218 163847 30454
rect 164083 30218 184916 30454
rect 185152 30218 190847 30454
rect 191083 30218 211916 30454
rect 212152 30218 217847 30454
rect 218083 30218 238916 30454
rect 239152 30218 244847 30454
rect 245083 30218 265916 30454
rect 266152 30218 271847 30454
rect 272083 30218 292916 30454
rect 293152 30218 298847 30454
rect 299083 30218 319916 30454
rect 320152 30218 325847 30454
rect 326083 30218 346916 30454
rect 347152 30218 352847 30454
rect 353083 30218 373916 30454
rect 374152 30218 379847 30454
rect 380083 30218 400916 30454
rect 401152 30218 406847 30454
rect 407083 30218 427916 30454
rect 428152 30218 433847 30454
rect 434083 30218 454916 30454
rect 455152 30218 460847 30454
rect 461083 30218 481916 30454
rect 482152 30218 487847 30454
rect 488083 30218 508916 30454
rect 509152 30218 514847 30454
rect 515083 30218 535916 30454
rect 536152 30218 541847 30454
rect 542083 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 586302 30454
rect 586538 30218 586622 30454
rect 586858 30218 586890 30454
rect -2966 30134 586890 30218
rect -2966 29898 -2934 30134
rect -2698 29898 -2614 30134
rect -2378 29898 10826 30134
rect 11062 29898 11146 30134
rect 11382 29898 22916 30134
rect 23152 29898 28847 30134
rect 29083 29898 49916 30134
rect 50152 29898 55847 30134
rect 56083 29898 76916 30134
rect 77152 29898 82847 30134
rect 83083 29898 103916 30134
rect 104152 29898 109847 30134
rect 110083 29898 130916 30134
rect 131152 29898 136847 30134
rect 137083 29898 157916 30134
rect 158152 29898 163847 30134
rect 164083 29898 184916 30134
rect 185152 29898 190847 30134
rect 191083 29898 211916 30134
rect 212152 29898 217847 30134
rect 218083 29898 238916 30134
rect 239152 29898 244847 30134
rect 245083 29898 265916 30134
rect 266152 29898 271847 30134
rect 272083 29898 292916 30134
rect 293152 29898 298847 30134
rect 299083 29898 319916 30134
rect 320152 29898 325847 30134
rect 326083 29898 346916 30134
rect 347152 29898 352847 30134
rect 353083 29898 373916 30134
rect 374152 29898 379847 30134
rect 380083 29898 400916 30134
rect 401152 29898 406847 30134
rect 407083 29898 427916 30134
rect 428152 29898 433847 30134
rect 434083 29898 454916 30134
rect 455152 29898 460847 30134
rect 461083 29898 481916 30134
rect 482152 29898 487847 30134
rect 488083 29898 508916 30134
rect 509152 29898 514847 30134
rect 515083 29898 535916 30134
rect 536152 29898 541847 30134
rect 542083 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 586302 30134
rect 586538 29898 586622 30134
rect 586858 29898 586890 30134
rect -2966 29866 586890 29898
rect -2966 21454 586890 21486
rect -2966 21218 -1974 21454
rect -1738 21218 -1654 21454
rect -1418 21218 1826 21454
rect 2062 21218 2146 21454
rect 2382 21218 19952 21454
rect 20188 21218 25882 21454
rect 26118 21218 31813 21454
rect 32049 21218 46952 21454
rect 47188 21218 52882 21454
rect 53118 21218 58813 21454
rect 59049 21218 73952 21454
rect 74188 21218 79882 21454
rect 80118 21218 85813 21454
rect 86049 21218 100952 21454
rect 101188 21218 106882 21454
rect 107118 21218 112813 21454
rect 113049 21218 127952 21454
rect 128188 21218 133882 21454
rect 134118 21218 139813 21454
rect 140049 21218 154952 21454
rect 155188 21218 160882 21454
rect 161118 21218 166813 21454
rect 167049 21218 181952 21454
rect 182188 21218 187882 21454
rect 188118 21218 193813 21454
rect 194049 21218 208952 21454
rect 209188 21218 214882 21454
rect 215118 21218 220813 21454
rect 221049 21218 235952 21454
rect 236188 21218 241882 21454
rect 242118 21218 247813 21454
rect 248049 21218 262952 21454
rect 263188 21218 268882 21454
rect 269118 21218 274813 21454
rect 275049 21218 289952 21454
rect 290188 21218 295882 21454
rect 296118 21218 301813 21454
rect 302049 21218 316952 21454
rect 317188 21218 322882 21454
rect 323118 21218 328813 21454
rect 329049 21218 343952 21454
rect 344188 21218 349882 21454
rect 350118 21218 355813 21454
rect 356049 21218 370952 21454
rect 371188 21218 376882 21454
rect 377118 21218 382813 21454
rect 383049 21218 397952 21454
rect 398188 21218 403882 21454
rect 404118 21218 409813 21454
rect 410049 21218 424952 21454
rect 425188 21218 430882 21454
rect 431118 21218 436813 21454
rect 437049 21218 451952 21454
rect 452188 21218 457882 21454
rect 458118 21218 463813 21454
rect 464049 21218 478952 21454
rect 479188 21218 484882 21454
rect 485118 21218 490813 21454
rect 491049 21218 505952 21454
rect 506188 21218 511882 21454
rect 512118 21218 517813 21454
rect 518049 21218 532952 21454
rect 533188 21218 538882 21454
rect 539118 21218 544813 21454
rect 545049 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 577826 21454
rect 578062 21218 578146 21454
rect 578382 21218 585342 21454
rect 585578 21218 585662 21454
rect 585898 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -1974 21134
rect -1738 20898 -1654 21134
rect -1418 20898 1826 21134
rect 2062 20898 2146 21134
rect 2382 20898 19952 21134
rect 20188 20898 25882 21134
rect 26118 20898 31813 21134
rect 32049 20898 46952 21134
rect 47188 20898 52882 21134
rect 53118 20898 58813 21134
rect 59049 20898 73952 21134
rect 74188 20898 79882 21134
rect 80118 20898 85813 21134
rect 86049 20898 100952 21134
rect 101188 20898 106882 21134
rect 107118 20898 112813 21134
rect 113049 20898 127952 21134
rect 128188 20898 133882 21134
rect 134118 20898 139813 21134
rect 140049 20898 154952 21134
rect 155188 20898 160882 21134
rect 161118 20898 166813 21134
rect 167049 20898 181952 21134
rect 182188 20898 187882 21134
rect 188118 20898 193813 21134
rect 194049 20898 208952 21134
rect 209188 20898 214882 21134
rect 215118 20898 220813 21134
rect 221049 20898 235952 21134
rect 236188 20898 241882 21134
rect 242118 20898 247813 21134
rect 248049 20898 262952 21134
rect 263188 20898 268882 21134
rect 269118 20898 274813 21134
rect 275049 20898 289952 21134
rect 290188 20898 295882 21134
rect 296118 20898 301813 21134
rect 302049 20898 316952 21134
rect 317188 20898 322882 21134
rect 323118 20898 328813 21134
rect 329049 20898 343952 21134
rect 344188 20898 349882 21134
rect 350118 20898 355813 21134
rect 356049 20898 370952 21134
rect 371188 20898 376882 21134
rect 377118 20898 382813 21134
rect 383049 20898 397952 21134
rect 398188 20898 403882 21134
rect 404118 20898 409813 21134
rect 410049 20898 424952 21134
rect 425188 20898 430882 21134
rect 431118 20898 436813 21134
rect 437049 20898 451952 21134
rect 452188 20898 457882 21134
rect 458118 20898 463813 21134
rect 464049 20898 478952 21134
rect 479188 20898 484882 21134
rect 485118 20898 490813 21134
rect 491049 20898 505952 21134
rect 506188 20898 511882 21134
rect 512118 20898 517813 21134
rect 518049 20898 532952 21134
rect 533188 20898 538882 21134
rect 539118 20898 544813 21134
rect 545049 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 577826 21134
rect 578062 20898 578146 21134
rect 578382 20898 585342 21134
rect 585578 20898 585662 21134
rect 585898 20898 586890 21134
rect -2966 20866 586890 20898
rect -2966 12454 586890 12486
rect -2966 12218 -2934 12454
rect -2698 12218 -2614 12454
rect -2378 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 28826 12454
rect 29062 12218 29146 12454
rect 29382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 64826 12454
rect 65062 12218 65146 12454
rect 65382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 100826 12454
rect 101062 12218 101146 12454
rect 101382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 136826 12454
rect 137062 12218 137146 12454
rect 137382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 172826 12454
rect 173062 12218 173146 12454
rect 173382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 208826 12454
rect 209062 12218 209146 12454
rect 209382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 244826 12454
rect 245062 12218 245146 12454
rect 245382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 280826 12454
rect 281062 12218 281146 12454
rect 281382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 316826 12454
rect 317062 12218 317146 12454
rect 317382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 352826 12454
rect 353062 12218 353146 12454
rect 353382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 388826 12454
rect 389062 12218 389146 12454
rect 389382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 424826 12454
rect 425062 12218 425146 12454
rect 425382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 460826 12454
rect 461062 12218 461146 12454
rect 461382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 496826 12454
rect 497062 12218 497146 12454
rect 497382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 532826 12454
rect 533062 12218 533146 12454
rect 533382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 568826 12454
rect 569062 12218 569146 12454
rect 569382 12218 586302 12454
rect 586538 12218 586622 12454
rect 586858 12218 586890 12454
rect -2966 12134 586890 12218
rect -2966 11898 -2934 12134
rect -2698 11898 -2614 12134
rect -2378 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 28826 12134
rect 29062 11898 29146 12134
rect 29382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 64826 12134
rect 65062 11898 65146 12134
rect 65382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 100826 12134
rect 101062 11898 101146 12134
rect 101382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 136826 12134
rect 137062 11898 137146 12134
rect 137382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 172826 12134
rect 173062 11898 173146 12134
rect 173382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 208826 12134
rect 209062 11898 209146 12134
rect 209382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 244826 12134
rect 245062 11898 245146 12134
rect 245382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 280826 12134
rect 281062 11898 281146 12134
rect 281382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 316826 12134
rect 317062 11898 317146 12134
rect 317382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 352826 12134
rect 353062 11898 353146 12134
rect 353382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 388826 12134
rect 389062 11898 389146 12134
rect 389382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 424826 12134
rect 425062 11898 425146 12134
rect 425382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 460826 12134
rect 461062 11898 461146 12134
rect 461382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 496826 12134
rect 497062 11898 497146 12134
rect 497382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 532826 12134
rect 533062 11898 533146 12134
rect 533382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 568826 12134
rect 569062 11898 569146 12134
rect 569382 11898 586302 12134
rect 586538 11898 586622 12134
rect 586858 11898 586890 12134
rect -2966 11866 586890 11898
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 19826 3454
rect 20062 3218 20146 3454
rect 20382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 55826 3454
rect 56062 3218 56146 3454
rect 56382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 91826 3454
rect 92062 3218 92146 3454
rect 92382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 127826 3454
rect 128062 3218 128146 3454
rect 128382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 163826 3454
rect 164062 3218 164146 3454
rect 164382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 199826 3454
rect 200062 3218 200146 3454
rect 200382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 235826 3454
rect 236062 3218 236146 3454
rect 236382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 271826 3454
rect 272062 3218 272146 3454
rect 272382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 307826 3454
rect 308062 3218 308146 3454
rect 308382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 343826 3454
rect 344062 3218 344146 3454
rect 344382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 379826 3454
rect 380062 3218 380146 3454
rect 380382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 415826 3454
rect 416062 3218 416146 3454
rect 416382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 451826 3454
rect 452062 3218 452146 3454
rect 452382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 487826 3454
rect 488062 3218 488146 3454
rect 488382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 523826 3454
rect 524062 3218 524146 3454
rect 524382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 559826 3454
rect 560062 3218 560146 3454
rect 560382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 19826 3134
rect 20062 2898 20146 3134
rect 20382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 55826 3134
rect 56062 2898 56146 3134
rect 56382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 91826 3134
rect 92062 2898 92146 3134
rect 92382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 127826 3134
rect 128062 2898 128146 3134
rect 128382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 163826 3134
rect 164062 2898 164146 3134
rect 164382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 199826 3134
rect 200062 2898 200146 3134
rect 200382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 235826 3134
rect 236062 2898 236146 3134
rect 236382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 271826 3134
rect 272062 2898 272146 3134
rect 272382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 307826 3134
rect 308062 2898 308146 3134
rect 308382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 343826 3134
rect 344062 2898 344146 3134
rect 344382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 379826 3134
rect 380062 2898 380146 3134
rect 380382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 415826 3134
rect 416062 2898 416146 3134
rect 416382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 451826 3134
rect 452062 2898 452146 3134
rect 452382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 487826 3134
rect 488062 2898 488146 3134
rect 488382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 523826 3134
rect 524062 2898 524146 3134
rect 524382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 559826 3134
rect 560062 2898 560146 3134
rect 560382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 19826 -346
rect 20062 -582 20146 -346
rect 20382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 55826 -346
rect 56062 -582 56146 -346
rect 56382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 91826 -346
rect 92062 -582 92146 -346
rect 92382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 127826 -346
rect 128062 -582 128146 -346
rect 128382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 163826 -346
rect 164062 -582 164146 -346
rect 164382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 199826 -346
rect 200062 -582 200146 -346
rect 200382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 235826 -346
rect 236062 -582 236146 -346
rect 236382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 271826 -346
rect 272062 -582 272146 -346
rect 272382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 307826 -346
rect 308062 -582 308146 -346
rect 308382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 343826 -346
rect 344062 -582 344146 -346
rect 344382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 379826 -346
rect 380062 -582 380146 -346
rect 380382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 415826 -346
rect 416062 -582 416146 -346
rect 416382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 451826 -346
rect 452062 -582 452146 -346
rect 452382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 487826 -346
rect 488062 -582 488146 -346
rect 488382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 523826 -346
rect 524062 -582 524146 -346
rect 524382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 559826 -346
rect 560062 -582 560146 -346
rect 560382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 19826 -666
rect 20062 -902 20146 -666
rect 20382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 55826 -666
rect 56062 -902 56146 -666
rect 56382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 91826 -666
rect 92062 -902 92146 -666
rect 92382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 127826 -666
rect 128062 -902 128146 -666
rect 128382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 163826 -666
rect 164062 -902 164146 -666
rect 164382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 199826 -666
rect 200062 -902 200146 -666
rect 200382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 235826 -666
rect 236062 -902 236146 -666
rect 236382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 271826 -666
rect 272062 -902 272146 -666
rect 272382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 307826 -666
rect 308062 -902 308146 -666
rect 308382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 343826 -666
rect 344062 -902 344146 -666
rect 344382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 379826 -666
rect 380062 -902 380146 -666
rect 380382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 415826 -666
rect 416062 -902 416146 -666
rect 416382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 451826 -666
rect 452062 -902 452146 -666
rect 452382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 487826 -666
rect 488062 -902 488146 -666
rect 488382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 523826 -666
rect 524062 -902 524146 -666
rect 524382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 559826 -666
rect 560062 -902 560146 -666
rect 560382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 10826 -1306
rect 11062 -1542 11146 -1306
rect 11382 -1542 28826 -1306
rect 29062 -1542 29146 -1306
rect 29382 -1542 46826 -1306
rect 47062 -1542 47146 -1306
rect 47382 -1542 64826 -1306
rect 65062 -1542 65146 -1306
rect 65382 -1542 82826 -1306
rect 83062 -1542 83146 -1306
rect 83382 -1542 100826 -1306
rect 101062 -1542 101146 -1306
rect 101382 -1542 118826 -1306
rect 119062 -1542 119146 -1306
rect 119382 -1542 136826 -1306
rect 137062 -1542 137146 -1306
rect 137382 -1542 154826 -1306
rect 155062 -1542 155146 -1306
rect 155382 -1542 172826 -1306
rect 173062 -1542 173146 -1306
rect 173382 -1542 190826 -1306
rect 191062 -1542 191146 -1306
rect 191382 -1542 208826 -1306
rect 209062 -1542 209146 -1306
rect 209382 -1542 226826 -1306
rect 227062 -1542 227146 -1306
rect 227382 -1542 244826 -1306
rect 245062 -1542 245146 -1306
rect 245382 -1542 262826 -1306
rect 263062 -1542 263146 -1306
rect 263382 -1542 280826 -1306
rect 281062 -1542 281146 -1306
rect 281382 -1542 298826 -1306
rect 299062 -1542 299146 -1306
rect 299382 -1542 316826 -1306
rect 317062 -1542 317146 -1306
rect 317382 -1542 334826 -1306
rect 335062 -1542 335146 -1306
rect 335382 -1542 352826 -1306
rect 353062 -1542 353146 -1306
rect 353382 -1542 370826 -1306
rect 371062 -1542 371146 -1306
rect 371382 -1542 388826 -1306
rect 389062 -1542 389146 -1306
rect 389382 -1542 406826 -1306
rect 407062 -1542 407146 -1306
rect 407382 -1542 424826 -1306
rect 425062 -1542 425146 -1306
rect 425382 -1542 442826 -1306
rect 443062 -1542 443146 -1306
rect 443382 -1542 460826 -1306
rect 461062 -1542 461146 -1306
rect 461382 -1542 478826 -1306
rect 479062 -1542 479146 -1306
rect 479382 -1542 496826 -1306
rect 497062 -1542 497146 -1306
rect 497382 -1542 514826 -1306
rect 515062 -1542 515146 -1306
rect 515382 -1542 532826 -1306
rect 533062 -1542 533146 -1306
rect 533382 -1542 550826 -1306
rect 551062 -1542 551146 -1306
rect 551382 -1542 568826 -1306
rect 569062 -1542 569146 -1306
rect 569382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 10826 -1626
rect 11062 -1862 11146 -1626
rect 11382 -1862 28826 -1626
rect 29062 -1862 29146 -1626
rect 29382 -1862 46826 -1626
rect 47062 -1862 47146 -1626
rect 47382 -1862 64826 -1626
rect 65062 -1862 65146 -1626
rect 65382 -1862 82826 -1626
rect 83062 -1862 83146 -1626
rect 83382 -1862 100826 -1626
rect 101062 -1862 101146 -1626
rect 101382 -1862 118826 -1626
rect 119062 -1862 119146 -1626
rect 119382 -1862 136826 -1626
rect 137062 -1862 137146 -1626
rect 137382 -1862 154826 -1626
rect 155062 -1862 155146 -1626
rect 155382 -1862 172826 -1626
rect 173062 -1862 173146 -1626
rect 173382 -1862 190826 -1626
rect 191062 -1862 191146 -1626
rect 191382 -1862 208826 -1626
rect 209062 -1862 209146 -1626
rect 209382 -1862 226826 -1626
rect 227062 -1862 227146 -1626
rect 227382 -1862 244826 -1626
rect 245062 -1862 245146 -1626
rect 245382 -1862 262826 -1626
rect 263062 -1862 263146 -1626
rect 263382 -1862 280826 -1626
rect 281062 -1862 281146 -1626
rect 281382 -1862 298826 -1626
rect 299062 -1862 299146 -1626
rect 299382 -1862 316826 -1626
rect 317062 -1862 317146 -1626
rect 317382 -1862 334826 -1626
rect 335062 -1862 335146 -1626
rect 335382 -1862 352826 -1626
rect 353062 -1862 353146 -1626
rect 353382 -1862 370826 -1626
rect 371062 -1862 371146 -1626
rect 371382 -1862 388826 -1626
rect 389062 -1862 389146 -1626
rect 389382 -1862 406826 -1626
rect 407062 -1862 407146 -1626
rect 407382 -1862 424826 -1626
rect 425062 -1862 425146 -1626
rect 425382 -1862 442826 -1626
rect 443062 -1862 443146 -1626
rect 443382 -1862 460826 -1626
rect 461062 -1862 461146 -1626
rect 461382 -1862 478826 -1626
rect 479062 -1862 479146 -1626
rect 479382 -1862 496826 -1626
rect 497062 -1862 497146 -1626
rect 497382 -1862 514826 -1626
rect 515062 -1862 515146 -1626
rect 515382 -1862 532826 -1626
rect 533062 -1862 533146 -1626
rect 533382 -1862 550826 -1626
rect 551062 -1862 551146 -1626
rect 551382 -1862 568826 -1626
rect 569062 -1862 569146 -1626
rect 569382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
use scan_wrapper_lesson_1  instance_0
timestamp 0
transform 1 0 16000 0 1 16000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_1
timestamp 0
transform 1 0 43000 0 1 16000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_2
timestamp 0
transform 1 0 70000 0 1 16000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_3
timestamp 0
transform 1 0 97000 0 1 16000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_4
timestamp 0
transform 1 0 124000 0 1 16000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_5
timestamp 0
transform 1 0 151000 0 1 16000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_6
timestamp 0
transform 1 0 178000 0 1 16000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_7
timestamp 0
transform 1 0 205000 0 1 16000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_8
timestamp 0
transform 1 0 232000 0 1 16000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_9
timestamp 0
transform 1 0 259000 0 1 16000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_10
timestamp 0
transform 1 0 286000 0 1 16000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_11
timestamp 0
transform 1 0 313000 0 1 16000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_12
timestamp 0
transform 1 0 340000 0 1 16000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_13
timestamp 0
transform 1 0 367000 0 1 16000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_14
timestamp 0
transform 1 0 394000 0 1 16000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_15
timestamp 0
transform 1 0 421000 0 1 16000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_16
timestamp 0
transform 1 0 448000 0 1 16000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_17
timestamp 0
transform 1 0 475000 0 1 16000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_18
timestamp 0
transform 1 0 502000 0 1 16000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_19
timestamp 0
transform 1 0 529000 0 1 16000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_20
timestamp 0
transform 1 0 16000 0 1 43000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_21
timestamp 0
transform 1 0 43000 0 1 43000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_22
timestamp 0
transform 1 0 70000 0 1 43000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_23
timestamp 0
transform 1 0 97000 0 1 43000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_24
timestamp 0
transform 1 0 124000 0 1 43000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_25
timestamp 0
transform 1 0 151000 0 1 43000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_26
timestamp 0
transform 1 0 178000 0 1 43000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_27
timestamp 0
transform 1 0 205000 0 1 43000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_28
timestamp 0
transform 1 0 232000 0 1 43000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_29
timestamp 0
transform 1 0 259000 0 1 43000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_30
timestamp 0
transform 1 0 286000 0 1 43000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_31
timestamp 0
transform 1 0 313000 0 1 43000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_32
timestamp 0
transform 1 0 340000 0 1 43000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_33
timestamp 0
transform 1 0 367000 0 1 43000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_34
timestamp 0
transform 1 0 394000 0 1 43000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_35
timestamp 0
transform 1 0 421000 0 1 43000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_36
timestamp 0
transform 1 0 448000 0 1 43000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_37
timestamp 0
transform 1 0 475000 0 1 43000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_38
timestamp 0
transform 1 0 502000 0 1 43000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_39
timestamp 0
transform 1 0 529000 0 1 43000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_40
timestamp 0
transform 1 0 16000 0 1 70000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_41
timestamp 0
transform 1 0 43000 0 1 70000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_42
timestamp 0
transform 1 0 70000 0 1 70000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_43
timestamp 0
transform 1 0 97000 0 1 70000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_44
timestamp 0
transform 1 0 124000 0 1 70000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_45
timestamp 0
transform 1 0 151000 0 1 70000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_46
timestamp 0
transform 1 0 178000 0 1 70000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_47
timestamp 0
transform 1 0 205000 0 1 70000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_48
timestamp 0
transform 1 0 232000 0 1 70000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_49
timestamp 0
transform 1 0 259000 0 1 70000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_50
timestamp 0
transform 1 0 286000 0 1 70000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_51
timestamp 0
transform 1 0 313000 0 1 70000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_52
timestamp 0
transform 1 0 340000 0 1 70000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_53
timestamp 0
transform 1 0 367000 0 1 70000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_54
timestamp 0
transform 1 0 394000 0 1 70000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_55
timestamp 0
transform 1 0 421000 0 1 70000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_56
timestamp 0
transform 1 0 448000 0 1 70000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_57
timestamp 0
transform 1 0 475000 0 1 70000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_58
timestamp 0
transform 1 0 502000 0 1 70000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_59
timestamp 0
transform 1 0 529000 0 1 70000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_60
timestamp 0
transform 1 0 16000 0 1 97000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_61
timestamp 0
transform 1 0 43000 0 1 97000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_62
timestamp 0
transform 1 0 70000 0 1 97000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_63
timestamp 0
transform 1 0 97000 0 1 97000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_64
timestamp 0
transform 1 0 124000 0 1 97000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_65
timestamp 0
transform 1 0 151000 0 1 97000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_66
timestamp 0
transform 1 0 178000 0 1 97000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_67
timestamp 0
transform 1 0 205000 0 1 97000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_68
timestamp 0
transform 1 0 232000 0 1 97000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_69
timestamp 0
transform 1 0 259000 0 1 97000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_70
timestamp 0
transform 1 0 286000 0 1 97000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_71
timestamp 0
transform 1 0 313000 0 1 97000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_72
timestamp 0
transform 1 0 340000 0 1 97000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_73
timestamp 0
transform 1 0 367000 0 1 97000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_74
timestamp 0
transform 1 0 394000 0 1 97000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_75
timestamp 0
transform 1 0 421000 0 1 97000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_76
timestamp 0
transform 1 0 448000 0 1 97000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_77
timestamp 0
transform 1 0 475000 0 1 97000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_78
timestamp 0
transform 1 0 502000 0 1 97000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_79
timestamp 0
transform 1 0 529000 0 1 97000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_80
timestamp 0
transform 1 0 16000 0 1 124000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_81
timestamp 0
transform 1 0 43000 0 1 124000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_82
timestamp 0
transform 1 0 70000 0 1 124000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_83
timestamp 0
transform 1 0 97000 0 1 124000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_84
timestamp 0
transform 1 0 124000 0 1 124000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_85
timestamp 0
transform 1 0 151000 0 1 124000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_86
timestamp 0
transform 1 0 178000 0 1 124000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_87
timestamp 0
transform 1 0 205000 0 1 124000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_88
timestamp 0
transform 1 0 232000 0 1 124000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_89
timestamp 0
transform 1 0 259000 0 1 124000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_90
timestamp 0
transform 1 0 286000 0 1 124000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_91
timestamp 0
transform 1 0 313000 0 1 124000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_92
timestamp 0
transform 1 0 340000 0 1 124000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_93
timestamp 0
transform 1 0 367000 0 1 124000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_94
timestamp 0
transform 1 0 394000 0 1 124000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_95
timestamp 0
transform 1 0 421000 0 1 124000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_96
timestamp 0
transform 1 0 448000 0 1 124000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_97
timestamp 0
transform 1 0 475000 0 1 124000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_98
timestamp 0
transform 1 0 502000 0 1 124000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_99
timestamp 0
transform 1 0 529000 0 1 124000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_100
timestamp 0
transform 1 0 16000 0 1 151000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_101
timestamp 0
transform 1 0 43000 0 1 151000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_102
timestamp 0
transform 1 0 70000 0 1 151000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_103
timestamp 0
transform 1 0 97000 0 1 151000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_104
timestamp 0
transform 1 0 124000 0 1 151000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_105
timestamp 0
transform 1 0 151000 0 1 151000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_106
timestamp 0
transform 1 0 178000 0 1 151000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_107
timestamp 0
transform 1 0 205000 0 1 151000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_108
timestamp 0
transform 1 0 232000 0 1 151000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_109
timestamp 0
transform 1 0 259000 0 1 151000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_110
timestamp 0
transform 1 0 286000 0 1 151000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_111
timestamp 0
transform 1 0 313000 0 1 151000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_112
timestamp 0
transform 1 0 340000 0 1 151000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_113
timestamp 0
transform 1 0 367000 0 1 151000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_114
timestamp 0
transform 1 0 394000 0 1 151000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_115
timestamp 0
transform 1 0 421000 0 1 151000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_116
timestamp 0
transform 1 0 448000 0 1 151000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_117
timestamp 0
transform 1 0 475000 0 1 151000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_118
timestamp 0
transform 1 0 502000 0 1 151000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_119
timestamp 0
transform 1 0 529000 0 1 151000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_120
timestamp 0
transform 1 0 16000 0 1 178000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_121
timestamp 0
transform 1 0 43000 0 1 178000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_122
timestamp 0
transform 1 0 70000 0 1 178000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_123
timestamp 0
transform 1 0 97000 0 1 178000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_124
timestamp 0
transform 1 0 124000 0 1 178000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_125
timestamp 0
transform 1 0 151000 0 1 178000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_126
timestamp 0
transform 1 0 178000 0 1 178000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_127
timestamp 0
transform 1 0 205000 0 1 178000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_128
timestamp 0
transform 1 0 232000 0 1 178000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_129
timestamp 0
transform 1 0 259000 0 1 178000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_130
timestamp 0
transform 1 0 286000 0 1 178000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_131
timestamp 0
transform 1 0 313000 0 1 178000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_132
timestamp 0
transform 1 0 340000 0 1 178000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_133
timestamp 0
transform 1 0 367000 0 1 178000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_134
timestamp 0
transform 1 0 394000 0 1 178000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_135
timestamp 0
transform 1 0 421000 0 1 178000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_136
timestamp 0
transform 1 0 448000 0 1 178000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_137
timestamp 0
transform 1 0 475000 0 1 178000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_138
timestamp 0
transform 1 0 502000 0 1 178000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_139
timestamp 0
transform 1 0 529000 0 1 178000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_140
timestamp 0
transform 1 0 16000 0 1 205000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_141
timestamp 0
transform 1 0 43000 0 1 205000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_142
timestamp 0
transform 1 0 70000 0 1 205000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_143
timestamp 0
transform 1 0 97000 0 1 205000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_144
timestamp 0
transform 1 0 124000 0 1 205000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_145
timestamp 0
transform 1 0 151000 0 1 205000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_146
timestamp 0
transform 1 0 178000 0 1 205000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_147
timestamp 0
transform 1 0 205000 0 1 205000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_148
timestamp 0
transform 1 0 232000 0 1 205000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_149
timestamp 0
transform 1 0 259000 0 1 205000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_150
timestamp 0
transform 1 0 286000 0 1 205000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_151
timestamp 0
transform 1 0 313000 0 1 205000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_152
timestamp 0
transform 1 0 340000 0 1 205000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_153
timestamp 0
transform 1 0 367000 0 1 205000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_154
timestamp 0
transform 1 0 394000 0 1 205000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_155
timestamp 0
transform 1 0 421000 0 1 205000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_156
timestamp 0
transform 1 0 448000 0 1 205000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_157
timestamp 0
transform 1 0 475000 0 1 205000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_158
timestamp 0
transform 1 0 502000 0 1 205000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_159
timestamp 0
transform 1 0 529000 0 1 205000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_160
timestamp 0
transform 1 0 16000 0 1 232000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_161
timestamp 0
transform 1 0 43000 0 1 232000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_162
timestamp 0
transform 1 0 70000 0 1 232000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_163
timestamp 0
transform 1 0 97000 0 1 232000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_164
timestamp 0
transform 1 0 124000 0 1 232000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_165
timestamp 0
transform 1 0 151000 0 1 232000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_166
timestamp 0
transform 1 0 178000 0 1 232000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_167
timestamp 0
transform 1 0 205000 0 1 232000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_168
timestamp 0
transform 1 0 232000 0 1 232000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_169
timestamp 0
transform 1 0 259000 0 1 232000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_170
timestamp 0
transform 1 0 286000 0 1 232000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_171
timestamp 0
transform 1 0 313000 0 1 232000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_172
timestamp 0
transform 1 0 340000 0 1 232000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_173
timestamp 0
transform 1 0 367000 0 1 232000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_174
timestamp 0
transform 1 0 394000 0 1 232000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_175
timestamp 0
transform 1 0 421000 0 1 232000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_176
timestamp 0
transform 1 0 448000 0 1 232000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_177
timestamp 0
transform 1 0 475000 0 1 232000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_178
timestamp 0
transform 1 0 502000 0 1 232000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_179
timestamp 0
transform 1 0 529000 0 1 232000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_180
timestamp 0
transform 1 0 16000 0 1 259000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_181
timestamp 0
transform 1 0 43000 0 1 259000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_182
timestamp 0
transform 1 0 70000 0 1 259000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_183
timestamp 0
transform 1 0 97000 0 1 259000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_184
timestamp 0
transform 1 0 124000 0 1 259000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_185
timestamp 0
transform 1 0 151000 0 1 259000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_186
timestamp 0
transform 1 0 178000 0 1 259000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_187
timestamp 0
transform 1 0 205000 0 1 259000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_188
timestamp 0
transform 1 0 232000 0 1 259000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_189
timestamp 0
transform 1 0 259000 0 1 259000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_190
timestamp 0
transform 1 0 286000 0 1 259000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_191
timestamp 0
transform 1 0 313000 0 1 259000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_192
timestamp 0
transform 1 0 340000 0 1 259000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_193
timestamp 0
transform 1 0 367000 0 1 259000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_194
timestamp 0
transform 1 0 394000 0 1 259000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_195
timestamp 0
transform 1 0 421000 0 1 259000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_196
timestamp 0
transform 1 0 448000 0 1 259000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_197
timestamp 0
transform 1 0 475000 0 1 259000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_198
timestamp 0
transform 1 0 502000 0 1 259000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_199
timestamp 0
transform 1 0 529000 0 1 259000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_200
timestamp 0
transform 1 0 16000 0 1 286000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_201
timestamp 0
transform 1 0 43000 0 1 286000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_202
timestamp 0
transform 1 0 70000 0 1 286000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_203
timestamp 0
transform 1 0 97000 0 1 286000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_204
timestamp 0
transform 1 0 124000 0 1 286000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_205
timestamp 0
transform 1 0 151000 0 1 286000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_206
timestamp 0
transform 1 0 178000 0 1 286000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_207
timestamp 0
transform 1 0 205000 0 1 286000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_208
timestamp 0
transform 1 0 232000 0 1 286000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_209
timestamp 0
transform 1 0 259000 0 1 286000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_210
timestamp 0
transform 1 0 286000 0 1 286000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_211
timestamp 0
transform 1 0 313000 0 1 286000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_212
timestamp 0
transform 1 0 340000 0 1 286000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_213
timestamp 0
transform 1 0 367000 0 1 286000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_214
timestamp 0
transform 1 0 394000 0 1 286000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_215
timestamp 0
transform 1 0 421000 0 1 286000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_216
timestamp 0
transform 1 0 448000 0 1 286000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_217
timestamp 0
transform 1 0 475000 0 1 286000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_218
timestamp 0
transform 1 0 502000 0 1 286000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_219
timestamp 0
transform 1 0 529000 0 1 286000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_220
timestamp 0
transform 1 0 16000 0 1 313000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_221
timestamp 0
transform 1 0 43000 0 1 313000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_222
timestamp 0
transform 1 0 70000 0 1 313000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_223
timestamp 0
transform 1 0 97000 0 1 313000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_224
timestamp 0
transform 1 0 124000 0 1 313000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_225
timestamp 0
transform 1 0 151000 0 1 313000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_226
timestamp 0
transform 1 0 178000 0 1 313000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_227
timestamp 0
transform 1 0 205000 0 1 313000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_228
timestamp 0
transform 1 0 232000 0 1 313000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_229
timestamp 0
transform 1 0 259000 0 1 313000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_230
timestamp 0
transform 1 0 286000 0 1 313000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_231
timestamp 0
transform 1 0 313000 0 1 313000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_232
timestamp 0
transform 1 0 340000 0 1 313000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_233
timestamp 0
transform 1 0 367000 0 1 313000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_234
timestamp 0
transform 1 0 394000 0 1 313000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_235
timestamp 0
transform 1 0 421000 0 1 313000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_236
timestamp 0
transform 1 0 448000 0 1 313000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_237
timestamp 0
transform 1 0 475000 0 1 313000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_238
timestamp 0
transform 1 0 502000 0 1 313000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_239
timestamp 0
transform 1 0 529000 0 1 313000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_240
timestamp 0
transform 1 0 16000 0 1 340000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_241
timestamp 0
transform 1 0 43000 0 1 340000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_242
timestamp 0
transform 1 0 70000 0 1 340000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_243
timestamp 0
transform 1 0 97000 0 1 340000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_244
timestamp 0
transform 1 0 124000 0 1 340000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_245
timestamp 0
transform 1 0 151000 0 1 340000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_246
timestamp 0
transform 1 0 178000 0 1 340000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_247
timestamp 0
transform 1 0 205000 0 1 340000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_248
timestamp 0
transform 1 0 232000 0 1 340000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_249
timestamp 0
transform 1 0 259000 0 1 340000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_250
timestamp 0
transform 1 0 286000 0 1 340000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_251
timestamp 0
transform 1 0 313000 0 1 340000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_252
timestamp 0
transform 1 0 340000 0 1 340000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_253
timestamp 0
transform 1 0 367000 0 1 340000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_254
timestamp 0
transform 1 0 394000 0 1 340000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_255
timestamp 0
transform 1 0 421000 0 1 340000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_256
timestamp 0
transform 1 0 448000 0 1 340000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_257
timestamp 0
transform 1 0 475000 0 1 340000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_258
timestamp 0
transform 1 0 502000 0 1 340000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_259
timestamp 0
transform 1 0 529000 0 1 340000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_260
timestamp 0
transform 1 0 16000 0 1 367000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_261
timestamp 0
transform 1 0 43000 0 1 367000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_262
timestamp 0
transform 1 0 70000 0 1 367000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_263
timestamp 0
transform 1 0 97000 0 1 367000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_264
timestamp 0
transform 1 0 124000 0 1 367000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_265
timestamp 0
transform 1 0 151000 0 1 367000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_266
timestamp 0
transform 1 0 178000 0 1 367000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_267
timestamp 0
transform 1 0 205000 0 1 367000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_268
timestamp 0
transform 1 0 232000 0 1 367000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_269
timestamp 0
transform 1 0 259000 0 1 367000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_270
timestamp 0
transform 1 0 286000 0 1 367000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_271
timestamp 0
transform 1 0 313000 0 1 367000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_272
timestamp 0
transform 1 0 340000 0 1 367000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_273
timestamp 0
transform 1 0 367000 0 1 367000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_274
timestamp 0
transform 1 0 394000 0 1 367000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_275
timestamp 0
transform 1 0 421000 0 1 367000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_276
timestamp 0
transform 1 0 448000 0 1 367000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_277
timestamp 0
transform 1 0 475000 0 1 367000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_278
timestamp 0
transform 1 0 502000 0 1 367000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_279
timestamp 0
transform 1 0 529000 0 1 367000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_280
timestamp 0
transform 1 0 16000 0 1 394000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_281
timestamp 0
transform 1 0 43000 0 1 394000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_282
timestamp 0
transform 1 0 70000 0 1 394000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_283
timestamp 0
transform 1 0 97000 0 1 394000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_284
timestamp 0
transform 1 0 124000 0 1 394000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_285
timestamp 0
transform 1 0 151000 0 1 394000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_286
timestamp 0
transform 1 0 178000 0 1 394000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_287
timestamp 0
transform 1 0 205000 0 1 394000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_288
timestamp 0
transform 1 0 232000 0 1 394000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_289
timestamp 0
transform 1 0 259000 0 1 394000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_290
timestamp 0
transform 1 0 286000 0 1 394000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_291
timestamp 0
transform 1 0 313000 0 1 394000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_292
timestamp 0
transform 1 0 340000 0 1 394000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_293
timestamp 0
transform 1 0 367000 0 1 394000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_294
timestamp 0
transform 1 0 394000 0 1 394000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_295
timestamp 0
transform 1 0 421000 0 1 394000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_296
timestamp 0
transform 1 0 448000 0 1 394000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_297
timestamp 0
transform 1 0 475000 0 1 394000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_298
timestamp 0
transform 1 0 502000 0 1 394000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_299
timestamp 0
transform 1 0 529000 0 1 394000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_300
timestamp 0
transform 1 0 16000 0 1 421000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_301
timestamp 0
transform 1 0 43000 0 1 421000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_302
timestamp 0
transform 1 0 70000 0 1 421000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_303
timestamp 0
transform 1 0 97000 0 1 421000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_304
timestamp 0
transform 1 0 124000 0 1 421000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_305
timestamp 0
transform 1 0 151000 0 1 421000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_306
timestamp 0
transform 1 0 178000 0 1 421000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_307
timestamp 0
transform 1 0 205000 0 1 421000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_308
timestamp 0
transform 1 0 232000 0 1 421000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_309
timestamp 0
transform 1 0 259000 0 1 421000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_310
timestamp 0
transform 1 0 286000 0 1 421000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_311
timestamp 0
transform 1 0 313000 0 1 421000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_312
timestamp 0
transform 1 0 340000 0 1 421000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_313
timestamp 0
transform 1 0 367000 0 1 421000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_314
timestamp 0
transform 1 0 394000 0 1 421000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_315
timestamp 0
transform 1 0 421000 0 1 421000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_316
timestamp 0
transform 1 0 448000 0 1 421000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_317
timestamp 0
transform 1 0 475000 0 1 421000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_318
timestamp 0
transform 1 0 502000 0 1 421000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_319
timestamp 0
transform 1 0 529000 0 1 421000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_320
timestamp 0
transform 1 0 16000 0 1 448000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_321
timestamp 0
transform 1 0 43000 0 1 448000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_322
timestamp 0
transform 1 0 70000 0 1 448000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_323
timestamp 0
transform 1 0 97000 0 1 448000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_324
timestamp 0
transform 1 0 124000 0 1 448000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_325
timestamp 0
transform 1 0 151000 0 1 448000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_326
timestamp 0
transform 1 0 178000 0 1 448000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_327
timestamp 0
transform 1 0 205000 0 1 448000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_328
timestamp 0
transform 1 0 232000 0 1 448000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_329
timestamp 0
transform 1 0 259000 0 1 448000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_330
timestamp 0
transform 1 0 286000 0 1 448000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_331
timestamp 0
transform 1 0 313000 0 1 448000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_332
timestamp 0
transform 1 0 340000 0 1 448000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_333
timestamp 0
transform 1 0 367000 0 1 448000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_334
timestamp 0
transform 1 0 394000 0 1 448000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_335
timestamp 0
transform 1 0 421000 0 1 448000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_336
timestamp 0
transform 1 0 448000 0 1 448000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_337
timestamp 0
transform 1 0 475000 0 1 448000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_338
timestamp 0
transform 1 0 502000 0 1 448000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_339
timestamp 0
transform 1 0 529000 0 1 448000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_340
timestamp 0
transform 1 0 16000 0 1 475000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_341
timestamp 0
transform 1 0 43000 0 1 475000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_342
timestamp 0
transform 1 0 70000 0 1 475000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_343
timestamp 0
transform 1 0 97000 0 1 475000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_344
timestamp 0
transform 1 0 124000 0 1 475000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_345
timestamp 0
transform 1 0 151000 0 1 475000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_346
timestamp 0
transform 1 0 178000 0 1 475000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_347
timestamp 0
transform 1 0 205000 0 1 475000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_348
timestamp 0
transform 1 0 232000 0 1 475000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_349
timestamp 0
transform 1 0 259000 0 1 475000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_350
timestamp 0
transform 1 0 286000 0 1 475000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_351
timestamp 0
transform 1 0 313000 0 1 475000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_352
timestamp 0
transform 1 0 340000 0 1 475000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_353
timestamp 0
transform 1 0 367000 0 1 475000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_354
timestamp 0
transform 1 0 394000 0 1 475000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_355
timestamp 0
transform 1 0 421000 0 1 475000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_356
timestamp 0
transform 1 0 448000 0 1 475000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_357
timestamp 0
transform 1 0 475000 0 1 475000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_358
timestamp 0
transform 1 0 502000 0 1 475000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_359
timestamp 0
transform 1 0 529000 0 1 475000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_360
timestamp 0
transform 1 0 16000 0 1 502000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_361
timestamp 0
transform 1 0 43000 0 1 502000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_362
timestamp 0
transform 1 0 70000 0 1 502000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_363
timestamp 0
transform 1 0 97000 0 1 502000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_364
timestamp 0
transform 1 0 124000 0 1 502000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_365
timestamp 0
transform 1 0 151000 0 1 502000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_366
timestamp 0
transform 1 0 178000 0 1 502000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_367
timestamp 0
transform 1 0 205000 0 1 502000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_368
timestamp 0
transform 1 0 232000 0 1 502000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_369
timestamp 0
transform 1 0 259000 0 1 502000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_370
timestamp 0
transform 1 0 286000 0 1 502000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_371
timestamp 0
transform 1 0 313000 0 1 502000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_372
timestamp 0
transform 1 0 340000 0 1 502000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_373
timestamp 0
transform 1 0 367000 0 1 502000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_374
timestamp 0
transform 1 0 394000 0 1 502000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_375
timestamp 0
transform 1 0 421000 0 1 502000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_376
timestamp 0
transform 1 0 448000 0 1 502000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_377
timestamp 0
transform 1 0 475000 0 1 502000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_378
timestamp 0
transform 1 0 502000 0 1 502000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_379
timestamp 0
transform 1 0 529000 0 1 502000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_380
timestamp 0
transform 1 0 16000 0 1 529000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_381
timestamp 0
transform 1 0 43000 0 1 529000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_382
timestamp 0
transform 1 0 70000 0 1 529000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_383
timestamp 0
transform 1 0 97000 0 1 529000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_384
timestamp 0
transform 1 0 124000 0 1 529000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_385
timestamp 0
transform 1 0 151000 0 1 529000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_386
timestamp 0
transform 1 0 178000 0 1 529000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_387
timestamp 0
transform 1 0 205000 0 1 529000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_388
timestamp 0
transform 1 0 232000 0 1 529000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_389
timestamp 0
transform 1 0 259000 0 1 529000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_390
timestamp 0
transform 1 0 286000 0 1 529000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_391
timestamp 0
transform 1 0 313000 0 1 529000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_392
timestamp 0
transform 1 0 340000 0 1 529000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_393
timestamp 0
transform 1 0 367000 0 1 529000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_394
timestamp 0
transform 1 0 394000 0 1 529000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_395
timestamp 0
transform 1 0 421000 0 1 529000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_396
timestamp 0
transform 1 0 448000 0 1 529000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_397
timestamp 0
transform 1 0 475000 0 1 529000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_398
timestamp 0
transform 1 0 502000 0 1 529000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_399
timestamp 0
transform 1 0 529000 0 1 529000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_400
timestamp 0
transform 1 0 16000 0 1 556000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_401
timestamp 0
transform 1 0 43000 0 1 556000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_402
timestamp 0
transform 1 0 70000 0 1 556000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_403
timestamp 0
transform 1 0 97000 0 1 556000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_404
timestamp 0
transform 1 0 124000 0 1 556000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_405
timestamp 0
transform 1 0 151000 0 1 556000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_406
timestamp 0
transform 1 0 178000 0 1 556000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_407
timestamp 0
transform 1 0 205000 0 1 556000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_408
timestamp 0
transform 1 0 232000 0 1 556000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_409
timestamp 0
transform 1 0 259000 0 1 556000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_410
timestamp 0
transform 1 0 286000 0 1 556000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_411
timestamp 0
transform 1 0 313000 0 1 556000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_412
timestamp 0
transform 1 0 340000 0 1 556000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_413
timestamp 0
transform 1 0 367000 0 1 556000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_414
timestamp 0
transform 1 0 394000 0 1 556000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_415
timestamp 0
transform 1 0 421000 0 1 556000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_416
timestamp 0
transform 1 0 448000 0 1 556000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_417
timestamp 0
transform 1 0 475000 0 1 556000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_418
timestamp 0
transform 1 0 502000 0 1 556000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_419
timestamp 0
transform 1 0 529000 0 1 556000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_420
timestamp 0
transform 1 0 16000 0 1 583000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_421
timestamp 0
transform 1 0 43000 0 1 583000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_422
timestamp 0
transform 1 0 70000 0 1 583000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_423
timestamp 0
transform 1 0 97000 0 1 583000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_424
timestamp 0
transform 1 0 124000 0 1 583000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_425
timestamp 0
transform 1 0 151000 0 1 583000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_426
timestamp 0
transform 1 0 178000 0 1 583000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_427
timestamp 0
transform 1 0 205000 0 1 583000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_428
timestamp 0
transform 1 0 232000 0 1 583000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_429
timestamp 0
transform 1 0 259000 0 1 583000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_430
timestamp 0
transform 1 0 286000 0 1 583000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_431
timestamp 0
transform 1 0 313000 0 1 583000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_432
timestamp 0
transform 1 0 340000 0 1 583000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_433
timestamp 0
transform 1 0 367000 0 1 583000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_434
timestamp 0
transform 1 0 394000 0 1 583000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_435
timestamp 0
transform 1 0 421000 0 1 583000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_436
timestamp 0
transform 1 0 448000 0 1 583000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_437
timestamp 0
transform 1 0 475000 0 1 583000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_438
timestamp 0
transform 1 0 502000 0 1 583000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_439
timestamp 0
transform 1 0 529000 0 1 583000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_440
timestamp 0
transform 1 0 16000 0 1 610000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_441
timestamp 0
transform 1 0 43000 0 1 610000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_442
timestamp 0
transform 1 0 70000 0 1 610000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_443
timestamp 0
transform 1 0 97000 0 1 610000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_444
timestamp 0
transform 1 0 124000 0 1 610000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_445
timestamp 0
transform 1 0 151000 0 1 610000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_446
timestamp 0
transform 1 0 178000 0 1 610000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_447
timestamp 0
transform 1 0 205000 0 1 610000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_448
timestamp 0
transform 1 0 232000 0 1 610000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_449
timestamp 0
transform 1 0 259000 0 1 610000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_450
timestamp 0
transform 1 0 286000 0 1 610000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_451
timestamp 0
transform 1 0 313000 0 1 610000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_452
timestamp 0
transform 1 0 340000 0 1 610000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_453
timestamp 0
transform 1 0 367000 0 1 610000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_454
timestamp 0
transform 1 0 394000 0 1 610000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_455
timestamp 0
transform 1 0 421000 0 1 610000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_456
timestamp 0
transform 1 0 448000 0 1 610000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_457
timestamp 0
transform 1 0 475000 0 1 610000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_458
timestamp 0
transform 1 0 502000 0 1 610000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_459
timestamp 0
transform 1 0 529000 0 1 610000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_460
timestamp 0
transform 1 0 16000 0 1 637000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_461
timestamp 0
transform 1 0 43000 0 1 637000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_462
timestamp 0
transform 1 0 70000 0 1 637000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_463
timestamp 0
transform 1 0 97000 0 1 637000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_464
timestamp 0
transform 1 0 124000 0 1 637000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_465
timestamp 0
transform 1 0 151000 0 1 637000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_466
timestamp 0
transform 1 0 178000 0 1 637000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_467
timestamp 0
transform 1 0 205000 0 1 637000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_468
timestamp 0
transform 1 0 232000 0 1 637000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_469
timestamp 0
transform 1 0 259000 0 1 637000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_470
timestamp 0
transform 1 0 286000 0 1 637000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_471
timestamp 0
transform 1 0 313000 0 1 637000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_472
timestamp 0
transform 1 0 340000 0 1 637000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_473
timestamp 0
transform 1 0 367000 0 1 637000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_474
timestamp 0
transform 1 0 394000 0 1 637000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_475
timestamp 0
transform 1 0 421000 0 1 637000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_476
timestamp 0
transform 1 0 448000 0 1 637000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_477
timestamp 0
transform 1 0 475000 0 1 637000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_478
timestamp 0
transform 1 0 502000 0 1 637000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_479
timestamp 0
transform 1 0 529000 0 1 637000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_480
timestamp 0
transform 1 0 16000 0 1 664000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_481
timestamp 0
transform 1 0 43000 0 1 664000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_482
timestamp 0
transform 1 0 70000 0 1 664000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_483
timestamp 0
transform 1 0 97000 0 1 664000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_484
timestamp 0
transform 1 0 124000 0 1 664000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_485
timestamp 0
transform 1 0 151000 0 1 664000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_486
timestamp 0
transform 1 0 178000 0 1 664000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_487
timestamp 0
transform 1 0 205000 0 1 664000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_488
timestamp 0
transform 1 0 232000 0 1 664000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_489
timestamp 0
transform 1 0 259000 0 1 664000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_490
timestamp 0
transform 1 0 286000 0 1 664000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_491
timestamp 0
transform 1 0 313000 0 1 664000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_492
timestamp 0
transform 1 0 340000 0 1 664000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_493
timestamp 0
transform 1 0 367000 0 1 664000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_494
timestamp 0
transform 1 0 394000 0 1 664000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_495
timestamp 0
transform 1 0 421000 0 1 664000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_496
timestamp 0
transform 1 0 448000 0 1 664000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_497
timestamp 0
transform 1 0 475000 0 1 664000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_498
timestamp 0
transform 1 0 502000 0 1 664000
box -10 0 20000 20000
use scan_wrapper_lesson_1  instance_499
timestamp 0
transform 1 0 529000 0 1 664000
box -10 0 20000 20000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 20866 586890 21486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 56866 586890 57486 6 vccd1
port 531 nsew power input
rlabel metal5 s 19794 66806 542414 67426 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 92866 586890 93486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s 19794 120806 542414 121426 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 128866 586890 129486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 164866 586890 165486 6 vccd1
port 531 nsew power input
rlabel metal5 s 19794 174806 542414 175426 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 200866 586890 201486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s 19794 228806 542414 229426 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 236866 586890 237486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 272866 586890 273486 6 vccd1
port 531 nsew power input
rlabel metal5 s 19794 282806 542414 283426 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 308866 586890 309486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s 19794 336806 542414 337426 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 344866 586890 345486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 380866 586890 381486 6 vccd1
port 531 nsew power input
rlabel metal5 s 19794 390806 542414 391426 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 416866 586890 417486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s 19794 444806 542414 445426 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 452866 586890 453486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 488866 586890 489486 6 vccd1
port 531 nsew power input
rlabel metal5 s 19794 498806 542414 499426 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 524866 586890 525486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s 19794 552806 542414 553426 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 560866 586890 561486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 596866 586890 597486 6 vccd1
port 531 nsew power input
rlabel metal5 s 19794 606806 542414 607426 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 632866 586890 633486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s 19794 660806 542414 661426 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 668866 586890 669486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 19794 -1894 20414 14000 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 14000 6 vccd1
port 531 nsew power input
rlabel metal4 s 55794 -1894 56414 14000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 14000 6 vccd1
port 531 nsew power input
rlabel metal4 s 91794 -1894 92414 14000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 14000 6 vccd1
port 531 nsew power input
rlabel metal4 s 127794 -1894 128414 14000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 14000 6 vccd1
port 531 nsew power input
rlabel metal4 s 163794 -1894 164414 14000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 14000 6 vccd1
port 531 nsew power input
rlabel metal4 s 199794 -1894 200414 14000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 14000 6 vccd1
port 531 nsew power input
rlabel metal4 s 235794 -1894 236414 14000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 14000 6 vccd1
port 531 nsew power input
rlabel metal4 s 271794 -1894 272414 14000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 14000 6 vccd1
port 531 nsew power input
rlabel metal4 s 307794 -1894 308414 14000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 14000 6 vccd1
port 531 nsew power input
rlabel metal4 s 343794 -1894 344414 14000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 14000 6 vccd1
port 531 nsew power input
rlabel metal4 s 379794 -1894 380414 14000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 14000 6 vccd1
port 531 nsew power input
rlabel metal4 s 415794 -1894 416414 14000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 14000 6 vccd1
port 531 nsew power input
rlabel metal4 s 451794 -1894 452414 14000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 14000 6 vccd1
port 531 nsew power input
rlabel metal4 s 487794 -1894 488414 14000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 14000 6 vccd1
port 531 nsew power input
rlabel metal4 s 523794 -1894 524414 14000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 14000 6 vccd1
port 531 nsew power input
rlabel metal4 s 19794 38000 20414 41000 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 38000 38414 41000 6 vccd1
port 531 nsew power input
rlabel metal4 s 55794 38000 56414 41000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 38000 74414 41000 6 vccd1
port 531 nsew power input
rlabel metal4 s 91794 38000 92414 41000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 38000 110414 41000 6 vccd1
port 531 nsew power input
rlabel metal4 s 127794 38000 128414 41000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 38000 146414 41000 6 vccd1
port 531 nsew power input
rlabel metal4 s 163794 38000 164414 41000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 38000 182414 41000 6 vccd1
port 531 nsew power input
rlabel metal4 s 199794 38000 200414 41000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 38000 218414 41000 6 vccd1
port 531 nsew power input
rlabel metal4 s 235794 38000 236414 41000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 38000 254414 41000 6 vccd1
port 531 nsew power input
rlabel metal4 s 271794 38000 272414 41000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 38000 290414 41000 6 vccd1
port 531 nsew power input
rlabel metal4 s 307794 38000 308414 41000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 38000 326414 41000 6 vccd1
port 531 nsew power input
rlabel metal4 s 343794 38000 344414 41000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 38000 362414 41000 6 vccd1
port 531 nsew power input
rlabel metal4 s 379794 38000 380414 41000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 38000 398414 41000 6 vccd1
port 531 nsew power input
rlabel metal4 s 415794 38000 416414 41000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 38000 434414 41000 6 vccd1
port 531 nsew power input
rlabel metal4 s 451794 38000 452414 41000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 38000 470414 41000 6 vccd1
port 531 nsew power input
rlabel metal4 s 487794 38000 488414 41000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 38000 506414 41000 6 vccd1
port 531 nsew power input
rlabel metal4 s 523794 38000 524414 41000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 38000 542414 41000 6 vccd1
port 531 nsew power input
rlabel metal4 s 19794 65000 20414 68000 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 65000 38414 68000 6 vccd1
port 531 nsew power input
rlabel metal4 s 55794 65000 56414 68000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 65000 74414 68000 6 vccd1
port 531 nsew power input
rlabel metal4 s 91794 65000 92414 68000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 65000 110414 68000 6 vccd1
port 531 nsew power input
rlabel metal4 s 127794 65000 128414 68000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 65000 146414 68000 6 vccd1
port 531 nsew power input
rlabel metal4 s 163794 65000 164414 68000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 65000 182414 68000 6 vccd1
port 531 nsew power input
rlabel metal4 s 199794 65000 200414 68000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 65000 218414 68000 6 vccd1
port 531 nsew power input
rlabel metal4 s 235794 65000 236414 68000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 65000 254414 68000 6 vccd1
port 531 nsew power input
rlabel metal4 s 271794 65000 272414 68000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 65000 290414 68000 6 vccd1
port 531 nsew power input
rlabel metal4 s 307794 65000 308414 68000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 65000 326414 68000 6 vccd1
port 531 nsew power input
rlabel metal4 s 343794 65000 344414 68000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 65000 362414 68000 6 vccd1
port 531 nsew power input
rlabel metal4 s 379794 65000 380414 68000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 65000 398414 68000 6 vccd1
port 531 nsew power input
rlabel metal4 s 415794 65000 416414 68000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 65000 434414 68000 6 vccd1
port 531 nsew power input
rlabel metal4 s 451794 65000 452414 68000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 65000 470414 68000 6 vccd1
port 531 nsew power input
rlabel metal4 s 487794 65000 488414 68000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 65000 506414 68000 6 vccd1
port 531 nsew power input
rlabel metal4 s 523794 65000 524414 68000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 65000 542414 68000 6 vccd1
port 531 nsew power input
rlabel metal4 s 19794 92000 20414 95000 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 92000 38414 95000 6 vccd1
port 531 nsew power input
rlabel metal4 s 55794 92000 56414 95000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 92000 74414 95000 6 vccd1
port 531 nsew power input
rlabel metal4 s 91794 92000 92414 95000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 92000 110414 95000 6 vccd1
port 531 nsew power input
rlabel metal4 s 127794 92000 128414 95000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 92000 146414 95000 6 vccd1
port 531 nsew power input
rlabel metal4 s 163794 92000 164414 95000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 92000 182414 95000 6 vccd1
port 531 nsew power input
rlabel metal4 s 199794 92000 200414 95000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 92000 218414 95000 6 vccd1
port 531 nsew power input
rlabel metal4 s 235794 92000 236414 95000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 92000 254414 95000 6 vccd1
port 531 nsew power input
rlabel metal4 s 271794 92000 272414 95000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 92000 290414 95000 6 vccd1
port 531 nsew power input
rlabel metal4 s 307794 92000 308414 95000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 92000 326414 95000 6 vccd1
port 531 nsew power input
rlabel metal4 s 343794 92000 344414 95000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 92000 362414 95000 6 vccd1
port 531 nsew power input
rlabel metal4 s 379794 92000 380414 95000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 92000 398414 95000 6 vccd1
port 531 nsew power input
rlabel metal4 s 415794 92000 416414 95000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 92000 434414 95000 6 vccd1
port 531 nsew power input
rlabel metal4 s 451794 92000 452414 95000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 92000 470414 95000 6 vccd1
port 531 nsew power input
rlabel metal4 s 487794 92000 488414 95000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 92000 506414 95000 6 vccd1
port 531 nsew power input
rlabel metal4 s 523794 92000 524414 95000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 92000 542414 95000 6 vccd1
port 531 nsew power input
rlabel metal4 s 19794 119000 20414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 119000 38414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 55794 119000 56414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 119000 74414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 91794 119000 92414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 119000 110414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 127794 119000 128414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 119000 146414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 163794 119000 164414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 119000 182414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 199794 119000 200414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 119000 218414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 235794 119000 236414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 119000 254414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 271794 119000 272414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 119000 290414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 307794 119000 308414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 119000 326414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 343794 119000 344414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 119000 362414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 379794 119000 380414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 119000 398414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 415794 119000 416414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 119000 434414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 451794 119000 452414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 119000 470414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 487794 119000 488414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 119000 506414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 523794 119000 524414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 119000 542414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 19794 146000 20414 149000 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 146000 38414 149000 6 vccd1
port 531 nsew power input
rlabel metal4 s 55794 146000 56414 149000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 146000 74414 149000 6 vccd1
port 531 nsew power input
rlabel metal4 s 91794 146000 92414 149000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 146000 110414 149000 6 vccd1
port 531 nsew power input
rlabel metal4 s 127794 146000 128414 149000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 146000 146414 149000 6 vccd1
port 531 nsew power input
rlabel metal4 s 163794 146000 164414 149000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 146000 182414 149000 6 vccd1
port 531 nsew power input
rlabel metal4 s 199794 146000 200414 149000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 146000 218414 149000 6 vccd1
port 531 nsew power input
rlabel metal4 s 235794 146000 236414 149000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 146000 254414 149000 6 vccd1
port 531 nsew power input
rlabel metal4 s 271794 146000 272414 149000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 146000 290414 149000 6 vccd1
port 531 nsew power input
rlabel metal4 s 307794 146000 308414 149000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 146000 326414 149000 6 vccd1
port 531 nsew power input
rlabel metal4 s 343794 146000 344414 149000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 146000 362414 149000 6 vccd1
port 531 nsew power input
rlabel metal4 s 379794 146000 380414 149000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 146000 398414 149000 6 vccd1
port 531 nsew power input
rlabel metal4 s 415794 146000 416414 149000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 146000 434414 149000 6 vccd1
port 531 nsew power input
rlabel metal4 s 451794 146000 452414 149000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 146000 470414 149000 6 vccd1
port 531 nsew power input
rlabel metal4 s 487794 146000 488414 149000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 146000 506414 149000 6 vccd1
port 531 nsew power input
rlabel metal4 s 523794 146000 524414 149000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 146000 542414 149000 6 vccd1
port 531 nsew power input
rlabel metal4 s 19794 173000 20414 176000 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 173000 38414 176000 6 vccd1
port 531 nsew power input
rlabel metal4 s 55794 173000 56414 176000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 173000 74414 176000 6 vccd1
port 531 nsew power input
rlabel metal4 s 91794 173000 92414 176000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 173000 110414 176000 6 vccd1
port 531 nsew power input
rlabel metal4 s 127794 173000 128414 176000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 173000 146414 176000 6 vccd1
port 531 nsew power input
rlabel metal4 s 163794 173000 164414 176000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 173000 182414 176000 6 vccd1
port 531 nsew power input
rlabel metal4 s 199794 173000 200414 176000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 173000 218414 176000 6 vccd1
port 531 nsew power input
rlabel metal4 s 235794 173000 236414 176000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 173000 254414 176000 6 vccd1
port 531 nsew power input
rlabel metal4 s 271794 173000 272414 176000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 173000 290414 176000 6 vccd1
port 531 nsew power input
rlabel metal4 s 307794 173000 308414 176000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 173000 326414 176000 6 vccd1
port 531 nsew power input
rlabel metal4 s 343794 173000 344414 176000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 173000 362414 176000 6 vccd1
port 531 nsew power input
rlabel metal4 s 379794 173000 380414 176000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 173000 398414 176000 6 vccd1
port 531 nsew power input
rlabel metal4 s 415794 173000 416414 176000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 173000 434414 176000 6 vccd1
port 531 nsew power input
rlabel metal4 s 451794 173000 452414 176000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 173000 470414 176000 6 vccd1
port 531 nsew power input
rlabel metal4 s 487794 173000 488414 176000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 173000 506414 176000 6 vccd1
port 531 nsew power input
rlabel metal4 s 523794 173000 524414 176000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 173000 542414 176000 6 vccd1
port 531 nsew power input
rlabel metal4 s 19794 200000 20414 203000 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 200000 38414 203000 6 vccd1
port 531 nsew power input
rlabel metal4 s 55794 200000 56414 203000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 200000 74414 203000 6 vccd1
port 531 nsew power input
rlabel metal4 s 91794 200000 92414 203000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 200000 110414 203000 6 vccd1
port 531 nsew power input
rlabel metal4 s 127794 200000 128414 203000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 200000 146414 203000 6 vccd1
port 531 nsew power input
rlabel metal4 s 163794 200000 164414 203000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 200000 182414 203000 6 vccd1
port 531 nsew power input
rlabel metal4 s 199794 200000 200414 203000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 200000 218414 203000 6 vccd1
port 531 nsew power input
rlabel metal4 s 235794 200000 236414 203000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 200000 254414 203000 6 vccd1
port 531 nsew power input
rlabel metal4 s 271794 200000 272414 203000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 200000 290414 203000 6 vccd1
port 531 nsew power input
rlabel metal4 s 307794 200000 308414 203000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 200000 326414 203000 6 vccd1
port 531 nsew power input
rlabel metal4 s 343794 200000 344414 203000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 200000 362414 203000 6 vccd1
port 531 nsew power input
rlabel metal4 s 379794 200000 380414 203000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 200000 398414 203000 6 vccd1
port 531 nsew power input
rlabel metal4 s 415794 200000 416414 203000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 200000 434414 203000 6 vccd1
port 531 nsew power input
rlabel metal4 s 451794 200000 452414 203000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 200000 470414 203000 6 vccd1
port 531 nsew power input
rlabel metal4 s 487794 200000 488414 203000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 200000 506414 203000 6 vccd1
port 531 nsew power input
rlabel metal4 s 523794 200000 524414 203000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 200000 542414 203000 6 vccd1
port 531 nsew power input
rlabel metal4 s 19794 227000 20414 230000 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 227000 38414 230000 6 vccd1
port 531 nsew power input
rlabel metal4 s 55794 227000 56414 230000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 227000 74414 230000 6 vccd1
port 531 nsew power input
rlabel metal4 s 91794 227000 92414 230000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 227000 110414 230000 6 vccd1
port 531 nsew power input
rlabel metal4 s 127794 227000 128414 230000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 227000 146414 230000 6 vccd1
port 531 nsew power input
rlabel metal4 s 163794 227000 164414 230000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 227000 182414 230000 6 vccd1
port 531 nsew power input
rlabel metal4 s 199794 227000 200414 230000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 227000 218414 230000 6 vccd1
port 531 nsew power input
rlabel metal4 s 235794 227000 236414 230000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 227000 254414 230000 6 vccd1
port 531 nsew power input
rlabel metal4 s 271794 227000 272414 230000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 227000 290414 230000 6 vccd1
port 531 nsew power input
rlabel metal4 s 307794 227000 308414 230000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 227000 326414 230000 6 vccd1
port 531 nsew power input
rlabel metal4 s 343794 227000 344414 230000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 227000 362414 230000 6 vccd1
port 531 nsew power input
rlabel metal4 s 379794 227000 380414 230000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 227000 398414 230000 6 vccd1
port 531 nsew power input
rlabel metal4 s 415794 227000 416414 230000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 227000 434414 230000 6 vccd1
port 531 nsew power input
rlabel metal4 s 451794 227000 452414 230000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 227000 470414 230000 6 vccd1
port 531 nsew power input
rlabel metal4 s 487794 227000 488414 230000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 227000 506414 230000 6 vccd1
port 531 nsew power input
rlabel metal4 s 523794 227000 524414 230000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 227000 542414 230000 6 vccd1
port 531 nsew power input
rlabel metal4 s 19794 254000 20414 257000 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 254000 38414 257000 6 vccd1
port 531 nsew power input
rlabel metal4 s 55794 254000 56414 257000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 254000 74414 257000 6 vccd1
port 531 nsew power input
rlabel metal4 s 91794 254000 92414 257000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 254000 110414 257000 6 vccd1
port 531 nsew power input
rlabel metal4 s 127794 254000 128414 257000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 254000 146414 257000 6 vccd1
port 531 nsew power input
rlabel metal4 s 163794 254000 164414 257000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 254000 182414 257000 6 vccd1
port 531 nsew power input
rlabel metal4 s 199794 254000 200414 257000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 254000 218414 257000 6 vccd1
port 531 nsew power input
rlabel metal4 s 235794 254000 236414 257000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 254000 254414 257000 6 vccd1
port 531 nsew power input
rlabel metal4 s 271794 254000 272414 257000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 254000 290414 257000 6 vccd1
port 531 nsew power input
rlabel metal4 s 307794 254000 308414 257000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 254000 326414 257000 6 vccd1
port 531 nsew power input
rlabel metal4 s 343794 254000 344414 257000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 254000 362414 257000 6 vccd1
port 531 nsew power input
rlabel metal4 s 379794 254000 380414 257000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 254000 398414 257000 6 vccd1
port 531 nsew power input
rlabel metal4 s 415794 254000 416414 257000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 254000 434414 257000 6 vccd1
port 531 nsew power input
rlabel metal4 s 451794 254000 452414 257000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 254000 470414 257000 6 vccd1
port 531 nsew power input
rlabel metal4 s 487794 254000 488414 257000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 254000 506414 257000 6 vccd1
port 531 nsew power input
rlabel metal4 s 523794 254000 524414 257000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 254000 542414 257000 6 vccd1
port 531 nsew power input
rlabel metal4 s 19794 281000 20414 284000 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 281000 38414 284000 6 vccd1
port 531 nsew power input
rlabel metal4 s 55794 281000 56414 284000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 281000 74414 284000 6 vccd1
port 531 nsew power input
rlabel metal4 s 91794 281000 92414 284000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 281000 110414 284000 6 vccd1
port 531 nsew power input
rlabel metal4 s 127794 281000 128414 284000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 281000 146414 284000 6 vccd1
port 531 nsew power input
rlabel metal4 s 163794 281000 164414 284000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 281000 182414 284000 6 vccd1
port 531 nsew power input
rlabel metal4 s 199794 281000 200414 284000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 281000 218414 284000 6 vccd1
port 531 nsew power input
rlabel metal4 s 235794 281000 236414 284000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 281000 254414 284000 6 vccd1
port 531 nsew power input
rlabel metal4 s 271794 281000 272414 284000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 281000 290414 284000 6 vccd1
port 531 nsew power input
rlabel metal4 s 307794 281000 308414 284000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 281000 326414 284000 6 vccd1
port 531 nsew power input
rlabel metal4 s 343794 281000 344414 284000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 281000 362414 284000 6 vccd1
port 531 nsew power input
rlabel metal4 s 379794 281000 380414 284000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 281000 398414 284000 6 vccd1
port 531 nsew power input
rlabel metal4 s 415794 281000 416414 284000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 281000 434414 284000 6 vccd1
port 531 nsew power input
rlabel metal4 s 451794 281000 452414 284000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 281000 470414 284000 6 vccd1
port 531 nsew power input
rlabel metal4 s 487794 281000 488414 284000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 281000 506414 284000 6 vccd1
port 531 nsew power input
rlabel metal4 s 523794 281000 524414 284000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 281000 542414 284000 6 vccd1
port 531 nsew power input
rlabel metal4 s 19794 308000 20414 311000 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 308000 38414 311000 6 vccd1
port 531 nsew power input
rlabel metal4 s 55794 308000 56414 311000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 308000 74414 311000 6 vccd1
port 531 nsew power input
rlabel metal4 s 91794 308000 92414 311000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 308000 110414 311000 6 vccd1
port 531 nsew power input
rlabel metal4 s 127794 308000 128414 311000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 308000 146414 311000 6 vccd1
port 531 nsew power input
rlabel metal4 s 163794 308000 164414 311000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 308000 182414 311000 6 vccd1
port 531 nsew power input
rlabel metal4 s 199794 308000 200414 311000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 308000 218414 311000 6 vccd1
port 531 nsew power input
rlabel metal4 s 235794 308000 236414 311000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 308000 254414 311000 6 vccd1
port 531 nsew power input
rlabel metal4 s 271794 308000 272414 311000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 308000 290414 311000 6 vccd1
port 531 nsew power input
rlabel metal4 s 307794 308000 308414 311000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 308000 326414 311000 6 vccd1
port 531 nsew power input
rlabel metal4 s 343794 308000 344414 311000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 308000 362414 311000 6 vccd1
port 531 nsew power input
rlabel metal4 s 379794 308000 380414 311000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 308000 398414 311000 6 vccd1
port 531 nsew power input
rlabel metal4 s 415794 308000 416414 311000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 308000 434414 311000 6 vccd1
port 531 nsew power input
rlabel metal4 s 451794 308000 452414 311000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 308000 470414 311000 6 vccd1
port 531 nsew power input
rlabel metal4 s 487794 308000 488414 311000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 308000 506414 311000 6 vccd1
port 531 nsew power input
rlabel metal4 s 523794 308000 524414 311000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 308000 542414 311000 6 vccd1
port 531 nsew power input
rlabel metal4 s 19794 335000 20414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 335000 38414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 55794 335000 56414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 335000 74414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 91794 335000 92414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 335000 110414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 127794 335000 128414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 335000 146414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 163794 335000 164414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 335000 182414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 199794 335000 200414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 335000 218414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 235794 335000 236414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 335000 254414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 271794 335000 272414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 335000 290414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 307794 335000 308414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 335000 326414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 343794 335000 344414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 335000 362414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 379794 335000 380414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 335000 398414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 415794 335000 416414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 335000 434414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 451794 335000 452414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 335000 470414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 487794 335000 488414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 335000 506414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 523794 335000 524414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 335000 542414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 19794 362000 20414 365000 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 362000 38414 365000 6 vccd1
port 531 nsew power input
rlabel metal4 s 55794 362000 56414 365000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 362000 74414 365000 6 vccd1
port 531 nsew power input
rlabel metal4 s 91794 362000 92414 365000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 362000 110414 365000 6 vccd1
port 531 nsew power input
rlabel metal4 s 127794 362000 128414 365000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 362000 146414 365000 6 vccd1
port 531 nsew power input
rlabel metal4 s 163794 362000 164414 365000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 362000 182414 365000 6 vccd1
port 531 nsew power input
rlabel metal4 s 199794 362000 200414 365000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 362000 218414 365000 6 vccd1
port 531 nsew power input
rlabel metal4 s 235794 362000 236414 365000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 362000 254414 365000 6 vccd1
port 531 nsew power input
rlabel metal4 s 271794 362000 272414 365000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 362000 290414 365000 6 vccd1
port 531 nsew power input
rlabel metal4 s 307794 362000 308414 365000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 362000 326414 365000 6 vccd1
port 531 nsew power input
rlabel metal4 s 343794 362000 344414 365000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 362000 362414 365000 6 vccd1
port 531 nsew power input
rlabel metal4 s 379794 362000 380414 365000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 362000 398414 365000 6 vccd1
port 531 nsew power input
rlabel metal4 s 415794 362000 416414 365000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 362000 434414 365000 6 vccd1
port 531 nsew power input
rlabel metal4 s 451794 362000 452414 365000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 362000 470414 365000 6 vccd1
port 531 nsew power input
rlabel metal4 s 487794 362000 488414 365000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 362000 506414 365000 6 vccd1
port 531 nsew power input
rlabel metal4 s 523794 362000 524414 365000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 362000 542414 365000 6 vccd1
port 531 nsew power input
rlabel metal4 s 19794 389000 20414 392000 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 389000 38414 392000 6 vccd1
port 531 nsew power input
rlabel metal4 s 55794 389000 56414 392000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 389000 74414 392000 6 vccd1
port 531 nsew power input
rlabel metal4 s 91794 389000 92414 392000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 389000 110414 392000 6 vccd1
port 531 nsew power input
rlabel metal4 s 127794 389000 128414 392000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 389000 146414 392000 6 vccd1
port 531 nsew power input
rlabel metal4 s 163794 389000 164414 392000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 389000 182414 392000 6 vccd1
port 531 nsew power input
rlabel metal4 s 199794 389000 200414 392000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 389000 218414 392000 6 vccd1
port 531 nsew power input
rlabel metal4 s 235794 389000 236414 392000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 389000 254414 392000 6 vccd1
port 531 nsew power input
rlabel metal4 s 271794 389000 272414 392000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 389000 290414 392000 6 vccd1
port 531 nsew power input
rlabel metal4 s 307794 389000 308414 392000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 389000 326414 392000 6 vccd1
port 531 nsew power input
rlabel metal4 s 343794 389000 344414 392000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 389000 362414 392000 6 vccd1
port 531 nsew power input
rlabel metal4 s 379794 389000 380414 392000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 389000 398414 392000 6 vccd1
port 531 nsew power input
rlabel metal4 s 415794 389000 416414 392000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 389000 434414 392000 6 vccd1
port 531 nsew power input
rlabel metal4 s 451794 389000 452414 392000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 389000 470414 392000 6 vccd1
port 531 nsew power input
rlabel metal4 s 487794 389000 488414 392000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 389000 506414 392000 6 vccd1
port 531 nsew power input
rlabel metal4 s 523794 389000 524414 392000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 389000 542414 392000 6 vccd1
port 531 nsew power input
rlabel metal4 s 19794 416000 20414 419000 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 416000 38414 419000 6 vccd1
port 531 nsew power input
rlabel metal4 s 55794 416000 56414 419000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 416000 74414 419000 6 vccd1
port 531 nsew power input
rlabel metal4 s 91794 416000 92414 419000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 416000 110414 419000 6 vccd1
port 531 nsew power input
rlabel metal4 s 127794 416000 128414 419000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 416000 146414 419000 6 vccd1
port 531 nsew power input
rlabel metal4 s 163794 416000 164414 419000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 416000 182414 419000 6 vccd1
port 531 nsew power input
rlabel metal4 s 199794 416000 200414 419000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 416000 218414 419000 6 vccd1
port 531 nsew power input
rlabel metal4 s 235794 416000 236414 419000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 416000 254414 419000 6 vccd1
port 531 nsew power input
rlabel metal4 s 271794 416000 272414 419000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 416000 290414 419000 6 vccd1
port 531 nsew power input
rlabel metal4 s 307794 416000 308414 419000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 416000 326414 419000 6 vccd1
port 531 nsew power input
rlabel metal4 s 343794 416000 344414 419000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 416000 362414 419000 6 vccd1
port 531 nsew power input
rlabel metal4 s 379794 416000 380414 419000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 416000 398414 419000 6 vccd1
port 531 nsew power input
rlabel metal4 s 415794 416000 416414 419000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 416000 434414 419000 6 vccd1
port 531 nsew power input
rlabel metal4 s 451794 416000 452414 419000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 416000 470414 419000 6 vccd1
port 531 nsew power input
rlabel metal4 s 487794 416000 488414 419000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 416000 506414 419000 6 vccd1
port 531 nsew power input
rlabel metal4 s 523794 416000 524414 419000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 416000 542414 419000 6 vccd1
port 531 nsew power input
rlabel metal4 s 19794 443000 20414 446000 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 443000 38414 446000 6 vccd1
port 531 nsew power input
rlabel metal4 s 55794 443000 56414 446000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 443000 74414 446000 6 vccd1
port 531 nsew power input
rlabel metal4 s 91794 443000 92414 446000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 443000 110414 446000 6 vccd1
port 531 nsew power input
rlabel metal4 s 127794 443000 128414 446000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 443000 146414 446000 6 vccd1
port 531 nsew power input
rlabel metal4 s 163794 443000 164414 446000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 443000 182414 446000 6 vccd1
port 531 nsew power input
rlabel metal4 s 199794 443000 200414 446000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 443000 218414 446000 6 vccd1
port 531 nsew power input
rlabel metal4 s 235794 443000 236414 446000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 443000 254414 446000 6 vccd1
port 531 nsew power input
rlabel metal4 s 271794 443000 272414 446000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 443000 290414 446000 6 vccd1
port 531 nsew power input
rlabel metal4 s 307794 443000 308414 446000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 443000 326414 446000 6 vccd1
port 531 nsew power input
rlabel metal4 s 343794 443000 344414 446000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 443000 362414 446000 6 vccd1
port 531 nsew power input
rlabel metal4 s 379794 443000 380414 446000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 443000 398414 446000 6 vccd1
port 531 nsew power input
rlabel metal4 s 415794 443000 416414 446000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 443000 434414 446000 6 vccd1
port 531 nsew power input
rlabel metal4 s 451794 443000 452414 446000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 443000 470414 446000 6 vccd1
port 531 nsew power input
rlabel metal4 s 487794 443000 488414 446000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 443000 506414 446000 6 vccd1
port 531 nsew power input
rlabel metal4 s 523794 443000 524414 446000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 443000 542414 446000 6 vccd1
port 531 nsew power input
rlabel metal4 s 19794 470000 20414 473000 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 470000 38414 473000 6 vccd1
port 531 nsew power input
rlabel metal4 s 55794 470000 56414 473000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 470000 74414 473000 6 vccd1
port 531 nsew power input
rlabel metal4 s 91794 470000 92414 473000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 470000 110414 473000 6 vccd1
port 531 nsew power input
rlabel metal4 s 127794 470000 128414 473000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 470000 146414 473000 6 vccd1
port 531 nsew power input
rlabel metal4 s 163794 470000 164414 473000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 470000 182414 473000 6 vccd1
port 531 nsew power input
rlabel metal4 s 199794 470000 200414 473000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 470000 218414 473000 6 vccd1
port 531 nsew power input
rlabel metal4 s 235794 470000 236414 473000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 470000 254414 473000 6 vccd1
port 531 nsew power input
rlabel metal4 s 271794 470000 272414 473000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 470000 290414 473000 6 vccd1
port 531 nsew power input
rlabel metal4 s 307794 470000 308414 473000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 470000 326414 473000 6 vccd1
port 531 nsew power input
rlabel metal4 s 343794 470000 344414 473000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 470000 362414 473000 6 vccd1
port 531 nsew power input
rlabel metal4 s 379794 470000 380414 473000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 470000 398414 473000 6 vccd1
port 531 nsew power input
rlabel metal4 s 415794 470000 416414 473000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 470000 434414 473000 6 vccd1
port 531 nsew power input
rlabel metal4 s 451794 470000 452414 473000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 470000 470414 473000 6 vccd1
port 531 nsew power input
rlabel metal4 s 487794 470000 488414 473000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 470000 506414 473000 6 vccd1
port 531 nsew power input
rlabel metal4 s 523794 470000 524414 473000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 470000 542414 473000 6 vccd1
port 531 nsew power input
rlabel metal4 s 19794 497000 20414 500000 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 497000 38414 500000 6 vccd1
port 531 nsew power input
rlabel metal4 s 55794 497000 56414 500000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 497000 74414 500000 6 vccd1
port 531 nsew power input
rlabel metal4 s 91794 497000 92414 500000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 497000 110414 500000 6 vccd1
port 531 nsew power input
rlabel metal4 s 127794 497000 128414 500000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 497000 146414 500000 6 vccd1
port 531 nsew power input
rlabel metal4 s 163794 497000 164414 500000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 497000 182414 500000 6 vccd1
port 531 nsew power input
rlabel metal4 s 199794 497000 200414 500000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 497000 218414 500000 6 vccd1
port 531 nsew power input
rlabel metal4 s 235794 497000 236414 500000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 497000 254414 500000 6 vccd1
port 531 nsew power input
rlabel metal4 s 271794 497000 272414 500000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 497000 290414 500000 6 vccd1
port 531 nsew power input
rlabel metal4 s 307794 497000 308414 500000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 497000 326414 500000 6 vccd1
port 531 nsew power input
rlabel metal4 s 343794 497000 344414 500000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 497000 362414 500000 6 vccd1
port 531 nsew power input
rlabel metal4 s 379794 497000 380414 500000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 497000 398414 500000 6 vccd1
port 531 nsew power input
rlabel metal4 s 415794 497000 416414 500000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 497000 434414 500000 6 vccd1
port 531 nsew power input
rlabel metal4 s 451794 497000 452414 500000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 497000 470414 500000 6 vccd1
port 531 nsew power input
rlabel metal4 s 487794 497000 488414 500000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 497000 506414 500000 6 vccd1
port 531 nsew power input
rlabel metal4 s 523794 497000 524414 500000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 497000 542414 500000 6 vccd1
port 531 nsew power input
rlabel metal4 s 19794 524000 20414 527000 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 524000 38414 527000 6 vccd1
port 531 nsew power input
rlabel metal4 s 55794 524000 56414 527000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 524000 74414 527000 6 vccd1
port 531 nsew power input
rlabel metal4 s 91794 524000 92414 527000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 524000 110414 527000 6 vccd1
port 531 nsew power input
rlabel metal4 s 127794 524000 128414 527000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 524000 146414 527000 6 vccd1
port 531 nsew power input
rlabel metal4 s 163794 524000 164414 527000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 524000 182414 527000 6 vccd1
port 531 nsew power input
rlabel metal4 s 199794 524000 200414 527000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 524000 218414 527000 6 vccd1
port 531 nsew power input
rlabel metal4 s 235794 524000 236414 527000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 524000 254414 527000 6 vccd1
port 531 nsew power input
rlabel metal4 s 271794 524000 272414 527000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 524000 290414 527000 6 vccd1
port 531 nsew power input
rlabel metal4 s 307794 524000 308414 527000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 524000 326414 527000 6 vccd1
port 531 nsew power input
rlabel metal4 s 343794 524000 344414 527000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 524000 362414 527000 6 vccd1
port 531 nsew power input
rlabel metal4 s 379794 524000 380414 527000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 524000 398414 527000 6 vccd1
port 531 nsew power input
rlabel metal4 s 415794 524000 416414 527000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 524000 434414 527000 6 vccd1
port 531 nsew power input
rlabel metal4 s 451794 524000 452414 527000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 524000 470414 527000 6 vccd1
port 531 nsew power input
rlabel metal4 s 487794 524000 488414 527000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 524000 506414 527000 6 vccd1
port 531 nsew power input
rlabel metal4 s 523794 524000 524414 527000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 524000 542414 527000 6 vccd1
port 531 nsew power input
rlabel metal4 s 19794 551000 20414 554000 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 551000 38414 554000 6 vccd1
port 531 nsew power input
rlabel metal4 s 55794 551000 56414 554000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 551000 74414 554000 6 vccd1
port 531 nsew power input
rlabel metal4 s 91794 551000 92414 554000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 551000 110414 554000 6 vccd1
port 531 nsew power input
rlabel metal4 s 127794 551000 128414 554000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 551000 146414 554000 6 vccd1
port 531 nsew power input
rlabel metal4 s 163794 551000 164414 554000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 551000 182414 554000 6 vccd1
port 531 nsew power input
rlabel metal4 s 199794 551000 200414 554000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 551000 218414 554000 6 vccd1
port 531 nsew power input
rlabel metal4 s 235794 551000 236414 554000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 551000 254414 554000 6 vccd1
port 531 nsew power input
rlabel metal4 s 271794 551000 272414 554000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 551000 290414 554000 6 vccd1
port 531 nsew power input
rlabel metal4 s 307794 551000 308414 554000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 551000 326414 554000 6 vccd1
port 531 nsew power input
rlabel metal4 s 343794 551000 344414 554000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 551000 362414 554000 6 vccd1
port 531 nsew power input
rlabel metal4 s 379794 551000 380414 554000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 551000 398414 554000 6 vccd1
port 531 nsew power input
rlabel metal4 s 415794 551000 416414 554000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 551000 434414 554000 6 vccd1
port 531 nsew power input
rlabel metal4 s 451794 551000 452414 554000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 551000 470414 554000 6 vccd1
port 531 nsew power input
rlabel metal4 s 487794 551000 488414 554000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 551000 506414 554000 6 vccd1
port 531 nsew power input
rlabel metal4 s 523794 551000 524414 554000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 551000 542414 554000 6 vccd1
port 531 nsew power input
rlabel metal4 s 19794 578000 20414 581000 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 578000 38414 581000 6 vccd1
port 531 nsew power input
rlabel metal4 s 55794 578000 56414 581000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 578000 74414 581000 6 vccd1
port 531 nsew power input
rlabel metal4 s 91794 578000 92414 581000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 578000 110414 581000 6 vccd1
port 531 nsew power input
rlabel metal4 s 127794 578000 128414 581000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 578000 146414 581000 6 vccd1
port 531 nsew power input
rlabel metal4 s 163794 578000 164414 581000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 578000 182414 581000 6 vccd1
port 531 nsew power input
rlabel metal4 s 199794 578000 200414 581000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 578000 218414 581000 6 vccd1
port 531 nsew power input
rlabel metal4 s 235794 578000 236414 581000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 578000 254414 581000 6 vccd1
port 531 nsew power input
rlabel metal4 s 271794 578000 272414 581000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 578000 290414 581000 6 vccd1
port 531 nsew power input
rlabel metal4 s 307794 578000 308414 581000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 578000 326414 581000 6 vccd1
port 531 nsew power input
rlabel metal4 s 343794 578000 344414 581000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 578000 362414 581000 6 vccd1
port 531 nsew power input
rlabel metal4 s 379794 578000 380414 581000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 578000 398414 581000 6 vccd1
port 531 nsew power input
rlabel metal4 s 415794 578000 416414 581000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 578000 434414 581000 6 vccd1
port 531 nsew power input
rlabel metal4 s 451794 578000 452414 581000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 578000 470414 581000 6 vccd1
port 531 nsew power input
rlabel metal4 s 487794 578000 488414 581000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 578000 506414 581000 6 vccd1
port 531 nsew power input
rlabel metal4 s 523794 578000 524414 581000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 578000 542414 581000 6 vccd1
port 531 nsew power input
rlabel metal4 s 19794 605000 20414 608000 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 605000 38414 608000 6 vccd1
port 531 nsew power input
rlabel metal4 s 55794 605000 56414 608000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 605000 74414 608000 6 vccd1
port 531 nsew power input
rlabel metal4 s 91794 605000 92414 608000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 605000 110414 608000 6 vccd1
port 531 nsew power input
rlabel metal4 s 127794 605000 128414 608000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 605000 146414 608000 6 vccd1
port 531 nsew power input
rlabel metal4 s 163794 605000 164414 608000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 605000 182414 608000 6 vccd1
port 531 nsew power input
rlabel metal4 s 199794 605000 200414 608000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 605000 218414 608000 6 vccd1
port 531 nsew power input
rlabel metal4 s 235794 605000 236414 608000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 605000 254414 608000 6 vccd1
port 531 nsew power input
rlabel metal4 s 271794 605000 272414 608000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 605000 290414 608000 6 vccd1
port 531 nsew power input
rlabel metal4 s 307794 605000 308414 608000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 605000 326414 608000 6 vccd1
port 531 nsew power input
rlabel metal4 s 343794 605000 344414 608000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 605000 362414 608000 6 vccd1
port 531 nsew power input
rlabel metal4 s 379794 605000 380414 608000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 605000 398414 608000 6 vccd1
port 531 nsew power input
rlabel metal4 s 415794 605000 416414 608000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 605000 434414 608000 6 vccd1
port 531 nsew power input
rlabel metal4 s 451794 605000 452414 608000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 605000 470414 608000 6 vccd1
port 531 nsew power input
rlabel metal4 s 487794 605000 488414 608000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 605000 506414 608000 6 vccd1
port 531 nsew power input
rlabel metal4 s 523794 605000 524414 608000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 605000 542414 608000 6 vccd1
port 531 nsew power input
rlabel metal4 s 19794 632000 20414 635000 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 632000 38414 635000 6 vccd1
port 531 nsew power input
rlabel metal4 s 55794 632000 56414 635000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 632000 74414 635000 6 vccd1
port 531 nsew power input
rlabel metal4 s 91794 632000 92414 635000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 632000 110414 635000 6 vccd1
port 531 nsew power input
rlabel metal4 s 127794 632000 128414 635000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 632000 146414 635000 6 vccd1
port 531 nsew power input
rlabel metal4 s 163794 632000 164414 635000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 632000 182414 635000 6 vccd1
port 531 nsew power input
rlabel metal4 s 199794 632000 200414 635000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 632000 218414 635000 6 vccd1
port 531 nsew power input
rlabel metal4 s 235794 632000 236414 635000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 632000 254414 635000 6 vccd1
port 531 nsew power input
rlabel metal4 s 271794 632000 272414 635000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 632000 290414 635000 6 vccd1
port 531 nsew power input
rlabel metal4 s 307794 632000 308414 635000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 632000 326414 635000 6 vccd1
port 531 nsew power input
rlabel metal4 s 343794 632000 344414 635000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 632000 362414 635000 6 vccd1
port 531 nsew power input
rlabel metal4 s 379794 632000 380414 635000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 632000 398414 635000 6 vccd1
port 531 nsew power input
rlabel metal4 s 415794 632000 416414 635000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 632000 434414 635000 6 vccd1
port 531 nsew power input
rlabel metal4 s 451794 632000 452414 635000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 632000 470414 635000 6 vccd1
port 531 nsew power input
rlabel metal4 s 487794 632000 488414 635000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 632000 506414 635000 6 vccd1
port 531 nsew power input
rlabel metal4 s 523794 632000 524414 635000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 632000 542414 635000 6 vccd1
port 531 nsew power input
rlabel metal4 s 19794 659000 20414 662000 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 659000 38414 662000 6 vccd1
port 531 nsew power input
rlabel metal4 s 55794 659000 56414 662000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 659000 74414 662000 6 vccd1
port 531 nsew power input
rlabel metal4 s 91794 659000 92414 662000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 659000 110414 662000 6 vccd1
port 531 nsew power input
rlabel metal4 s 127794 659000 128414 662000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 659000 146414 662000 6 vccd1
port 531 nsew power input
rlabel metal4 s 163794 659000 164414 662000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 659000 182414 662000 6 vccd1
port 531 nsew power input
rlabel metal4 s 199794 659000 200414 662000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 659000 218414 662000 6 vccd1
port 531 nsew power input
rlabel metal4 s 235794 659000 236414 662000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 659000 254414 662000 6 vccd1
port 531 nsew power input
rlabel metal4 s 271794 659000 272414 662000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 659000 290414 662000 6 vccd1
port 531 nsew power input
rlabel metal4 s 307794 659000 308414 662000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 659000 326414 662000 6 vccd1
port 531 nsew power input
rlabel metal4 s 343794 659000 344414 662000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 659000 362414 662000 6 vccd1
port 531 nsew power input
rlabel metal4 s 379794 659000 380414 662000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 659000 398414 662000 6 vccd1
port 531 nsew power input
rlabel metal4 s 415794 659000 416414 662000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 659000 434414 662000 6 vccd1
port 531 nsew power input
rlabel metal4 s 451794 659000 452414 662000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 659000 470414 662000 6 vccd1
port 531 nsew power input
rlabel metal4 s 487794 659000 488414 662000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 659000 506414 662000 6 vccd1
port 531 nsew power input
rlabel metal4 s 523794 659000 524414 662000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 659000 542414 662000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 19794 686000 20414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 686000 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 55794 686000 56414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 686000 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 91794 686000 92414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 686000 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 127794 686000 128414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 686000 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 163794 686000 164414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 686000 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 199794 686000 200414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 686000 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 235794 686000 236414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 686000 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 271794 686000 272414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 686000 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 307794 686000 308414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 686000 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 343794 686000 344414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 686000 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 379794 686000 380414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 686000 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 415794 686000 416414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 686000 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 451794 686000 452414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 686000 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 487794 686000 488414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 686000 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 523794 686000 524414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 686000 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 559794 -1894 560414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 11866 586890 12486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 29866 586890 30486 6 vssd1
port 532 nsew ground input
rlabel metal5 s 28794 39806 551414 40426 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 47866 586890 48486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 65866 586890 66486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 83866 586890 84486 6 vssd1
port 532 nsew ground input
rlabel metal5 s 28794 93806 551414 94426 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 101866 586890 102486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 119866 586890 120486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 137866 586890 138486 6 vssd1
port 532 nsew ground input
rlabel metal5 s 28794 147806 551414 148426 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 155866 586890 156486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 173866 586890 174486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 191866 586890 192486 6 vssd1
port 532 nsew ground input
rlabel metal5 s 28794 201806 551414 202426 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 209866 586890 210486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 227866 586890 228486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 245866 586890 246486 6 vssd1
port 532 nsew ground input
rlabel metal5 s 28794 255806 551414 256426 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 263866 586890 264486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 281866 586890 282486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 299866 586890 300486 6 vssd1
port 532 nsew ground input
rlabel metal5 s 28794 309806 551414 310426 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 317866 586890 318486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 335866 586890 336486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 353866 586890 354486 6 vssd1
port 532 nsew ground input
rlabel metal5 s 28794 363806 551414 364426 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 371866 586890 372486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 389866 586890 390486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 407866 586890 408486 6 vssd1
port 532 nsew ground input
rlabel metal5 s 28794 417806 551414 418426 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 425866 586890 426486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 443866 586890 444486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 461866 586890 462486 6 vssd1
port 532 nsew ground input
rlabel metal5 s 28794 471806 551414 472426 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 479866 586890 480486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 497866 586890 498486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 515866 586890 516486 6 vssd1
port 532 nsew ground input
rlabel metal5 s 28794 525806 551414 526426 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 533866 586890 534486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 551866 586890 552486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 569866 586890 570486 6 vssd1
port 532 nsew ground input
rlabel metal5 s 28794 579806 551414 580426 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 587866 586890 588486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 605866 586890 606486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 623866 586890 624486 6 vssd1
port 532 nsew ground input
rlabel metal5 s 28794 633806 551414 634426 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 641866 586890 642486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 659866 586890 660486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 677866 586890 678486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 695866 586890 696486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 28794 -1894 29414 14000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 46794 -1894 47414 14000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 64794 -1894 65414 14000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 82794 -1894 83414 14000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 100794 -1894 101414 14000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 118794 -1894 119414 14000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 136794 -1894 137414 14000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 154794 -1894 155414 14000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 172794 -1894 173414 14000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 190794 -1894 191414 14000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 208794 -1894 209414 14000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 226794 -1894 227414 14000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 244794 -1894 245414 14000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 262794 -1894 263414 14000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 280794 -1894 281414 14000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 298794 -1894 299414 14000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 316794 -1894 317414 14000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 334794 -1894 335414 14000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 352794 -1894 353414 14000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 370794 -1894 371414 14000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 388794 -1894 389414 14000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 406794 -1894 407414 14000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 424794 -1894 425414 14000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 442794 -1894 443414 14000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 460794 -1894 461414 14000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 478794 -1894 479414 14000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 496794 -1894 497414 14000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 514794 -1894 515414 14000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 532794 -1894 533414 14000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 550794 -1894 551414 14000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 28794 38000 29414 41000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 46794 38000 47414 41000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 64794 38000 65414 41000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 82794 38000 83414 41000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 100794 38000 101414 41000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 118794 38000 119414 41000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 136794 38000 137414 41000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 154794 38000 155414 41000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 172794 38000 173414 41000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 190794 38000 191414 41000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 208794 38000 209414 41000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 226794 38000 227414 41000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 244794 38000 245414 41000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 262794 38000 263414 41000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 280794 38000 281414 41000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 298794 38000 299414 41000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 316794 38000 317414 41000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 334794 38000 335414 41000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 352794 38000 353414 41000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 370794 38000 371414 41000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 388794 38000 389414 41000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 406794 38000 407414 41000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 424794 38000 425414 41000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 442794 38000 443414 41000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 460794 38000 461414 41000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 478794 38000 479414 41000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 496794 38000 497414 41000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 514794 38000 515414 41000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 532794 38000 533414 41000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 550794 38000 551414 41000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 28794 65000 29414 68000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 46794 65000 47414 68000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 64794 65000 65414 68000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 82794 65000 83414 68000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 100794 65000 101414 68000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 118794 65000 119414 68000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 136794 65000 137414 68000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 154794 65000 155414 68000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 172794 65000 173414 68000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 190794 65000 191414 68000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 208794 65000 209414 68000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 226794 65000 227414 68000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 244794 65000 245414 68000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 262794 65000 263414 68000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 280794 65000 281414 68000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 298794 65000 299414 68000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 316794 65000 317414 68000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 334794 65000 335414 68000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 352794 65000 353414 68000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 370794 65000 371414 68000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 388794 65000 389414 68000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 406794 65000 407414 68000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 424794 65000 425414 68000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 442794 65000 443414 68000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 460794 65000 461414 68000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 478794 65000 479414 68000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 496794 65000 497414 68000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 514794 65000 515414 68000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 532794 65000 533414 68000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 550794 65000 551414 68000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 28794 92000 29414 95000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 46794 92000 47414 95000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 64794 92000 65414 95000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 82794 92000 83414 95000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 100794 92000 101414 95000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 118794 92000 119414 95000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 136794 92000 137414 95000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 154794 92000 155414 95000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 172794 92000 173414 95000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 190794 92000 191414 95000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 208794 92000 209414 95000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 226794 92000 227414 95000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 244794 92000 245414 95000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 262794 92000 263414 95000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 280794 92000 281414 95000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 298794 92000 299414 95000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 316794 92000 317414 95000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 334794 92000 335414 95000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 352794 92000 353414 95000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 370794 92000 371414 95000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 388794 92000 389414 95000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 406794 92000 407414 95000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 424794 92000 425414 95000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 442794 92000 443414 95000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 460794 92000 461414 95000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 478794 92000 479414 95000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 496794 92000 497414 95000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 514794 92000 515414 95000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 532794 92000 533414 95000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 550794 92000 551414 95000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 28794 119000 29414 122000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 46794 119000 47414 122000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 64794 119000 65414 122000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 82794 119000 83414 122000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 100794 119000 101414 122000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 118794 119000 119414 122000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 136794 119000 137414 122000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 154794 119000 155414 122000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 172794 119000 173414 122000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 190794 119000 191414 122000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 208794 119000 209414 122000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 226794 119000 227414 122000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 244794 119000 245414 122000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 262794 119000 263414 122000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 280794 119000 281414 122000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 298794 119000 299414 122000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 316794 119000 317414 122000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 334794 119000 335414 122000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 352794 119000 353414 122000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 370794 119000 371414 122000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 388794 119000 389414 122000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 406794 119000 407414 122000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 424794 119000 425414 122000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 442794 119000 443414 122000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 460794 119000 461414 122000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 478794 119000 479414 122000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 496794 119000 497414 122000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 514794 119000 515414 122000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 532794 119000 533414 122000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 550794 119000 551414 122000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 28794 146000 29414 149000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 46794 146000 47414 149000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 64794 146000 65414 149000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 82794 146000 83414 149000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 100794 146000 101414 149000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 118794 146000 119414 149000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 136794 146000 137414 149000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 154794 146000 155414 149000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 172794 146000 173414 149000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 190794 146000 191414 149000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 208794 146000 209414 149000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 226794 146000 227414 149000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 244794 146000 245414 149000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 262794 146000 263414 149000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 280794 146000 281414 149000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 298794 146000 299414 149000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 316794 146000 317414 149000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 334794 146000 335414 149000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 352794 146000 353414 149000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 370794 146000 371414 149000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 388794 146000 389414 149000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 406794 146000 407414 149000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 424794 146000 425414 149000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 442794 146000 443414 149000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 460794 146000 461414 149000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 478794 146000 479414 149000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 496794 146000 497414 149000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 514794 146000 515414 149000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 532794 146000 533414 149000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 550794 146000 551414 149000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 28794 173000 29414 176000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 46794 173000 47414 176000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 64794 173000 65414 176000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 82794 173000 83414 176000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 100794 173000 101414 176000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 118794 173000 119414 176000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 136794 173000 137414 176000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 154794 173000 155414 176000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 172794 173000 173414 176000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 190794 173000 191414 176000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 208794 173000 209414 176000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 226794 173000 227414 176000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 244794 173000 245414 176000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 262794 173000 263414 176000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 280794 173000 281414 176000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 298794 173000 299414 176000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 316794 173000 317414 176000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 334794 173000 335414 176000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 352794 173000 353414 176000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 370794 173000 371414 176000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 388794 173000 389414 176000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 406794 173000 407414 176000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 424794 173000 425414 176000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 442794 173000 443414 176000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 460794 173000 461414 176000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 478794 173000 479414 176000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 496794 173000 497414 176000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 514794 173000 515414 176000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 532794 173000 533414 176000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 550794 173000 551414 176000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 28794 200000 29414 203000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 46794 200000 47414 203000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 64794 200000 65414 203000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 82794 200000 83414 203000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 100794 200000 101414 203000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 118794 200000 119414 203000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 136794 200000 137414 203000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 154794 200000 155414 203000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 172794 200000 173414 203000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 190794 200000 191414 203000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 208794 200000 209414 203000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 226794 200000 227414 203000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 244794 200000 245414 203000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 262794 200000 263414 203000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 280794 200000 281414 203000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 298794 200000 299414 203000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 316794 200000 317414 203000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 334794 200000 335414 203000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 352794 200000 353414 203000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 370794 200000 371414 203000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 388794 200000 389414 203000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 406794 200000 407414 203000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 424794 200000 425414 203000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 442794 200000 443414 203000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 460794 200000 461414 203000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 478794 200000 479414 203000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 496794 200000 497414 203000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 514794 200000 515414 203000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 532794 200000 533414 203000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 550794 200000 551414 203000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 28794 227000 29414 230000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 46794 227000 47414 230000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 64794 227000 65414 230000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 82794 227000 83414 230000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 100794 227000 101414 230000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 118794 227000 119414 230000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 136794 227000 137414 230000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 154794 227000 155414 230000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 172794 227000 173414 230000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 190794 227000 191414 230000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 208794 227000 209414 230000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 226794 227000 227414 230000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 244794 227000 245414 230000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 262794 227000 263414 230000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 280794 227000 281414 230000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 298794 227000 299414 230000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 316794 227000 317414 230000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 334794 227000 335414 230000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 352794 227000 353414 230000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 370794 227000 371414 230000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 388794 227000 389414 230000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 406794 227000 407414 230000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 424794 227000 425414 230000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 442794 227000 443414 230000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 460794 227000 461414 230000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 478794 227000 479414 230000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 496794 227000 497414 230000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 514794 227000 515414 230000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 532794 227000 533414 230000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 550794 227000 551414 230000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 28794 254000 29414 257000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 46794 254000 47414 257000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 64794 254000 65414 257000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 82794 254000 83414 257000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 100794 254000 101414 257000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 118794 254000 119414 257000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 136794 254000 137414 257000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 154794 254000 155414 257000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 172794 254000 173414 257000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 190794 254000 191414 257000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 208794 254000 209414 257000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 226794 254000 227414 257000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 244794 254000 245414 257000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 262794 254000 263414 257000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 280794 254000 281414 257000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 298794 254000 299414 257000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 316794 254000 317414 257000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 334794 254000 335414 257000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 352794 254000 353414 257000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 370794 254000 371414 257000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 388794 254000 389414 257000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 406794 254000 407414 257000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 424794 254000 425414 257000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 442794 254000 443414 257000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 460794 254000 461414 257000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 478794 254000 479414 257000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 496794 254000 497414 257000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 514794 254000 515414 257000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 532794 254000 533414 257000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 550794 254000 551414 257000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 28794 281000 29414 284000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 46794 281000 47414 284000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 64794 281000 65414 284000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 82794 281000 83414 284000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 100794 281000 101414 284000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 118794 281000 119414 284000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 136794 281000 137414 284000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 154794 281000 155414 284000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 172794 281000 173414 284000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 190794 281000 191414 284000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 208794 281000 209414 284000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 226794 281000 227414 284000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 244794 281000 245414 284000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 262794 281000 263414 284000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 280794 281000 281414 284000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 298794 281000 299414 284000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 316794 281000 317414 284000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 334794 281000 335414 284000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 352794 281000 353414 284000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 370794 281000 371414 284000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 388794 281000 389414 284000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 406794 281000 407414 284000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 424794 281000 425414 284000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 442794 281000 443414 284000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 460794 281000 461414 284000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 478794 281000 479414 284000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 496794 281000 497414 284000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 514794 281000 515414 284000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 532794 281000 533414 284000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 550794 281000 551414 284000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 28794 308000 29414 311000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 46794 308000 47414 311000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 64794 308000 65414 311000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 82794 308000 83414 311000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 100794 308000 101414 311000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 118794 308000 119414 311000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 136794 308000 137414 311000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 154794 308000 155414 311000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 172794 308000 173414 311000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 190794 308000 191414 311000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 208794 308000 209414 311000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 226794 308000 227414 311000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 244794 308000 245414 311000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 262794 308000 263414 311000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 280794 308000 281414 311000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 298794 308000 299414 311000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 316794 308000 317414 311000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 334794 308000 335414 311000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 352794 308000 353414 311000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 370794 308000 371414 311000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 388794 308000 389414 311000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 406794 308000 407414 311000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 424794 308000 425414 311000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 442794 308000 443414 311000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 460794 308000 461414 311000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 478794 308000 479414 311000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 496794 308000 497414 311000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 514794 308000 515414 311000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 532794 308000 533414 311000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 550794 308000 551414 311000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 28794 335000 29414 338000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 46794 335000 47414 338000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 64794 335000 65414 338000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 82794 335000 83414 338000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 100794 335000 101414 338000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 118794 335000 119414 338000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 136794 335000 137414 338000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 154794 335000 155414 338000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 172794 335000 173414 338000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 190794 335000 191414 338000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 208794 335000 209414 338000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 226794 335000 227414 338000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 244794 335000 245414 338000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 262794 335000 263414 338000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 280794 335000 281414 338000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 298794 335000 299414 338000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 316794 335000 317414 338000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 334794 335000 335414 338000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 352794 335000 353414 338000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 370794 335000 371414 338000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 388794 335000 389414 338000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 406794 335000 407414 338000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 424794 335000 425414 338000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 442794 335000 443414 338000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 460794 335000 461414 338000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 478794 335000 479414 338000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 496794 335000 497414 338000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 514794 335000 515414 338000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 532794 335000 533414 338000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 550794 335000 551414 338000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 28794 362000 29414 365000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 46794 362000 47414 365000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 64794 362000 65414 365000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 82794 362000 83414 365000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 100794 362000 101414 365000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 118794 362000 119414 365000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 136794 362000 137414 365000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 154794 362000 155414 365000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 172794 362000 173414 365000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 190794 362000 191414 365000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 208794 362000 209414 365000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 226794 362000 227414 365000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 244794 362000 245414 365000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 262794 362000 263414 365000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 280794 362000 281414 365000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 298794 362000 299414 365000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 316794 362000 317414 365000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 334794 362000 335414 365000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 352794 362000 353414 365000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 370794 362000 371414 365000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 388794 362000 389414 365000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 406794 362000 407414 365000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 424794 362000 425414 365000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 442794 362000 443414 365000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 460794 362000 461414 365000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 478794 362000 479414 365000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 496794 362000 497414 365000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 514794 362000 515414 365000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 532794 362000 533414 365000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 550794 362000 551414 365000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 28794 389000 29414 392000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 46794 389000 47414 392000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 64794 389000 65414 392000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 82794 389000 83414 392000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 100794 389000 101414 392000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 118794 389000 119414 392000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 136794 389000 137414 392000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 154794 389000 155414 392000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 172794 389000 173414 392000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 190794 389000 191414 392000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 208794 389000 209414 392000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 226794 389000 227414 392000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 244794 389000 245414 392000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 262794 389000 263414 392000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 280794 389000 281414 392000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 298794 389000 299414 392000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 316794 389000 317414 392000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 334794 389000 335414 392000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 352794 389000 353414 392000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 370794 389000 371414 392000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 388794 389000 389414 392000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 406794 389000 407414 392000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 424794 389000 425414 392000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 442794 389000 443414 392000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 460794 389000 461414 392000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 478794 389000 479414 392000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 496794 389000 497414 392000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 514794 389000 515414 392000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 532794 389000 533414 392000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 550794 389000 551414 392000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 28794 416000 29414 419000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 46794 416000 47414 419000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 64794 416000 65414 419000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 82794 416000 83414 419000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 100794 416000 101414 419000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 118794 416000 119414 419000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 136794 416000 137414 419000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 154794 416000 155414 419000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 172794 416000 173414 419000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 190794 416000 191414 419000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 208794 416000 209414 419000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 226794 416000 227414 419000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 244794 416000 245414 419000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 262794 416000 263414 419000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 280794 416000 281414 419000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 298794 416000 299414 419000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 316794 416000 317414 419000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 334794 416000 335414 419000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 352794 416000 353414 419000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 370794 416000 371414 419000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 388794 416000 389414 419000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 406794 416000 407414 419000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 424794 416000 425414 419000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 442794 416000 443414 419000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 460794 416000 461414 419000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 478794 416000 479414 419000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 496794 416000 497414 419000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 514794 416000 515414 419000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 532794 416000 533414 419000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 550794 416000 551414 419000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 28794 443000 29414 446000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 46794 443000 47414 446000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 64794 443000 65414 446000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 82794 443000 83414 446000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 100794 443000 101414 446000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 118794 443000 119414 446000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 136794 443000 137414 446000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 154794 443000 155414 446000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 172794 443000 173414 446000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 190794 443000 191414 446000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 208794 443000 209414 446000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 226794 443000 227414 446000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 244794 443000 245414 446000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 262794 443000 263414 446000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 280794 443000 281414 446000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 298794 443000 299414 446000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 316794 443000 317414 446000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 334794 443000 335414 446000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 352794 443000 353414 446000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 370794 443000 371414 446000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 388794 443000 389414 446000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 406794 443000 407414 446000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 424794 443000 425414 446000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 442794 443000 443414 446000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 460794 443000 461414 446000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 478794 443000 479414 446000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 496794 443000 497414 446000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 514794 443000 515414 446000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 532794 443000 533414 446000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 550794 443000 551414 446000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 28794 470000 29414 473000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 46794 470000 47414 473000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 64794 470000 65414 473000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 82794 470000 83414 473000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 100794 470000 101414 473000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 118794 470000 119414 473000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 136794 470000 137414 473000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 154794 470000 155414 473000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 172794 470000 173414 473000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 190794 470000 191414 473000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 208794 470000 209414 473000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 226794 470000 227414 473000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 244794 470000 245414 473000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 262794 470000 263414 473000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 280794 470000 281414 473000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 298794 470000 299414 473000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 316794 470000 317414 473000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 334794 470000 335414 473000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 352794 470000 353414 473000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 370794 470000 371414 473000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 388794 470000 389414 473000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 406794 470000 407414 473000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 424794 470000 425414 473000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 442794 470000 443414 473000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 460794 470000 461414 473000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 478794 470000 479414 473000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 496794 470000 497414 473000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 514794 470000 515414 473000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 532794 470000 533414 473000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 550794 470000 551414 473000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 28794 497000 29414 500000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 46794 497000 47414 500000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 64794 497000 65414 500000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 82794 497000 83414 500000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 100794 497000 101414 500000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 118794 497000 119414 500000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 136794 497000 137414 500000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 154794 497000 155414 500000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 172794 497000 173414 500000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 190794 497000 191414 500000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 208794 497000 209414 500000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 226794 497000 227414 500000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 244794 497000 245414 500000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 262794 497000 263414 500000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 280794 497000 281414 500000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 298794 497000 299414 500000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 316794 497000 317414 500000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 334794 497000 335414 500000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 352794 497000 353414 500000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 370794 497000 371414 500000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 388794 497000 389414 500000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 406794 497000 407414 500000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 424794 497000 425414 500000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 442794 497000 443414 500000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 460794 497000 461414 500000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 478794 497000 479414 500000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 496794 497000 497414 500000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 514794 497000 515414 500000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 532794 497000 533414 500000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 550794 497000 551414 500000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 28794 524000 29414 527000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 46794 524000 47414 527000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 64794 524000 65414 527000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 82794 524000 83414 527000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 100794 524000 101414 527000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 118794 524000 119414 527000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 136794 524000 137414 527000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 154794 524000 155414 527000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 172794 524000 173414 527000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 190794 524000 191414 527000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 208794 524000 209414 527000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 226794 524000 227414 527000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 244794 524000 245414 527000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 262794 524000 263414 527000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 280794 524000 281414 527000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 298794 524000 299414 527000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 316794 524000 317414 527000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 334794 524000 335414 527000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 352794 524000 353414 527000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 370794 524000 371414 527000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 388794 524000 389414 527000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 406794 524000 407414 527000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 424794 524000 425414 527000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 442794 524000 443414 527000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 460794 524000 461414 527000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 478794 524000 479414 527000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 496794 524000 497414 527000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 514794 524000 515414 527000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 532794 524000 533414 527000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 550794 524000 551414 527000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 28794 551000 29414 554000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 46794 551000 47414 554000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 64794 551000 65414 554000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 82794 551000 83414 554000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 100794 551000 101414 554000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 118794 551000 119414 554000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 136794 551000 137414 554000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 154794 551000 155414 554000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 172794 551000 173414 554000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 190794 551000 191414 554000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 208794 551000 209414 554000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 226794 551000 227414 554000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 244794 551000 245414 554000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 262794 551000 263414 554000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 280794 551000 281414 554000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 298794 551000 299414 554000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 316794 551000 317414 554000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 334794 551000 335414 554000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 352794 551000 353414 554000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 370794 551000 371414 554000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 388794 551000 389414 554000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 406794 551000 407414 554000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 424794 551000 425414 554000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 442794 551000 443414 554000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 460794 551000 461414 554000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 478794 551000 479414 554000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 496794 551000 497414 554000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 514794 551000 515414 554000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 532794 551000 533414 554000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 550794 551000 551414 554000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 28794 578000 29414 581000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 46794 578000 47414 581000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 64794 578000 65414 581000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 82794 578000 83414 581000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 100794 578000 101414 581000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 118794 578000 119414 581000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 136794 578000 137414 581000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 154794 578000 155414 581000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 172794 578000 173414 581000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 190794 578000 191414 581000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 208794 578000 209414 581000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 226794 578000 227414 581000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 244794 578000 245414 581000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 262794 578000 263414 581000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 280794 578000 281414 581000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 298794 578000 299414 581000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 316794 578000 317414 581000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 334794 578000 335414 581000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 352794 578000 353414 581000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 370794 578000 371414 581000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 388794 578000 389414 581000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 406794 578000 407414 581000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 424794 578000 425414 581000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 442794 578000 443414 581000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 460794 578000 461414 581000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 478794 578000 479414 581000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 496794 578000 497414 581000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 514794 578000 515414 581000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 532794 578000 533414 581000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 550794 578000 551414 581000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 28794 605000 29414 608000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 46794 605000 47414 608000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 64794 605000 65414 608000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 82794 605000 83414 608000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 100794 605000 101414 608000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 118794 605000 119414 608000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 136794 605000 137414 608000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 154794 605000 155414 608000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 172794 605000 173414 608000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 190794 605000 191414 608000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 208794 605000 209414 608000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 226794 605000 227414 608000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 244794 605000 245414 608000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 262794 605000 263414 608000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 280794 605000 281414 608000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 298794 605000 299414 608000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 316794 605000 317414 608000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 334794 605000 335414 608000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 352794 605000 353414 608000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 370794 605000 371414 608000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 388794 605000 389414 608000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 406794 605000 407414 608000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 424794 605000 425414 608000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 442794 605000 443414 608000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 460794 605000 461414 608000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 478794 605000 479414 608000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 496794 605000 497414 608000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 514794 605000 515414 608000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 532794 605000 533414 608000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 550794 605000 551414 608000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 28794 632000 29414 635000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 46794 632000 47414 635000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 64794 632000 65414 635000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 82794 632000 83414 635000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 100794 632000 101414 635000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 118794 632000 119414 635000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 136794 632000 137414 635000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 154794 632000 155414 635000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 172794 632000 173414 635000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 190794 632000 191414 635000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 208794 632000 209414 635000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 226794 632000 227414 635000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 244794 632000 245414 635000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 262794 632000 263414 635000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 280794 632000 281414 635000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 298794 632000 299414 635000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 316794 632000 317414 635000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 334794 632000 335414 635000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 352794 632000 353414 635000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 370794 632000 371414 635000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 388794 632000 389414 635000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 406794 632000 407414 635000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 424794 632000 425414 635000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 442794 632000 443414 635000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 460794 632000 461414 635000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 478794 632000 479414 635000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 496794 632000 497414 635000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 514794 632000 515414 635000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 532794 632000 533414 635000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 550794 632000 551414 635000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 28794 659000 29414 662000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 46794 659000 47414 662000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 64794 659000 65414 662000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 82794 659000 83414 662000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 100794 659000 101414 662000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 118794 659000 119414 662000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 136794 659000 137414 662000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 154794 659000 155414 662000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 172794 659000 173414 662000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 190794 659000 191414 662000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 208794 659000 209414 662000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 226794 659000 227414 662000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 244794 659000 245414 662000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 262794 659000 263414 662000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 280794 659000 281414 662000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 298794 659000 299414 662000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 316794 659000 317414 662000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 334794 659000 335414 662000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 352794 659000 353414 662000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 370794 659000 371414 662000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 388794 659000 389414 662000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 406794 659000 407414 662000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 424794 659000 425414 662000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 442794 659000 443414 662000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 460794 659000 461414 662000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 478794 659000 479414 662000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 496794 659000 497414 662000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 514794 659000 515414 662000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 532794 659000 533414 662000 6 vssd1
port 532 nsew ground input
rlabel metal4 s 550794 659000 551414 662000 6 vssd1
port 532 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 532 nsew ground input
rlabel metal4 s 10794 -1894 11414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 28794 686000 29414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 46794 686000 47414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 64794 686000 65414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 82794 686000 83414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 100794 686000 101414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 118794 686000 119414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 136794 686000 137414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 154794 686000 155414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 172794 686000 173414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 190794 686000 191414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 208794 686000 209414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 226794 686000 227414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 244794 686000 245414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 262794 686000 263414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 280794 686000 281414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 298794 686000 299414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 316794 686000 317414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 334794 686000 335414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 352794 686000 353414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 370794 686000 371414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 388794 686000 389414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 406794 686000 407414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 424794 686000 425414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 442794 686000 443414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 460794 686000 461414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 478794 686000 479414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 496794 686000 497414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 514794 686000 515414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 532794 686000 533414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 550794 686000 551414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 568794 -1894 569414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 532 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 533 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 534 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 535 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 536 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 537 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 538 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 539 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 540 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 541 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 542 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 543 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 544 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 545 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 546 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 547 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 548 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 549 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 550 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 551 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 552 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 553 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 554 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 555 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 556 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 557 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 558 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 559 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 560 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 561 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 562 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 563 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 564 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 565 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 566 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 567 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 568 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 569 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 570 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 571 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 572 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 573 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 574 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 575 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 576 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 577 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 578 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 579 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 580 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 581 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 582 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 583 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 584 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 585 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 586 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 587 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 588 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 589 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 590 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 591 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 592 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 593 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 594 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 595 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 596 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 597 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 598 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 599 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 600 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 601 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 602 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 603 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 604 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 605 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 606 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 607 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 608 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 609 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 610 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 611 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 612 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 613 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 614 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 615 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 616 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 617 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 618 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 619 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 620 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 621 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 622 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 623 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 624 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 625 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 626 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 627 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 628 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 629 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 630 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 631 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 632 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 633 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 634 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 635 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 636 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 637 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 638 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
